module real_aes_2712_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_0), .B(n_151), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_159), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_2), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_3), .B(n_151), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_4), .B(n_178), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_5), .B(n_178), .Y(n_509) );
INVx1_ASAP7_75t_L g147 ( .A(n_6), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_7), .B(n_178), .Y(n_538) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_9), .A2(n_463), .B1(n_758), .B2(n_762), .Y(n_757) );
NAND2xp33_ASAP7_75t_L g579 ( .A(n_10), .B(n_176), .Y(n_579) );
AND2x2_ASAP7_75t_L g181 ( .A(n_11), .B(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g192 ( .A(n_12), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g138 ( .A(n_13), .Y(n_138) );
AOI221x1_ASAP7_75t_L g484 ( .A1(n_14), .A2(n_26), .B1(n_151), .B2(n_159), .C(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_15), .B(n_178), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_16), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_17), .B(n_151), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_18), .A2(n_89), .B1(n_466), .B2(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_18), .Y(n_466) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_19), .A2(n_193), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_20), .B(n_136), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_21), .B(n_178), .Y(n_562) );
AO21x1_ASAP7_75t_L g504 ( .A1(n_22), .A2(n_151), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_23), .B(n_151), .Y(n_232) );
INVx1_ASAP7_75t_L g115 ( .A(n_24), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_25), .A2(n_93), .B1(n_142), .B2(n_151), .Y(n_141) );
NAND2x1_ASAP7_75t_L g496 ( .A(n_27), .B(n_178), .Y(n_496) );
NAND2x1_ASAP7_75t_L g537 ( .A(n_28), .B(n_176), .Y(n_537) );
OR2x2_ASAP7_75t_L g139 ( .A(n_29), .B(n_90), .Y(n_139) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_29), .A2(n_90), .B(n_138), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_30), .B(n_176), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_31), .B(n_178), .Y(n_578) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_32), .A2(n_182), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_33), .B(n_176), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_34), .A2(n_159), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_35), .B(n_178), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_36), .A2(n_159), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g149 ( .A(n_37), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g157 ( .A(n_37), .B(n_147), .Y(n_157) );
INVx1_ASAP7_75t_L g163 ( .A(n_37), .Y(n_163) );
OR2x6_ASAP7_75t_L g113 ( .A(n_38), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_39), .B(n_151), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_40), .A2(n_445), .B1(n_446), .B2(n_449), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_40), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_41), .B(n_151), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_42), .B(n_178), .Y(n_217) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_43), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_44), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_45), .B(n_176), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_46), .B(n_151), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_47), .A2(n_159), .B(n_174), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_48), .A2(n_63), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_48), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_49), .A2(n_159), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_50), .B(n_176), .Y(n_204) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_51), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_52), .B(n_176), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_53), .B(n_151), .Y(n_244) );
INVx1_ASAP7_75t_L g145 ( .A(n_54), .Y(n_145) );
INVx1_ASAP7_75t_L g154 ( .A(n_54), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_55), .B(n_178), .Y(n_177) );
INVxp33_ASAP7_75t_L g770 ( .A(n_56), .Y(n_770) );
AND2x2_ASAP7_75t_L g212 ( .A(n_57), .B(n_136), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_58), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_59), .B(n_178), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_60), .B(n_176), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_61), .A2(n_159), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_62), .B(n_151), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_63), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_64), .B(n_151), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_65), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_66), .A2(n_159), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g238 ( .A(n_67), .B(n_137), .Y(n_238) );
AO21x1_ASAP7_75t_L g506 ( .A1(n_68), .A2(n_159), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_69), .B(n_151), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_70), .B(n_176), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_71), .B(n_151), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_72), .B(n_176), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_73), .A2(n_97), .B1(n_159), .B2(n_161), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_74), .B(n_178), .Y(n_235) );
AND2x2_ASAP7_75t_L g520 ( .A(n_75), .B(n_137), .Y(n_520) );
INVx1_ASAP7_75t_L g150 ( .A(n_76), .Y(n_150) );
INVx1_ASAP7_75t_L g156 ( .A(n_76), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_77), .A2(n_123), .B1(n_451), .B2(n_452), .Y(n_122) );
INVxp33_ASAP7_75t_L g452 ( .A(n_77), .Y(n_452) );
AND2x2_ASAP7_75t_L g540 ( .A(n_77), .B(n_182), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_78), .B(n_176), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_79), .A2(n_159), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_80), .A2(n_159), .B(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_81), .A2(n_159), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g229 ( .A(n_82), .B(n_137), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_83), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g116 ( .A(n_84), .Y(n_116) );
AND2x2_ASAP7_75t_L g525 ( .A(n_85), .B(n_182), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_86), .B(n_151), .Y(n_564) );
AND2x2_ASAP7_75t_L g205 ( .A(n_87), .B(n_193), .Y(n_205) );
AND2x2_ASAP7_75t_L g505 ( .A(n_88), .B(n_219), .Y(n_505) );
INVx1_ASAP7_75t_L g467 ( .A(n_89), .Y(n_467) );
AND2x2_ASAP7_75t_L g499 ( .A(n_91), .B(n_182), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_92), .B(n_176), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_94), .B(n_178), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_95), .B(n_176), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_96), .A2(n_159), .B(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_98), .A2(n_159), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_99), .B(n_178), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_100), .B(n_178), .Y(n_530) );
BUFx2_ASAP7_75t_L g237 ( .A(n_101), .Y(n_237) );
OA22x2_ASAP7_75t_L g120 ( .A1(n_102), .A2(n_121), .B1(n_460), .B2(n_764), .Y(n_120) );
BUFx2_ASAP7_75t_L g768 ( .A(n_102), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_103), .A2(n_159), .B(n_577), .Y(n_576) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_120), .B(n_769), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_109), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_117), .Y(n_109) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g763 ( .A(n_111), .Y(n_763) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_112), .B(n_456), .Y(n_455) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_112), .B(n_113), .Y(n_472) );
OR2x6_ASAP7_75t_SL g475 ( .A(n_112), .B(n_456), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_113), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_453), .B(n_457), .Y(n_121) );
INVx2_ASAP7_75t_L g451 ( .A(n_123), .Y(n_451) );
AOI22x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_444), .B2(n_450), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_124), .A2(n_469), .B1(n_473), .B2(n_476), .Y(n_468) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_125), .A2(n_477), .B1(n_759), .B2(n_760), .Y(n_758) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_381), .Y(n_125) );
NAND3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_297), .C(n_334), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_265), .C(n_280), .Y(n_127) );
OAI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_209), .B1(n_239), .B2(n_251), .C(n_252), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_131), .B(n_194), .Y(n_130) );
OAI22xp33_ASAP7_75t_SL g325 ( .A1(n_131), .A2(n_289), .B1(n_326), .B2(n_329), .Y(n_325) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
OAI21xp33_ASAP7_75t_SL g335 ( .A1(n_132), .A2(n_336), .B(n_342), .Y(n_335) );
OR2x2_ASAP7_75t_L g364 ( .A(n_132), .B(n_196), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_132), .B(n_284), .Y(n_365) );
INVx2_ASAP7_75t_L g396 ( .A(n_132), .Y(n_396) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_133), .B(n_256), .Y(n_377) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g251 ( .A(n_134), .B(n_169), .Y(n_251) );
BUFx3_ASAP7_75t_L g277 ( .A(n_134), .Y(n_277) );
AND2x2_ASAP7_75t_L g413 ( .A(n_134), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g436 ( .A(n_134), .B(n_197), .Y(n_436) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
AND2x4_ASAP7_75t_L g208 ( .A(n_135), .B(n_140), .Y(n_208) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_136), .A2(n_141), .B(n_158), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_136), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_136), .A2(n_200), .B(n_201), .Y(n_199) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_136), .A2(n_484), .B(n_488), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_136), .A2(n_527), .B(n_528), .Y(n_526) );
OA21x2_ASAP7_75t_L g627 ( .A1(n_136), .A2(n_484), .B(n_488), .Y(n_627) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g219 ( .A(n_138), .B(n_139), .Y(n_219) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g160 ( .A(n_145), .B(n_147), .Y(n_160) );
AND2x4_ASAP7_75t_L g178 ( .A(n_145), .B(n_155), .Y(n_178) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x6_ASAP7_75t_L g159 ( .A(n_149), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
AND2x6_ASAP7_75t_L g176 ( .A(n_150), .B(n_153), .Y(n_176) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_157), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx5_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
AND2x4_ASAP7_75t_L g161 ( .A(n_160), .B(n_162), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_167), .B(n_197), .Y(n_356) );
INVx1_ASAP7_75t_L g393 ( .A(n_167), .Y(n_393) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_183), .Y(n_167) );
AND2x2_ASAP7_75t_L g207 ( .A(n_168), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g414 ( .A(n_168), .Y(n_414) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g257 ( .A(n_169), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_169), .B(n_183), .Y(n_258) );
AND2x2_ASAP7_75t_L g279 ( .A(n_169), .B(n_198), .Y(n_279) );
AND2x2_ASAP7_75t_L g361 ( .A(n_169), .B(n_184), .Y(n_361) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_172), .B(n_181), .Y(n_169) );
INVx4_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_180), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_177), .B(n_179), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_176), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_179), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_179), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_179), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_179), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_179), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_179), .A2(n_247), .B(n_248), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_179), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_179), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_179), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_179), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_179), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_179), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_179), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_179), .A2(n_578), .B(n_579), .Y(n_577) );
INVx3_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
AND2x4_ASAP7_75t_SL g254 ( .A(n_183), .B(n_198), .Y(n_254) );
INVx1_ASAP7_75t_L g285 ( .A(n_183), .Y(n_285) );
INVx2_ASAP7_75t_L g293 ( .A(n_183), .Y(n_293) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_183), .Y(n_317) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_184), .Y(n_206) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_192), .Y(n_184) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_185), .A2(n_534), .B(n_540), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_191), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_193), .A2(n_232), .B(n_233), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
AND2x2_ASAP7_75t_L g432 ( .A(n_195), .B(n_295), .Y(n_432) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g291 ( .A(n_197), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g343 ( .A(n_197), .B(n_258), .Y(n_343) );
AND2x2_ASAP7_75t_L g360 ( .A(n_197), .B(n_361), .Y(n_360) );
INVx4_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x4_ASAP7_75t_L g284 ( .A(n_198), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g300 ( .A(n_198), .Y(n_300) );
AND2x2_ASAP7_75t_L g344 ( .A(n_198), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g351 ( .A(n_198), .B(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_198), .B(n_257), .Y(n_366) );
BUFx2_ASAP7_75t_L g376 ( .A(n_198), .Y(n_376) );
AND2x2_ASAP7_75t_L g401 ( .A(n_198), .B(n_361), .Y(n_401) );
AND2x2_ASAP7_75t_L g422 ( .A(n_198), .B(n_423), .Y(n_422) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
INVx1_ASAP7_75t_L g353 ( .A(n_206), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_207), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g383 ( .A(n_207), .B(n_254), .Y(n_383) );
INVx3_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
AND2x2_ASAP7_75t_L g423 ( .A(n_208), .B(n_345), .Y(n_423) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_210), .A2(n_253), .B1(n_258), .B2(n_259), .Y(n_252) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_220), .Y(n_210) );
INVx4_ASAP7_75t_L g250 ( .A(n_211), .Y(n_250) );
INVx2_ASAP7_75t_L g287 ( .A(n_211), .Y(n_287) );
NAND2x1_ASAP7_75t_L g313 ( .A(n_211), .B(n_230), .Y(n_313) );
OR2x2_ASAP7_75t_L g328 ( .A(n_211), .B(n_263), .Y(n_328) );
OR2x2_ASAP7_75t_SL g355 ( .A(n_211), .B(n_327), .Y(n_355) );
AND2x2_ASAP7_75t_L g368 ( .A(n_211), .B(n_242), .Y(n_368) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_211), .Y(n_389) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_219), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_219), .A2(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_219), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_SL g558 ( .A(n_219), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_219), .A2(n_575), .B(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g268 ( .A(n_220), .Y(n_268) );
AND2x2_ASAP7_75t_L g400 ( .A(n_220), .B(n_374), .Y(n_400) );
NOR2x1_ASAP7_75t_SL g220 ( .A(n_221), .B(n_230), .Y(n_220) );
AND2x2_ASAP7_75t_L g241 ( .A(n_221), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g417 ( .A(n_221), .B(n_340), .Y(n_417) );
AO21x1_ASAP7_75t_SL g221 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_221) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_222), .A2(n_223), .B(n_229), .Y(n_264) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_222), .A2(n_493), .B(n_499), .Y(n_492) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_222), .A2(n_514), .B(n_520), .Y(n_513) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_222), .A2(n_514), .B(n_520), .Y(n_547) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_222), .A2(n_493), .B(n_499), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_228), .Y(n_223) );
OR2x2_ASAP7_75t_L g249 ( .A(n_230), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g260 ( .A(n_230), .B(n_250), .Y(n_260) );
AND2x2_ASAP7_75t_L g306 ( .A(n_230), .B(n_263), .Y(n_306) );
OR2x2_ASAP7_75t_L g327 ( .A(n_230), .B(n_242), .Y(n_327) );
INVx2_ASAP7_75t_SL g333 ( .A(n_230), .Y(n_333) );
AND2x2_ASAP7_75t_L g339 ( .A(n_230), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_230), .B(n_332), .Y(n_349) );
BUFx2_ASAP7_75t_L g371 ( .A(n_230), .Y(n_371) );
OR2x6_ASAP7_75t_L g230 ( .A(n_231), .B(n_238), .Y(n_230) );
INVx2_ASAP7_75t_L g418 ( .A(n_239), .Y(n_418) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
OR2x2_ASAP7_75t_L g443 ( .A(n_240), .B(n_287), .Y(n_443) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_241), .B(n_250), .Y(n_309) );
AND2x2_ASAP7_75t_L g380 ( .A(n_241), .B(n_260), .Y(n_380) );
INVx1_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_242), .Y(n_271) );
INVx1_ASAP7_75t_L g304 ( .A(n_242), .Y(n_304) );
INVx2_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_250), .B(n_271), .Y(n_270) );
BUFx2_ASAP7_75t_L g330 ( .A(n_250), .Y(n_330) );
INVx2_ASAP7_75t_SL g406 ( .A(n_251), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_253), .A2(n_308), .B1(n_310), .B2(n_314), .Y(n_307) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g434 ( .A(n_254), .B(n_290), .Y(n_434) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_256), .B(n_300), .Y(n_379) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g345 ( .A(n_257), .B(n_293), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_258), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g288 ( .A(n_259), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_259), .A2(n_403), .B1(n_407), .B2(n_409), .C(n_411), .Y(n_402) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g272 ( .A(n_260), .B(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_260), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_260), .B(n_303), .Y(n_358) );
INVx1_ASAP7_75t_SL g354 ( .A(n_261), .Y(n_354) );
AOI221xp5_ASAP7_75t_SL g382 ( .A1(n_261), .A2(n_272), .B1(n_383), .B2(n_384), .C(n_387), .Y(n_382) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_261), .A2(n_333), .A3(n_360), .B1(n_416), .B2(n_418), .C1(n_419), .C2(n_422), .Y(n_415) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
BUFx2_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_263), .Y(n_274) );
INVx2_ASAP7_75t_L g332 ( .A(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g373 ( .A(n_263), .B(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OA21x2_ASAP7_75t_SL g265 ( .A1(n_266), .A2(n_272), .B(n_275), .Y(n_265) );
AOI211xp5_ASAP7_75t_L g435 ( .A1(n_266), .A2(n_436), .B(n_437), .C(n_441), .Y(n_435) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
OR2x2_ASAP7_75t_L g324 ( .A(n_268), .B(n_286), .Y(n_324) );
OR2x2_ASAP7_75t_L g408 ( .A(n_268), .B(n_303), .Y(n_408) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g426 ( .A(n_273), .Y(n_426) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g281 ( .A(n_277), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g316 ( .A(n_279), .B(n_317), .Y(n_316) );
OAI322xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .A3(n_286), .B1(n_288), .B2(n_289), .C1(n_294), .C2(n_296), .Y(n_280) );
INVx1_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
OR2x2_ASAP7_75t_L g294 ( .A(n_283), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_283), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
OAI32xp33_ASAP7_75t_L g350 ( .A1(n_287), .A2(n_351), .A3(n_354), .B1(n_355), .B2(n_356), .Y(n_350) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g295 ( .A(n_290), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_290), .B(n_353), .Y(n_352) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_290), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g416 ( .A(n_290), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g337 ( .A(n_291), .Y(n_337) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_295), .B(n_361), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_318), .Y(n_297) );
OAI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_307), .Y(n_298) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g367 ( .A(n_306), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_309), .A2(n_329), .B1(n_431), .B2(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_311), .A2(n_358), .B(n_359), .C(n_362), .Y(n_357) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx3_ASAP7_75t_L g439 ( .A(n_313), .Y(n_439) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g320 ( .A(n_317), .Y(n_320) );
AO21x1_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_325), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g385 ( .A(n_320), .Y(n_385) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_326), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g341 ( .A(n_328), .Y(n_341) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NOR3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_357), .C(n_369), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_338), .A2(n_400), .B(n_401), .Y(n_399) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
O2A1O1Ixp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_344), .B(n_346), .C(n_350), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
INVx2_ASAP7_75t_L g427 ( .A(n_355), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g441 ( .A1(n_356), .A2(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g421 ( .A(n_361), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .A3(n_366), .B(n_367), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g440 ( .A(n_368), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_375), .B(n_378), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
BUFx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g390 ( .A(n_373), .Y(n_390) );
AOI21xp33_ASAP7_75t_SL g437 ( .A1(n_375), .A2(n_438), .B(n_440), .Y(n_437) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_376), .B(n_396), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_376), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g386 ( .A(n_377), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND5xp2_ASAP7_75t_L g381 ( .A(n_382), .B(n_402), .C(n_415), .D(n_424), .E(n_435), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_391), .B1(n_394), .B2(n_397), .C(n_399), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_428), .B(n_430), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g459 ( .A(n_455), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_457), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_757), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
CKINVDCx11_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
CKINVDCx6p67_ASAP7_75t_R g759 ( .A(n_470), .Y(n_759) );
INVx3_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_474), .Y(n_761) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND4xp75_ASAP7_75t_L g477 ( .A(n_478), .B(n_667), .C(n_707), .D(n_736), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_629), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_586), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_521), .B(n_541), .Y(n_480) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_482), .B(n_489), .Y(n_481) );
AND2x4_ASAP7_75t_L g585 ( .A(n_482), .B(n_546), .Y(n_585) );
INVx1_ASAP7_75t_SL g638 ( .A(n_482), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_482), .A2(n_674), .B(n_677), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_SL g677 ( .A1(n_482), .A2(n_678), .B(n_679), .C(n_680), .Y(n_677) );
NAND2x1_ASAP7_75t_L g718 ( .A(n_482), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_482), .B(n_679), .Y(n_740) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g544 ( .A(n_483), .Y(n_544) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_483), .Y(n_617) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_500), .Y(n_489) );
AND2x2_ASAP7_75t_L g609 ( .A(n_490), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g690 ( .A(n_490), .B(n_546), .Y(n_690) );
INVx1_ASAP7_75t_L g750 ( .A(n_490), .Y(n_750) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g594 ( .A(n_491), .B(n_512), .Y(n_594) );
AND2x2_ASAP7_75t_L g719 ( .A(n_491), .B(n_513), .Y(n_719) );
AND2x2_ASAP7_75t_L g724 ( .A(n_491), .B(n_684), .Y(n_724) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
BUFx3_ASAP7_75t_L g633 ( .A(n_492), .Y(n_633) );
AND2x2_ASAP7_75t_L g679 ( .A(n_492), .B(n_513), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
AND2x2_ASAP7_75t_L g664 ( .A(n_500), .B(n_543), .Y(n_664) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
AND2x4_ASAP7_75t_L g546 ( .A(n_501), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g656 ( .A(n_501), .B(n_640), .Y(n_656) );
AND2x2_ASAP7_75t_SL g699 ( .A(n_501), .B(n_627), .Y(n_699) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g635 ( .A(n_502), .Y(n_635) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g596 ( .A(n_503), .Y(n_596) );
OAI21x1_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g511 ( .A(n_505), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_512), .B(n_596), .Y(n_599) );
AND2x2_ASAP7_75t_L g684 ( .A(n_512), .B(n_627), .Y(n_684) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g681 ( .A(n_513), .B(n_544), .Y(n_681) );
AND2x2_ASAP7_75t_L g701 ( .A(n_513), .B(n_627), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_519), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_521), .B(n_590), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_521), .A2(n_713), .B1(n_714), .B2(n_715), .C(n_717), .Y(n_712) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI332xp33_ASAP7_75t_L g746 ( .A1(n_522), .A2(n_606), .A3(n_613), .B1(n_672), .B2(n_747), .B3(n_748), .C1(n_749), .C2(n_751), .Y(n_746) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
AND2x2_ASAP7_75t_L g552 ( .A(n_523), .B(n_533), .Y(n_552) );
AND2x2_ASAP7_75t_L g569 ( .A(n_523), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g581 ( .A(n_523), .Y(n_581) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_523), .B(n_582), .Y(n_641) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NOR2x1_ASAP7_75t_SL g603 ( .A(n_524), .B(n_570), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_524), .B(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g614 ( .A(n_524), .B(n_533), .Y(n_614) );
BUFx2_ASAP7_75t_L g649 ( .A(n_524), .Y(n_649) );
AND2x2_ASAP7_75t_L g704 ( .A(n_524), .B(n_573), .Y(n_704) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
OR2x2_ASAP7_75t_L g572 ( .A(n_532), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g582 ( .A(n_532), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g622 ( .A(n_532), .Y(n_622) );
AND2x2_ASAP7_75t_L g692 ( .A(n_532), .B(n_591), .Y(n_692) );
AND2x2_ASAP7_75t_L g705 ( .A(n_532), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_532), .B(n_706), .Y(n_723) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_533), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_548), .A3(n_553), .B1(n_567), .B2(n_584), .Y(n_541) );
INVx2_ASAP7_75t_L g650 ( .A(n_542), .Y(n_650) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g661 ( .A(n_543), .Y(n_661) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g595 ( .A(n_544), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g728 ( .A(n_544), .B(n_633), .Y(n_728) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g640 ( .A(n_547), .Y(n_640) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx2_ASAP7_75t_L g628 ( .A(n_550), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_550), .B(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_551), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g716 ( .A(n_551), .Y(n_716) );
AND2x2_ASAP7_75t_L g734 ( .A(n_551), .B(n_596), .Y(n_734) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp67_ASAP7_75t_SL g678 ( .A(n_554), .B(n_607), .Y(n_678) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_555), .B(n_589), .Y(n_676) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g752 ( .A(n_556), .B(n_622), .Y(n_752) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
INVx2_ASAP7_75t_L g624 ( .A(n_557), .Y(n_624) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_558), .B(n_566), .Y(n_565) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_580), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_568), .B(n_626), .Y(n_711) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND3x2_ASAP7_75t_L g666 ( .A(n_569), .B(n_613), .C(n_622), .Y(n_666) );
AND2x2_ASAP7_75t_L g590 ( .A(n_570), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_570), .B(n_573), .Y(n_647) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g601 ( .A(n_572), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g591 ( .A(n_573), .Y(n_591) );
INVx1_ASAP7_75t_L g606 ( .A(n_573), .Y(n_606) );
BUFx3_ASAP7_75t_L g613 ( .A(n_573), .Y(n_613) );
AND2x2_ASAP7_75t_L g623 ( .A(n_573), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x4_ASAP7_75t_L g632 ( .A(n_581), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_581), .B(n_591), .Y(n_675) );
AND2x2_ASAP7_75t_L g631 ( .A(n_582), .B(n_606), .Y(n_631) );
INVx2_ASAP7_75t_L g658 ( .A(n_582), .Y(n_658) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_592), .B(n_597), .C(n_618), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_587), .A2(n_714), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_590), .B(n_649), .Y(n_648) );
AOI211xp5_ASAP7_75t_SL g668 ( .A1(n_590), .A2(n_669), .B(n_673), .C(n_682), .Y(n_668) );
AND2x2_ASAP7_75t_L g654 ( .A(n_591), .B(n_614), .Y(n_654) );
OR2x2_ASAP7_75t_L g657 ( .A(n_591), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_594), .B(n_699), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_595), .B(n_640), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_595), .A2(n_621), .B1(n_701), .B2(n_704), .C(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g626 ( .A(n_596), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g672 ( .A(n_596), .B(n_627), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_601), .B1(n_604), .B2(n_608), .C(n_611), .Y(n_597) );
AND2x2_ASAP7_75t_L g743 ( .A(n_598), .B(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g610 ( .A(n_599), .Y(n_610) );
INVx1_ASAP7_75t_L g696 ( .A(n_600), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_601), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_603), .B(n_606), .Y(n_615) );
AND2x2_ASAP7_75t_L g691 ( .A(n_603), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g616 ( .A(n_610), .B(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_615), .B(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g735 ( .A(n_612), .Y(n_735) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g714 ( .A(n_613), .B(n_641), .Y(n_714) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_614), .B(n_623), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B(n_625), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_653), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g725 ( .A(n_619), .Y(n_725) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
INVx1_ASAP7_75t_L g706 ( .A(n_624), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_626), .B(n_696), .Y(n_747) );
AND2x2_ASAP7_75t_L g715 ( .A(n_627), .B(n_716), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_628), .A2(n_709), .B(n_712), .C(n_720), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_651), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .A3(n_634), .B1(n_636), .B2(n_641), .C1(n_642), .C2(n_650), .Y(n_630) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_632), .Y(n_748) );
AND2x2_ASAP7_75t_L g698 ( .A(n_633), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g732 ( .A(n_633), .Y(n_732) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_SL g683 ( .A(n_635), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_SL g689 ( .A(n_635), .B(n_681), .Y(n_689) );
AND2x2_ASAP7_75t_L g713 ( .A(n_635), .B(n_679), .Y(n_713) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g685 ( .A(n_639), .Y(n_685) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_SL g688 ( .A1(n_644), .A2(n_689), .B1(n_690), .B2(n_691), .C(n_693), .Y(n_688) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g755 ( .A(n_647), .Y(n_755) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_659), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g730 ( .A(n_654), .Y(n_730) );
INVx1_ASAP7_75t_L g662 ( .A(n_656), .Y(n_662) );
OR2x2_ASAP7_75t_L g749 ( .A(n_656), .B(n_750), .Y(n_749) );
INVx2_ASAP7_75t_SL g745 ( .A(n_657), .Y(n_745) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_665), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_661), .B(n_679), .Y(n_756) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_688), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_671), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OR2x2_ASAP7_75t_L g722 ( .A(n_675), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_686), .Y(n_682) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_697), .A3(n_700), .B(n_702), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_699), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_724), .B1(n_725), .B2(n_726), .C(n_729), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_746), .C(n_753), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_738), .B(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_745), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
BUFx4f_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
endmodule