module fake_jpeg_21790_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_48),
.B1(n_50),
.B2(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_26),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_56),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_55),
.Y(n_69)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_26),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_39),
.C(n_34),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_75),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_35),
.CI(n_34),
.CON(n_75),
.SN(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_82),
.B1(n_38),
.B2(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_17),
.B(n_36),
.C(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_101),
.B1(n_68),
.B2(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_98),
.Y(n_113)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.C(n_35),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_75),
.B1(n_77),
.B2(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_43),
.B1(n_35),
.B2(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_106),
.B1(n_21),
.B2(n_23),
.Y(n_131)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_108),
.Y(n_112)
);

AOI22x1_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_109),
.B1(n_81),
.B2(n_62),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_43),
.B1(n_58),
.B2(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_47),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_111),
.B(n_126),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_118),
.Y(n_148)
);

AO21x2_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_76),
.B(n_41),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_41),
.B(n_61),
.C(n_30),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_31),
.C(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_132),
.B(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_102),
.B1(n_93),
.B2(n_104),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_68),
.B1(n_81),
.B2(n_36),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_33),
.B1(n_36),
.B2(n_73),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_73),
.B1(n_60),
.B2(n_42),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_91),
.B1(n_99),
.B2(n_30),
.Y(n_146)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_29),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_29),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_99),
.B(n_10),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_60),
.B1(n_42),
.B2(n_25),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_78),
.B1(n_74),
.B2(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_138),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_153),
.B1(n_154),
.B2(n_115),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_105),
.B1(n_92),
.B2(n_96),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_127),
.B1(n_125),
.B2(n_118),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_120),
.B(n_112),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_155),
.B(n_157),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_91),
.B1(n_25),
.B2(n_95),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_152),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_149),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_131),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_41),
.B(n_30),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_149),
.B(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_114),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_164),
.B(n_165),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_180),
.B1(n_10),
.B2(n_13),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_116),
.C(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_148),
.C(n_136),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_128),
.B1(n_126),
.B2(n_119),
.Y(n_164)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_134),
.B(n_122),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_169),
.B(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_160),
.B(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_152),
.A2(n_132),
.B1(n_30),
.B2(n_24),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_179),
.B1(n_139),
.B2(n_156),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_1),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_24),
.B1(n_15),
.B2(n_2),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_24),
.B1(n_15),
.B2(n_2),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_185),
.Y(n_187)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_190),
.C(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_159),
.C(n_136),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_203),
.B1(n_172),
.B2(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_150),
.C(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_150),
.C(n_146),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_200),
.C(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_24),
.C(n_15),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_15),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_180),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_177),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_207),
.A2(n_179),
.B1(n_175),
.B2(n_164),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_3),
.C(n_5),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_204),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_170),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_217),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_189),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_177),
.B(n_182),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_178),
.B1(n_168),
.B2(n_184),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_225),
.B1(n_188),
.B2(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_223),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_184),
.B1(n_170),
.B2(n_183),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_166),
.B(n_181),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_186),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_232),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_230),
.A2(n_241),
.B1(n_244),
.B2(n_228),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_188),
.C(n_201),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_214),
.C(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_185),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_200),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_167),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_245),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_214),
.C(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_218),
.C(n_217),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_218),
.C(n_211),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.C(n_11),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_167),
.C(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_205),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_231),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_206),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_202),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_262),
.B(n_263),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_267),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_9),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_220),
.B1(n_207),
.B2(n_229),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_249),
.A2(n_173),
.B1(n_193),
.B2(n_199),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_176),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_270),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_11),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_246),
.B(n_11),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_260),
.B(n_271),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_14),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_13),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_9),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_12),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_288),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_265),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_273),
.B(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_279),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_14),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_285),
.B(n_289),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_295),
.C(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_292),
.C(n_278),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_286),
.B(n_14),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_7),
.B(n_8),
.Y(n_300)
);


endmodule