module real_jpeg_12511_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_2),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_3),
.A2(n_33),
.B1(n_68),
.B2(n_70),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_4),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_6),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_63),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_7),
.A2(n_56),
.B1(n_68),
.B2(n_70),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_68),
.B1(n_70),
.B2(n_87),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_37),
.B(n_38),
.C(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_13),
.A2(n_40),
.B1(n_68),
.B2(n_70),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_81),
.B1(n_85),
.B2(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_13),
.B(n_74),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_14),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_68),
.B1(n_70),
.B2(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_136)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_108),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_47),
.B1(n_48),
.B2(n_77),
.Y(n_21)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_24)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_25),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_25),
.A2(n_84),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_25),
.A2(n_30),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_26),
.A2(n_27),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_26),
.B(n_40),
.C(n_90),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_26),
.B(n_171),
.Y(n_170)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_30),
.B(n_136),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_32),
.A2(n_85),
.B(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_53)
);

OAI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_40),
.B(n_42),
.CON(n_133),
.SN(n_133)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_40),
.B(n_85),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_40),
.B(n_89),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_67),
.B2(n_71),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_41),
.B(n_68),
.C(n_71),
.Y(n_134)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_60),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_55),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_73),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_65),
.B1(n_74),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_64),
.A2(n_66),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_65),
.A2(n_74),
.B1(n_121),
.B2(n_133),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OA22x2_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_66)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_67),
.A2(n_70),
.B(n_132),
.C(n_134),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_70),
.B1(n_90),
.B2(n_92),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_70),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_99),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_88),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_81),
.A2(n_85),
.B1(n_165),
.B2(n_173),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_81),
.A2(n_167),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_93),
.B(n_94),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_SL g92 ( 
.A(n_90),
.Y(n_92)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_140),
.B1(n_142),
.B2(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_142),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_97),
.A2(n_142),
.B1(n_150),
.B2(n_160),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.C(n_105),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_113),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_109),
.B(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_111),
.B(n_113),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_119),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_119),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_196),
.B(n_200),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_151),
.B(n_195),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_146),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_143),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_137),
.C(n_143),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_135),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_141),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_149),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_190),
.B(n_194),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_179),
.B(n_189),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_168),
.B(n_178),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_163),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_161),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_177),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_185),
.C(n_188),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);


endmodule