module fake_jpeg_7982_n_263 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_17),
.Y(n_54)
);

AO21x1_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_17),
.B(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_32),
.B1(n_31),
.B2(n_37),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_71),
.B1(n_48),
.B2(n_42),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_30),
.B(n_36),
.C(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_53),
.B1(n_52),
.B2(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_28),
.B1(n_21),
.B2(n_17),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_28),
.B1(n_13),
.B2(n_26),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_45),
.C(n_42),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_90),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_81),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_94),
.B(n_22),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_94),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_50),
.B1(n_49),
.B2(n_46),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_33),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_41),
.B1(n_43),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_71),
.B1(n_82),
.B2(n_84),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_23),
.B(n_20),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_107),
.B1(n_79),
.B2(n_92),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_70),
.B1(n_41),
.B2(n_39),
.Y(n_97)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_76),
.B1(n_91),
.B2(n_56),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_77),
.A2(n_65),
.B(n_15),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_112),
.B(n_14),
.Y(n_117)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_111),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_109),
.B1(n_74),
.B2(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_74),
.B1(n_66),
.B2(n_65),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_110),
.B1(n_69),
.B2(n_38),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_66),
.B1(n_73),
.B2(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_15),
.B(n_22),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_21),
.B(n_14),
.C(n_19),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_19),
.B(n_12),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_83),
.B(n_80),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_123),
.B(n_97),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_129),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_90),
.B1(n_82),
.B2(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_126),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_75),
.B(n_76),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_130),
.B1(n_97),
.B2(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_12),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_127),
.B(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_93),
.B1(n_74),
.B2(n_23),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_35),
.C(n_56),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_110),
.C(n_108),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_69),
.B1(n_38),
.B2(n_16),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_137),
.B1(n_26),
.B2(n_24),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_105),
.B1(n_103),
.B2(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_27),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_69),
.B1(n_38),
.B2(n_16),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_109),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_139),
.C(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_155),
.B1(n_131),
.B2(n_120),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_145),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_148),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_35),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_153),
.C(n_156),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_158),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_26),
.Y(n_156)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_24),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_24),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_122),
.C(n_118),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_135),
.B1(n_126),
.B2(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_116),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_117),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_139),
.C(n_151),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_124),
.B(n_128),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_1),
.B(n_2),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_18),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_18),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_180),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_145),
.B(n_18),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_164),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_198),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_SL g188 ( 
.A(n_167),
.B(n_147),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_153),
.C(n_143),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_152),
.C(n_1),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_0),
.C(n_1),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_1),
.C(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_2),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_175),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_204),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_188),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_3),
.C(n_5),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_189),
.B1(n_168),
.B2(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_178),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_214),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_180),
.B1(n_169),
.B2(n_170),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_2),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_195),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_219),
.C(n_202),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_194),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_193),
.B1(n_4),
.B2(n_5),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_199),
.B1(n_8),
.B2(n_9),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_3),
.B(n_5),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_3),
.B(n_6),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_227),
.B1(n_212),
.B2(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_204),
.B(n_202),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_7),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.C(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_218),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_7),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_7),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_244),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_7),
.B(n_8),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_250),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_229),
.B1(n_237),
.B2(n_232),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_229),
.B1(n_236),
.B2(n_10),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_8),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_239),
.B1(n_10),
.B2(n_11),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

AOI21x1_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_9),
.B(n_11),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_254),
.B(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_254),
.C(n_255),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_256),
.B(n_258),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_247),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_9),
.B(n_11),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_11),
.Y(n_263)
);


endmodule