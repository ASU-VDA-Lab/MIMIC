module fake_jpeg_3702_n_481 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_481);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_481;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_16),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_57),
.Y(n_151)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_70),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_60),
.B(n_67),
.Y(n_123)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_61),
.Y(n_163)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_62),
.Y(n_184)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_63),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_87),
.Y(n_132)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_84),
.B(n_93),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_85),
.Y(n_130)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_86),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_89),
.Y(n_157)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_25),
.B(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_98),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_14),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_100),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_22),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_103),
.Y(n_190)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_102),
.B(n_104),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_12),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_22),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_108),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_22),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_36),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_110),
.Y(n_174)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_112),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_36),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_113),
.B(n_116),
.Y(n_191)
);

BUFx4f_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_114),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_52),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_117),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_36),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g118 ( 
.A(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_41),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_33),
.B1(n_49),
.B2(n_47),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_121),
.A2(n_124),
.B1(n_153),
.B2(n_154),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_48),
.B1(n_38),
.B2(n_31),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_51),
.B1(n_50),
.B2(n_41),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_125),
.A2(n_129),
.B1(n_138),
.B2(n_143),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_115),
.B1(n_119),
.B2(n_117),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_38),
.B1(n_50),
.B2(n_51),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_133),
.A2(n_152),
.B1(n_167),
.B2(n_137),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_46),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_137),
.B(n_150),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_62),
.A2(n_46),
.B1(n_38),
.B2(n_49),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_63),
.A2(n_48),
.B1(n_30),
.B2(n_23),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_139),
.A2(n_171),
.B1(n_156),
.B2(n_133),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_64),
.A2(n_47),
.B1(n_20),
.B2(n_33),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_32),
.B1(n_20),
.B2(n_30),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_147),
.A2(n_149),
.B1(n_194),
.B2(n_115),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_32),
.B1(n_30),
.B2(n_23),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_24),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_79),
.A2(n_24),
.B1(n_30),
.B2(n_23),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_152),
.B(n_167),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_69),
.A2(n_30),
.B1(n_23),
.B2(n_35),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_73),
.A2(n_35),
.B1(n_18),
.B2(n_2),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_83),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_155),
.A2(n_160),
.B1(n_164),
.B2(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_65),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_158),
.B(n_151),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_0),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_159),
.B(n_170),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_111),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_96),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_92),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_168),
.A2(n_94),
.B(n_195),
.C(n_193),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_72),
.A2(n_80),
.B1(n_104),
.B2(n_89),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_176),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_74),
.A2(n_8),
.B1(n_9),
.B2(n_107),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_118),
.A2(n_92),
.B1(n_88),
.B2(n_110),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_192),
.B1(n_151),
.B2(n_180),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_57),
.B1(n_77),
.B2(n_78),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_77),
.A2(n_29),
.B1(n_26),
.B2(n_55),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_78),
.C(n_94),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_197),
.B(n_217),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_120),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_198),
.B(n_218),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_201),
.A2(n_206),
.B1(n_224),
.B2(n_249),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_202),
.Y(n_306)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_195),
.B(n_168),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_208),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_209),
.B(n_210),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_141),
.B(n_165),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_211),
.B(n_212),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_123),
.B(n_132),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_150),
.A2(n_174),
.B(n_171),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_213),
.B(n_221),
.Y(n_292)
);

BUFx4f_ASAP7_75t_SL g214 ( 
.A(n_127),
.Y(n_214)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_159),
.A2(n_139),
.B1(n_134),
.B2(n_185),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_215),
.A2(n_217),
.B1(n_227),
.B2(n_244),
.Y(n_302)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_186),
.A2(n_185),
.B1(n_184),
.B2(n_163),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_145),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_127),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_223),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_248),
.Y(n_277)
);

OR2x2_ASAP7_75t_SL g221 ( 
.A(n_157),
.B(n_181),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_131),
.B(n_181),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_162),
.A2(n_183),
.B1(n_182),
.B2(n_163),
.Y(n_224)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_148),
.A2(n_184),
.B1(n_162),
.B2(n_170),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_230),
.B(n_234),
.Y(n_291)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_231),
.Y(n_276)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_235),
.B(n_236),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_240),
.Y(n_294)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_239),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_189),
.B(n_187),
.Y(n_240)
);

INVx6_ASAP7_75t_SL g241 ( 
.A(n_180),
.Y(n_241)
);

INVx2_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

BUFx16f_ASAP7_75t_L g242 ( 
.A(n_126),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_242),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_243),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_161),
.A2(n_172),
.B1(n_135),
.B2(n_173),
.Y(n_244)
);

BUFx6f_ASAP7_75t_SL g245 ( 
.A(n_140),
.Y(n_245)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_131),
.B(n_157),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_247),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_142),
.B(n_135),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_172),
.A2(n_177),
.B1(n_140),
.B2(n_128),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_252),
.Y(n_293)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_254),
.Y(n_301)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_224),
.B1(n_245),
.B2(n_222),
.Y(n_280)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_257),
.Y(n_303)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_121),
.A2(n_137),
.B1(n_150),
.B2(n_133),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_213),
.B1(n_260),
.B2(n_206),
.Y(n_271)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_144),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_261),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_131),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_262),
.A2(n_272),
.B(n_292),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_269),
.B(n_272),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_271),
.A2(n_305),
.B1(n_302),
.B2(n_270),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_199),
.B(n_221),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_229),
.A2(n_201),
.B1(n_225),
.B2(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_275),
.A2(n_234),
.B1(n_243),
.B2(n_266),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_280),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g282 ( 
.A(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_284),
.Y(n_313)
);

AOI32xp33_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_200),
.A3(n_233),
.B1(n_255),
.B2(n_241),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_234),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_197),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_296),
.B(n_309),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_307),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_200),
.A2(n_231),
.B1(n_202),
.B2(n_237),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_226),
.B(n_257),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_214),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_275),
.A2(n_271),
.B1(n_266),
.B2(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_311),
.A2(n_329),
.B1(n_346),
.B2(n_270),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_269),
.B(n_207),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_312),
.B(n_315),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_204),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_322),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_214),
.B(n_216),
.C(n_256),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_263),
.B(n_340),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_336),
.C(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_320),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_321),
.A2(n_339),
.B1(n_341),
.B2(n_343),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_243),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_323),
.A2(n_335),
.B(n_340),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_278),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_327),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_293),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_284),
.A2(n_285),
.B(n_296),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_328),
.A2(n_313),
.B(n_326),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_297),
.A2(n_295),
.B1(n_277),
.B2(n_299),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_279),
.Y(n_330)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_290),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_333),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_301),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_264),
.C(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_265),
.Y(n_338)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_309),
.B(n_308),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_267),
.B(n_303),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_342),
.A2(n_345),
.B(n_276),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_286),
.B(n_288),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_288),
.B(n_277),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_273),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_267),
.B(n_287),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_349),
.B(n_363),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_273),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_357),
.C(n_360),
.Y(n_388)
);

OAI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_356),
.A2(n_353),
.B1(n_366),
.B2(n_348),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_287),
.Y(n_357)
);

A2O1A1O1Ixp25_ASAP7_75t_L g358 ( 
.A1(n_313),
.A2(n_283),
.B(n_263),
.C(n_274),
.D(n_304),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_358),
.A2(n_371),
.B(n_314),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_283),
.C(n_300),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_315),
.C(n_324),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_321),
.A2(n_276),
.B1(n_289),
.B2(n_300),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_362),
.A2(n_366),
.B1(n_367),
.B2(n_373),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_311),
.A2(n_289),
.B1(n_306),
.B2(n_310),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_346),
.A2(n_306),
.B1(n_310),
.B2(n_274),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_340),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_328),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_336),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_333),
.A2(n_316),
.B1(n_326),
.B2(n_329),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_334),
.Y(n_375)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_347),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_374),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g400 ( 
.A(n_378),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_380),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_356),
.A2(n_318),
.B1(n_334),
.B2(n_319),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_373),
.A2(n_318),
.B1(n_327),
.B2(n_340),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_385),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_369),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_384),
.Y(n_414)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_387),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_339),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_389),
.B(n_396),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_399),
.C(n_388),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_353),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_393),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_392),
.B(n_368),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_342),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_335),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_394),
.B(n_397),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_395),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_371),
.A2(n_322),
.B1(n_332),
.B2(n_325),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_350),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_398),
.B(n_399),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_312),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_399),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_388),
.B(n_360),
.C(n_361),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_405),
.C(n_406),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_354),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_354),
.C(n_348),
.Y(n_406)
);

OAI322xp33_ASAP7_75t_L g407 ( 
.A1(n_391),
.A2(n_350),
.A3(n_374),
.B1(n_372),
.B2(n_343),
.C1(n_358),
.C2(n_344),
.Y(n_407)
);

AOI321xp33_ASAP7_75t_L g435 ( 
.A1(n_407),
.A2(n_395),
.A3(n_387),
.B1(n_317),
.B2(n_393),
.C(n_385),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_349),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_417),
.C(n_376),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_SL g418 ( 
.A(n_394),
.B(n_375),
.C(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_418),
.B(n_420),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_410),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_433),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_397),
.Y(n_423)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_412),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_428),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_429),
.C(n_431),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_386),
.Y(n_447)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_402),
.C(n_405),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_383),
.C(n_396),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_401),
.A2(n_398),
.B(n_384),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_432),
.A2(n_414),
.B(n_380),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_L g433 ( 
.A1(n_406),
.A2(n_376),
.B(n_381),
.Y(n_433)
);

AO221x1_ASAP7_75t_L g434 ( 
.A1(n_418),
.A2(n_367),
.B1(n_362),
.B2(n_389),
.C(n_317),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_434),
.A2(n_435),
.B1(n_380),
.B2(n_411),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_416),
.A2(n_408),
.B1(n_415),
.B2(n_411),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_436),
.A2(n_408),
.B1(n_379),
.B2(n_403),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_432),
.A2(n_395),
.B(n_415),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_439),
.A2(n_446),
.B(n_436),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_417),
.C(n_420),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_442),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_445),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_412),
.B1(n_379),
.B2(n_409),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_447),
.B(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_452),
.Y(n_459)
);

AOI321xp33_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_435),
.A3(n_430),
.B1(n_428),
.B2(n_431),
.C(n_423),
.Y(n_450)
);

INVx11_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_438),
.B(n_400),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_438),
.B(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_454),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_422),
.C(n_426),
.Y(n_454)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_455),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_437),
.A2(n_424),
.B1(n_414),
.B2(n_382),
.Y(n_456)
);

MAJx2_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_443),
.C(n_444),
.Y(n_462)
);

OA21x2_ASAP7_75t_SL g457 ( 
.A1(n_440),
.A2(n_414),
.B(n_345),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_457),
.B(n_439),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_461),
.B(n_462),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_454),
.B(n_445),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_465),
.B(n_466),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_458),
.B(n_451),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_464),
.A2(n_455),
.B1(n_456),
.B2(n_443),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_441),
.B(n_446),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_470),
.A2(n_471),
.B1(n_463),
.B2(n_459),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g471 ( 
.A(n_462),
.B(n_450),
.CI(n_451),
.CON(n_471),
.SN(n_471)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_472),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_468),
.A2(n_463),
.B(n_424),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_467),
.B(n_471),
.C(n_414),
.Y(n_476)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_469),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_468),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_475),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g479 ( 
.A(n_476),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_478),
.B(n_477),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_480),
.B(n_479),
.Y(n_481)
);


endmodule