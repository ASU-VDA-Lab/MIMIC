module real_jpeg_4073_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_86),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_189),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_1),
.A2(n_189),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_1),
.A2(n_189),
.B1(n_213),
.B2(n_215),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_38),
.B1(n_61),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_46),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_3),
.A2(n_46),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_5),
.A2(n_85),
.B1(n_86),
.B2(n_90),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_5),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_85),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_5),
.A2(n_85),
.B1(n_165),
.B2(n_335),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_5),
.A2(n_47),
.B1(n_85),
.B2(n_158),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_6),
.A2(n_246),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_6),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_6),
.A2(n_273),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_6),
.A2(n_273),
.B1(n_342),
.B2(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_6),
.A2(n_86),
.B1(n_273),
.B2(n_431),
.Y(n_430)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_8),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_9),
.A2(n_231),
.B1(n_234),
.B2(n_237),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_9),
.B(n_248),
.C(n_252),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_9),
.B(n_133),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_9),
.B(n_170),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_9),
.B(n_79),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_9),
.B(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_12),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_13),
.A2(n_74),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_13),
.A2(n_74),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_14),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_14),
.A2(n_50),
.B1(n_146),
.B2(n_173),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_14),
.A2(n_146),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_14),
.A2(n_146),
.B1(n_262),
.B2(n_368),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_16),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_16),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_16),
.A2(n_104),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_16),
.A2(n_104),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_16),
.A2(n_104),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_221),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_219),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_191),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_20),
.B(n_191),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_116),
.C(n_161),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_21),
.A2(n_22),
.B1(n_116),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_23),
.A2(n_24),
.B(n_82),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_24),
.A2(n_81),
.B1(n_82),
.B2(n_115),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_24),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_24),
.A2(n_44),
.B1(n_115),
.B2(n_420),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_35),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_25),
.A2(n_37),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_257),
.B(n_263),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_25),
.A2(n_237),
.B(n_263),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_25),
.A2(n_390),
.B1(n_391),
.B2(n_392),
.Y(n_389)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_26),
.B(n_266),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_26),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_26),
.A2(n_334),
.B1(n_367),
.B2(n_370),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_26),
.A2(n_393),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_33),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_35),
.A2(n_290),
.B(n_294),
.Y(n_289)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_35),
.Y(n_370)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_40),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_43),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_44),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_53),
.B1(n_73),
.B2(n_79),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_45),
.A2(n_53),
.B1(n_79),
.B2(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_48),
.Y(n_276)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_49),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_51),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_53),
.A2(n_73),
.B1(n_79),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_53),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_53),
.B(n_239),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_55),
.Y(n_173)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_58),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_63),
.A2(n_272),
.B(n_277),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_69),
.Y(n_165)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_69),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_69),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_69),
.Y(n_336)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_70),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_71),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_71),
.Y(n_398)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_75),
.Y(n_343)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_76),
.Y(n_240)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_79),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_79),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_102),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_84),
.Y(n_197)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_92),
.B(n_103),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_93),
.B(n_237),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_93),
.A2(n_184),
.B1(n_185),
.B2(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_93)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_94),
.Y(n_386)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_97),
.Y(n_329)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_98),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_98),
.Y(n_216)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_100),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_102),
.A2(n_198),
.B(n_430),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_107),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_107),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_110),
.Y(n_384)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_116),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_154),
.B(n_160),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_155),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_133),
.B1(n_139),
.B2(n_147),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_119),
.A2(n_322),
.B(n_326),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_119),
.B(n_363),
.Y(n_362)
);

AOI22x1_ASAP7_75t_L g433 ( 
.A1(n_119),
.A2(n_133),
.B1(n_363),
.B2(n_434),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_119),
.A2(n_326),
.B(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_140),
.B1(n_175),
.B2(n_182),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_120),
.A2(n_182),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_120),
.A2(n_182),
.B1(n_359),
.B2(n_409),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_133),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_126),
.Y(n_325)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_132),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_133),
.Y(n_182)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_135),
.Y(n_345)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_137),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_144),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_148),
.A2(n_380),
.A3(n_384),
.B1(n_385),
.B2(n_387),
.Y(n_379)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_161),
.B(n_436),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_174),
.C(n_183),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_162),
.B(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_171),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_163),
.B(n_171),
.Y(n_444)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_164),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_170),
.Y(n_427)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_172),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_174),
.B(n_183),
.Y(n_418)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_175),
.Y(n_434)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_182),
.B(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_182),
.A2(n_359),
.B(n_362),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B(n_190),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_187),
.B(n_237),
.Y(n_387)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_188),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_190),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_205),
.B2(n_218),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_217),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_207),
.A2(n_230),
.B(n_238),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_207),
.A2(n_208),
.B1(n_272),
.B2(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_207),
.A2(n_238),
.B(n_315),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_207),
.A2(n_208),
.B1(n_411),
.B2(n_424),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_208),
.A2(n_277),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_SL g322 ( 
.A1(n_215),
.A2(n_237),
.B(n_323),
.Y(n_322)
);

INVx6_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI311xp33_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_414),
.A3(n_452),
.B1(n_470),
.C1(n_471),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_373),
.B(n_413),
.Y(n_223)
);

AO21x1_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_350),
.B(n_372),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_309),
.B(n_349),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_280),
.B(n_308),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_255),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_243),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_229),
.A2(n_243),
.B1(n_244),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g405 ( 
.A1(n_237),
.A2(n_381),
.B(n_387),
.Y(n_405)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_269),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_270),
.C(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_264),
.Y(n_391)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_267),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_278),
.B2(n_279),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_297),
.B(n_307),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_288),
.B(n_296),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_295),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_295),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_291),
.Y(n_369)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_294),
.A2(n_333),
.B(n_337),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_305),
.Y(n_307)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_311),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_331),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_320),
.B2(n_321),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_320),
.C(n_331),
.Y(n_351)
);

INVx3_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_341),
.A3(n_343),
.B1(n_344),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_328),
.B(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_345),
.B(n_347),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_351),
.B(n_352),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_357),
.B2(n_371),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_356),
.C(n_371),
.Y(n_374)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_364),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_365),
.C(n_366),
.Y(n_399)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_374),
.B(n_375),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_402),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_399),
.B1(n_400),
.B2(n_401),
.Y(n_376)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_379),
.B1(n_388),
.B2(n_389),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_379),
.B(n_388),
.Y(n_448)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_399),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_400),
.C(n_402),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_407),
.B2(n_412),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_408),
.C(n_410),
.Y(n_461)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_407),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_438),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_SL g471 ( 
.A1(n_415),
.A2(n_438),
.B(n_472),
.C(n_475),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_435),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_435),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.C(n_421),
.Y(n_416)
);

FAx1_ASAP7_75t_SL g451 ( 
.A(n_417),
.B(n_419),
.CI(n_421),
.CON(n_451),
.SN(n_451)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_428),
.C(n_433),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_425),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_428),
.A2(n_429),
.B1(n_433),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_433),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_451),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_451),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_444),
.C(n_445),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_440),
.A2(n_441),
.B1(n_444),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_463),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.C(n_449),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_446),
.A2(n_447),
.B1(n_449),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_451),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_465),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_454),
.A2(n_473),
.B(n_474),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_462),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_462),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.C(n_461),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_468),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_460),
.B1(n_461),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_461),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_467),
.Y(n_473)
);


endmodule