module fake_jpeg_13175_n_554 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_554);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_554;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_9),
.B(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_54),
.B(n_67),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_56),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_16),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_73),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_1),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_78),
.Y(n_171)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_23),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_82),
.A2(n_39),
.B1(n_28),
.B2(n_36),
.Y(n_163)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_93),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_1),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_25),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_100),
.Y(n_109)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_27),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_102),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_16),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g103 ( 
.A(n_48),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_103),
.Y(n_146)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_44),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_33),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_131),
.B(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_82),
.B(n_33),
.C(n_50),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_58),
.A2(n_23),
.B1(n_42),
.B2(n_40),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_153),
.Y(n_204)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_155),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_66),
.B(n_39),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_65),
.B(n_51),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_38),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_203)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_147),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_173),
.B(n_192),
.C(n_139),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_108),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_175),
.B(n_178),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_176),
.A2(n_196),
.B1(n_222),
.B2(n_226),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_64),
.B1(n_75),
.B2(n_24),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_179),
.B(n_95),
.Y(n_250)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_122),
.A2(n_24),
.B1(n_51),
.B2(n_50),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_119),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_110),
.B(n_45),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_202),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_106),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_109),
.B(n_49),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_193),
.B(n_194),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_128),
.B(n_49),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_63),
.B1(n_87),
.B2(n_80),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_138),
.B(n_124),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_230),
.B1(n_137),
.B2(n_133),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_113),
.A2(n_31),
.B1(n_45),
.B2(n_29),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_206),
.Y(n_280)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g270 ( 
.A(n_210),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_128),
.B(n_49),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_211),
.B(n_215),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_158),
.A2(n_29),
.B1(n_31),
.B2(n_79),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_213),
.A2(n_228),
.B1(n_231),
.B2(n_170),
.Y(n_260)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_146),
.B(n_37),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_149),
.B(n_21),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_221),
.B(n_223),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_161),
.A2(n_72),
.B1(n_62),
.B2(n_77),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_151),
.B(n_20),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_133),
.B(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_4),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_171),
.A2(n_74),
.B1(n_71),
.B2(n_94),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_119),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_229),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_142),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_111),
.A2(n_105),
.B1(n_19),
.B2(n_44),
.Y(n_230)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_142),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_116),
.A2(n_88),
.B1(n_95),
.B2(n_44),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_92),
.B(n_20),
.Y(n_237)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_26),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_236),
.A2(n_261),
.B1(n_262),
.B2(n_266),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_120),
.B1(n_125),
.B2(n_150),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_274),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_173),
.B(n_132),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_242),
.B(n_253),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_246),
.B(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_267),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_202),
.B(n_88),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_252),
.B(n_275),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_260),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_174),
.A2(n_136),
.B1(n_118),
.B2(n_162),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_195),
.A2(n_136),
.B1(n_118),
.B2(n_162),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_191),
.A2(n_170),
.B1(n_115),
.B2(n_92),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_207),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_273),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_173),
.B(n_26),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_242),
.C(n_264),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_180),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_225),
.B(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_189),
.B(n_26),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_26),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_277),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_192),
.B(n_21),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_208),
.B(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_285),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_190),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_13),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_21),
.B(n_20),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_284),
.A2(n_224),
.B(n_186),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_5),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_246),
.Y(n_327)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_226),
.B1(n_210),
.B2(n_231),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_290),
.A2(n_270),
.B1(n_241),
.B2(n_258),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_235),
.A2(n_214),
.B1(n_216),
.B2(n_233),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_293),
.B(n_331),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_245),
.A2(n_182),
.B1(n_197),
.B2(n_229),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_295),
.A2(n_299),
.B1(n_301),
.B2(n_306),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_182),
.B1(n_187),
.B2(n_185),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_296),
.A2(n_325),
.B1(n_241),
.B2(n_257),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_249),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_298),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_245),
.A2(n_228),
.B1(n_181),
.B2(n_219),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_253),
.A2(n_199),
.B1(n_201),
.B2(n_187),
.Y(n_301)
);

OAI22x1_ASAP7_75t_L g302 ( 
.A1(n_235),
.A2(n_200),
.B1(n_172),
.B2(n_217),
.Y(n_302)
);

OAI21xp33_ASAP7_75t_SL g350 ( 
.A1(n_302),
.A2(n_238),
.B(n_268),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_265),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_321),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_259),
.A2(n_185),
.B1(n_205),
.B2(n_204),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_212),
.C(n_172),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_307),
.B(n_318),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_309),
.A2(n_268),
.B(n_238),
.Y(n_348)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_311),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_280),
.A2(n_198),
.B1(n_184),
.B2(n_200),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_259),
.A2(n_212),
.B(n_218),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_317),
.A2(n_243),
.B(n_248),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_21),
.C(n_7),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_6),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_319),
.B(n_285),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_243),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_334),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_273),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_256),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_324),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_262),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_330),
.Y(n_373)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_280),
.A2(n_7),
.B(n_10),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_284),
.B(n_237),
.Y(n_338)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_7),
.C(n_10),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_274),
.B(n_10),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_333),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_239),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_279),
.B1(n_241),
.B2(n_255),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_338),
.A2(n_341),
.B(n_344),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_346),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_309),
.A2(n_281),
.B(n_250),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_343),
.B(n_332),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_329),
.A2(n_252),
.B(n_267),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_345),
.A2(n_352),
.B1(n_356),
.B2(n_367),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_348),
.A2(n_355),
.B(n_360),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_364),
.B1(n_320),
.B2(n_335),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_299),
.A2(n_239),
.B1(n_255),
.B2(n_258),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_323),
.A2(n_239),
.B(n_254),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_315),
.A2(n_254),
.B(n_248),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_361),
.A2(n_368),
.B(n_374),
.Y(n_402)
);

OAI32xp33_ASAP7_75t_L g363 ( 
.A1(n_315),
.A2(n_278),
.A3(n_263),
.B1(n_286),
.B2(n_240),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_365),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_313),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_295),
.A2(n_257),
.B1(n_263),
.B2(n_286),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_317),
.A2(n_14),
.B(n_15),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_240),
.B1(n_15),
.B2(n_16),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_372),
.A2(n_378),
.B1(n_325),
.B2(n_294),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_297),
.A2(n_15),
.B1(n_305),
.B2(n_322),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_306),
.B(n_301),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_377),
.A2(n_328),
.B(n_355),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_297),
.A2(n_333),
.B1(n_294),
.B2(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_381),
.A2(n_386),
.B1(n_390),
.B2(n_407),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_288),
.C(n_293),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_382),
.B(n_389),
.C(n_393),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_349),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_383),
.B(n_387),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_384),
.A2(n_399),
.B1(n_346),
.B2(n_365),
.Y(n_416)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_351),
.Y(n_385)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_378),
.A2(n_312),
.B1(n_296),
.B2(n_316),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_349),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_288),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_342),
.A2(n_312),
.B1(n_316),
.B2(n_327),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_400),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_307),
.C(n_308),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_298),
.C(n_318),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_403),
.C(n_404),
.Y(n_429)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_337),
.B(n_300),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_398),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_337),
.B(n_331),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_289),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_304),
.C(n_310),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_342),
.A2(n_326),
.B1(n_336),
.B2(n_311),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_410),
.Y(n_442)
);

OAI32xp33_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_334),
.A3(n_302),
.B1(n_303),
.B2(n_330),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_302),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_377),
.C(n_338),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_340),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_414),
.Y(n_445)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_415),
.A2(n_361),
.B(n_368),
.Y(n_420)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_416),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_369),
.B1(n_352),
.B2(n_345),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_417),
.A2(n_386),
.B1(n_381),
.B2(n_407),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_388),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_447),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_420),
.A2(n_410),
.B(n_373),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_347),
.C(n_360),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_402),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_384),
.A2(n_374),
.B1(n_354),
.B2(n_371),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_389),
.B(n_341),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_432),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_403),
.B(n_371),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_426),
.B(n_424),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_354),
.B1(n_339),
.B2(n_379),
.Y(n_427)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_405),
.A2(n_353),
.B1(n_343),
.B2(n_344),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_377),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_437),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_415),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_439),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_408),
.A2(n_368),
.B(n_350),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_436),
.A2(n_340),
.B(n_375),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_363),
.Y(n_437)
);

OAI22x1_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_377),
.B1(n_367),
.B2(n_372),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_392),
.A2(n_373),
.B1(n_377),
.B2(n_375),
.Y(n_441)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_441),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_395),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_449),
.A2(n_463),
.B1(n_464),
.B2(n_448),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_423),
.A2(n_406),
.B1(n_390),
.B2(n_402),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_450),
.A2(n_420),
.B1(n_442),
.B2(n_432),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_393),
.C(n_406),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_456),
.B(n_457),
.C(n_460),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_411),
.C(n_414),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_458),
.B(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_385),
.C(n_409),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_380),
.C(n_400),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_474),
.C(n_421),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_364),
.B1(n_413),
.B2(n_391),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_467),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_434),
.A2(n_340),
.B(n_375),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_436),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_445),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_469),
.B(n_472),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_438),
.B(n_362),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_473),
.B(n_423),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_362),
.C(n_433),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_475),
.A2(n_471),
.B1(n_476),
.B2(n_479),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_453),
.A2(n_442),
.B1(n_435),
.B2(n_431),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g509 ( 
.A(n_476),
.B(n_455),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_444),
.B1(n_431),
.B2(n_439),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_479),
.A2(n_487),
.B1(n_493),
.B2(n_467),
.Y(n_511)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_482),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_492),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_468),
.Y(n_485)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_454),
.Y(n_486)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_452),
.A2(n_440),
.B1(n_425),
.B2(n_443),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_490),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_489),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_426),
.C(n_447),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_461),
.B(n_446),
.C(n_440),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_491),
.B(n_495),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_446),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_464),
.A2(n_425),
.B1(n_443),
.B2(n_459),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_449),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_466),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_457),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_456),
.C(n_474),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_505),
.B(n_512),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_485),
.A2(n_450),
.B1(n_462),
.B2(n_458),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_475),
.B(n_462),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_509),
.Y(n_525)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_508),
.Y(n_514)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_511),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_455),
.C(n_451),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_513),
.A2(n_490),
.B1(n_495),
.B2(n_477),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_491),
.C(n_484),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_526),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_480),
.Y(n_516)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_478),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_519),
.B(n_527),
.Y(n_534)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_499),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_521),
.A2(n_513),
.B1(n_493),
.B2(n_507),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_498),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_522),
.B(n_523),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_502),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_524),
.B(n_497),
.C(n_501),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_477),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_486),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_504),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_536),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_514),
.A2(n_500),
.B(n_506),
.Y(n_530)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_530),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_533),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_520),
.C(n_524),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_519),
.B(n_497),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_512),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_520),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_516),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_541),
.A2(n_534),
.B(n_531),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_542),
.B(n_528),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_543),
.B(n_539),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g544 ( 
.A1(n_541),
.A2(n_534),
.B(n_536),
.Y(n_544)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_544),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_546),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_549),
.B(n_547),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_550),
.A2(n_548),
.B(n_518),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_538),
.B(n_540),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_552),
.A2(n_525),
.B(n_526),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_553),
.A2(n_483),
.B1(n_525),
.B2(n_549),
.Y(n_554)
);


endmodule