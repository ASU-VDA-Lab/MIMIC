module fake_netlist_6_1740_n_1777 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1777);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1777;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_69),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_81),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_28),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_22),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_59),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_74),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_92),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_56),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_32),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_21),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_95),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_51),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_19),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_10),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_106),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_42),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_18),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_46),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_26),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_48),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_9),
.Y(n_206)
);

BUFx8_ASAP7_75t_SL g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_110),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_38),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_126),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_151),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_138),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_36),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_101),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_26),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_13),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_109),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_137),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_5),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_50),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_147),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_67),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_128),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_31),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_88),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_39),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_58),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_3),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_54),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_122),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_102),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_104),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_99),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_113),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_12),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_3),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_115),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_19),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_2),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_78),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_84),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_89),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_90),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_50),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_97),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_49),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_15),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_134),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_54),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_105),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_82),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_35),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_108),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_41),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_77),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_52),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_57),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_120),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_43),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_91),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_30),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_21),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_37),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_16),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_86),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_131),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_18),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_33),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_156),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_87),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_7),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_73),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_145),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_79),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_83),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_29),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_100),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_15),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_207),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_160),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_209),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_191),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_210),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_191),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_191),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_248),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_191),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_215),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_261),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_216),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_164),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

NOR2xp67_ASAP7_75t_L g333 ( 
.A(n_163),
.B(n_0),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_167),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_250),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_191),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_280),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_177),
.B(n_0),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_241),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_172),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_174),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_229),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_175),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_280),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_305),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_250),
.B(n_1),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_R g353 ( 
.A(n_176),
.B(n_179),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_163),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_218),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_234),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_182),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_298),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_218),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_243),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_177),
.B(n_1),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_187),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_251),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_251),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_180),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_181),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_274),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_183),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_185),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_158),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_190),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_195),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_196),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_158),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_168),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_170),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_168),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_208),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_171),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_171),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_211),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_170),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_304),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_304),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_205),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_313),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_345),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_347),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_308),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_351),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_315),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_316),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_316),
.A2(n_322),
.B(n_320),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_320),
.B(n_205),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_L g413 ( 
.A(n_338),
.B(n_308),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_352),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_322),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_323),
.B(n_217),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_326),
.B(n_221),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_326),
.A2(n_192),
.B(n_189),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_332),
.B(n_221),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_336),
.B(n_219),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_336),
.B(n_224),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

CKINVDCx11_ASAP7_75t_R g431 ( 
.A(n_359),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_338),
.B(n_232),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_333),
.B(n_265),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_333),
.B(n_265),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_381),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_349),
.A2(n_235),
.B1(n_203),
.B2(n_292),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_385),
.B(n_230),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_354),
.A2(n_192),
.B(n_189),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_357),
.B(n_275),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_386),
.B(n_240),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_354),
.B(n_288),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_355),
.B(n_288),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_344),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_360),
.B(n_300),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_361),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_383),
.B(n_244),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_363),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_443),
.B(n_317),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_321),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_406),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_411),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_390),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_401),
.A2(n_348),
.B1(n_328),
.B2(n_325),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_330),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_390),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_414),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_408),
.A2(n_159),
.B(n_157),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_417),
.B(n_331),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_406),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_414),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_394),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_438),
.A2(n_325),
.B1(n_364),
.B2(n_358),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_401),
.B(n_367),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_358),
.Y(n_480)
);

BUFx4f_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_414),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_391),
.B(n_334),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_391),
.B(n_340),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_411),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_388),
.B(n_412),
.Y(n_488)
);

BUFx8_ASAP7_75t_SL g489 ( 
.A(n_397),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_365),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_428),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_452),
.B(n_342),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_346),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_438),
.B(n_369),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_427),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_365),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_424),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_431),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_414),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_429),
.B(n_375),
.Y(n_503)
);

CKINVDCx11_ASAP7_75t_R g504 ( 
.A(n_431),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_429),
.B(n_380),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_427),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_392),
.B(n_384),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_419),
.B(n_300),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_445),
.B(n_366),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_392),
.B(n_387),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_419),
.B(n_246),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_413),
.B(n_169),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_455),
.B(n_378),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_393),
.B(n_446),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_399),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_433),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_448),
.B(n_324),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_399),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_455),
.B(n_377),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_393),
.B(n_446),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_442),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_448),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_412),
.B(n_423),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_413),
.A2(n_290),
.B1(n_178),
.B2(n_198),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_439),
.B(n_312),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_442),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_393),
.B(n_366),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_442),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_169),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_412),
.B(n_254),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_418),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_446),
.B(n_368),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_449),
.B(n_371),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_395),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_412),
.B(n_260),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_439),
.B(n_444),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_388),
.B(n_423),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_395),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_395),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_444),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_423),
.A2(n_178),
.B1(n_290),
.B2(n_212),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_423),
.B(n_425),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_423),
.B(n_319),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_389),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_389),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_449),
.A2(n_266),
.B1(n_236),
.B2(n_233),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_449),
.B(n_201),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_389),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_416),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_425),
.B(n_327),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_418),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_418),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_437),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_416),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_425),
.B(n_263),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_416),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_446),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_449),
.B(n_157),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_425),
.B(n_269),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_416),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_437),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_433),
.B(n_434),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_446),
.B(n_368),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_418),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_425),
.A2(n_212),
.B1(n_198),
.B2(n_310),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_440),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_433),
.A2(n_222),
.B1(n_204),
.B2(n_200),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_409),
.B(n_370),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_433),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_434),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_418),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_426),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_409),
.B(n_329),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_440),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_426),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_410),
.B(n_343),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_408),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_418),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_388),
.Y(n_600)
);

NAND3xp33_ASAP7_75t_L g601 ( 
.A(n_410),
.B(n_159),
.C(n_245),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_388),
.B(n_276),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_R g603 ( 
.A(n_434),
.B(n_188),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_440),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_422),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_396),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_492),
.B(n_434),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_500),
.B(n_257),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_519),
.A2(n_388),
.B1(n_434),
.B2(n_293),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_523),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_523),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_530),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_479),
.B(n_356),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_524),
.B(n_422),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_524),
.B(n_422),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_524),
.B(n_422),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_556),
.A2(n_247),
.B1(n_249),
.B2(n_245),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_481),
.B(n_422),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_519),
.A2(n_293),
.B1(n_283),
.B2(n_184),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_507),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_530),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_598),
.B(n_422),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_600),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_458),
.B(n_420),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_598),
.B(n_422),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_489),
.B(n_201),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_465),
.B(n_193),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_510),
.B(n_199),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_494),
.B(n_422),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_576),
.A2(n_247),
.B1(n_249),
.B2(n_262),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_481),
.B(n_257),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_481),
.B(n_257),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_L g636 ( 
.A1(n_546),
.A2(n_471),
.B1(n_503),
.B2(n_499),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_487),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_506),
.B(n_206),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_551),
.B(n_415),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_488),
.B(n_257),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_600),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_486),
.B(n_220),
.Y(n_643)
);

INVxp33_ASAP7_75t_L g644 ( 
.A(n_527),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_460),
.B(n_415),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_457),
.B(n_226),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g647 ( 
.A1(n_459),
.A2(n_253),
.B1(n_264),
.B2(n_259),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_545),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_497),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_460),
.B(n_415),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_476),
.A2(n_242),
.B1(n_239),
.B2(n_238),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_463),
.B(n_353),
.C(n_258),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_583),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_488),
.B(n_257),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_600),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_461),
.B(n_415),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_470),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_461),
.B(n_415),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_480),
.B(n_194),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_532),
.B(n_420),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_464),
.B(n_396),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_464),
.B(n_398),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_519),
.A2(n_238),
.B1(n_173),
.B2(n_165),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_583),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_497),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_497),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_589),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_483),
.B(n_398),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_483),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_500),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_520),
.B(n_400),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_496),
.B(n_421),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_490),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_520),
.B(n_400),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_480),
.B(n_201),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_488),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_505),
.B(n_257),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_488),
.A2(n_184),
.B1(n_173),
.B2(n_165),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_495),
.B(n_227),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_552),
.B(n_257),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_526),
.B(n_402),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_552),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_552),
.B(n_281),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_526),
.B(n_402),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_505),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_533),
.B(n_299),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_558),
.B(n_303),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_590),
.B(n_403),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_594),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_515),
.B(n_231),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_490),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_531),
.A2(n_228),
.B1(n_284),
.B2(n_225),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_517),
.B(n_403),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_517),
.B(n_404),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_591),
.B(n_225),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_591),
.A2(n_228),
.B1(n_284),
.B2(n_295),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_509),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_511),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_531),
.B(n_239),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_493),
.B(n_256),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_511),
.B(n_404),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_504),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_581),
.A2(n_273),
.B1(n_295),
.B2(n_262),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_538),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_485),
.B(n_270),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_513),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_498),
.B(n_421),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_536),
.B(n_242),
.Y(n_710)
);

AND2x4_ASAP7_75t_SL g711 ( 
.A(n_577),
.B(n_201),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_597),
.B(n_271),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_538),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_498),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_473),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_535),
.B(n_277),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_513),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_603),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_509),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_514),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_541),
.A2(n_267),
.B1(n_283),
.B2(n_278),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_516),
.B(n_405),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_606),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_516),
.B(n_405),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_606),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_535),
.B(n_279),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_501),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_509),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_536),
.B(n_537),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_477),
.B(n_285),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_537),
.B(n_451),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_539),
.B(n_451),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_522),
.B(n_296),
.C(n_307),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_512),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_559),
.B(n_430),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_529),
.B(n_194),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_527),
.B(n_286),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_567),
.A2(n_267),
.B1(n_278),
.B2(n_273),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_539),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_548),
.B(n_451),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_548),
.A2(n_306),
.B1(n_272),
.B2(n_451),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_462),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_476),
.B(n_287),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_521),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_550),
.B(n_272),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_297),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_L g748 ( 
.A(n_574),
.B(n_430),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_540),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_578),
.B(n_306),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_540),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_518),
.B(n_451),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_521),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_588),
.B(n_301),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_540),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_602),
.B(n_440),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_467),
.B(n_435),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_467),
.B(n_472),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_462),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_525),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_564),
.B(n_302),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_SL g762 ( 
.A(n_577),
.B(n_202),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_491),
.B(n_202),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_525),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_601),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_601),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_466),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_491),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_474),
.B(n_309),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_467),
.B(n_435),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_491),
.B(n_202),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_466),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_436),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_491),
.B(n_202),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_528),
.Y(n_775)
);

OR2x2_ASAP7_75t_SL g776 ( 
.A(n_534),
.B(n_213),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_540),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_528),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_549),
.Y(n_779)
);

INVxp33_ASAP7_75t_L g780 ( 
.A(n_557),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_655),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_636),
.B(n_585),
.Y(n_782)
);

O2A1O1Ixp5_ASAP7_75t_L g783 ( 
.A1(n_746),
.A2(n_469),
.B(n_549),
.C(n_553),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_634),
.A2(n_555),
.B(n_554),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_607),
.A2(n_474),
.B(n_568),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_610),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_626),
.B(n_577),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_632),
.A2(n_474),
.B(n_568),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_615),
.A2(n_474),
.B(n_568),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_631),
.B(n_577),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_615),
.A2(n_508),
.B(n_568),
.Y(n_792)
);

BUFx8_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_616),
.A2(n_508),
.B(n_592),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_691),
.B(n_577),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_629),
.B(n_467),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_616),
.A2(n_508),
.B(n_592),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_644),
.B(n_780),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_643),
.B(n_605),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_719),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_747),
.A2(n_605),
.B(n_544),
.C(n_599),
.Y(n_801)
);

OAI21xp33_ASAP7_75t_L g802 ( 
.A1(n_712),
.A2(n_311),
.B(n_223),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_618),
.A2(n_508),
.B(n_592),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_637),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

AO21x1_ASAP7_75t_L g806 ( 
.A1(n_701),
.A2(n_469),
.B(n_553),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_634),
.A2(n_566),
.B(n_555),
.Y(n_807)
);

INVx6_ASAP7_75t_L g808 ( 
.A(n_622),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_639),
.B(n_472),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_735),
.B(n_472),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_612),
.A2(n_540),
.B1(n_544),
.B2(n_599),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_638),
.B(n_491),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_655),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_635),
.A2(n_582),
.B(n_554),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_622),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_618),
.A2(n_566),
.B(n_582),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_620),
.A2(n_592),
.B(n_547),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_638),
.B(n_614),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_620),
.A2(n_547),
.B(n_584),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_645),
.A2(n_656),
.B(n_650),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_736),
.B(n_605),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_623),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_655),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_622),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_658),
.A2(n_547),
.B(n_584),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_660),
.B(n_436),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_726),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_644),
.B(n_472),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_677),
.A2(n_540),
.B1(n_599),
.B2(n_482),
.Y(n_829)
);

CKINVDCx10_ASAP7_75t_R g830 ( 
.A(n_728),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_683),
.A2(n_540),
.B1(n_599),
.B2(n_482),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_765),
.B(n_482),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_614),
.B(n_482),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_686),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_617),
.B(n_502),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_766),
.A2(n_596),
.B(n_573),
.C(n_593),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_617),
.B(n_502),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_649),
.B(n_502),
.Y(n_838)
);

CKINVDCx10_ASAP7_75t_R g839 ( 
.A(n_704),
.Y(n_839)
);

INVx11_ASAP7_75t_L g840 ( 
.A(n_715),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_699),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_699),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_635),
.A2(n_573),
.B(n_596),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_649),
.B(n_502),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_624),
.A2(n_627),
.B(n_752),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_756),
.A2(n_547),
.B(n_584),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_756),
.A2(n_547),
.B(n_584),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_701),
.A2(n_575),
.B(n_593),
.C(n_587),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_710),
.A2(n_575),
.B(n_587),
.C(n_579),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_665),
.B(n_542),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_640),
.A2(n_584),
.B(n_563),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_709),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_710),
.A2(n_579),
.B(n_441),
.C(n_475),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_743),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_673),
.B(n_441),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_674),
.B(n_447),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_730),
.A2(n_542),
.B(n_544),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_743),
.Y(n_858)
);

OAI21xp33_ASAP7_75t_L g859 ( 
.A1(n_744),
.A2(n_213),
.B(n_214),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_665),
.B(n_666),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_693),
.Y(n_861)
);

NOR2x1p5_ASAP7_75t_L g862 ( 
.A(n_652),
.B(n_214),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_657),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_746),
.A2(n_475),
.B(n_478),
.C(n_484),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_730),
.A2(n_542),
.B(n_544),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_758),
.A2(n_569),
.B(n_542),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_751),
.A2(n_563),
.B(n_569),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_613),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_608),
.A2(n_563),
.B(n_569),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_659),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_759),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_628),
.B(n_762),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_780),
.B(n_563),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_663),
.A2(n_621),
.B1(n_700),
.B2(n_671),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_666),
.B(n_569),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_661),
.A2(n_468),
.B(n_478),
.Y(n_876)
);

AO21x1_ASAP7_75t_L g877 ( 
.A1(n_608),
.A2(n_223),
.B(n_252),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_759),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_678),
.A2(n_604),
.B(n_595),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_709),
.B(n_630),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_738),
.B(n_447),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_638),
.A2(n_468),
.B1(n_484),
.B2(n_586),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_709),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_767),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_699),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_659),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_751),
.A2(n_571),
.B(n_595),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_680),
.A2(n_604),
.B(n_586),
.C(n_580),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_646),
.A2(n_580),
.B(n_572),
.C(n_571),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_642),
.B(n_543),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_648),
.B(n_543),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_699),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_669),
.A2(n_572),
.B1(n_570),
.B2(n_561),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_659),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_751),
.A2(n_570),
.B(n_561),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_653),
.B(n_560),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_664),
.B(n_560),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_776),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_748),
.A2(n_565),
.B1(n_456),
.B2(n_454),
.Y(n_899)
);

AO21x1_ASAP7_75t_L g900 ( 
.A1(n_678),
.A2(n_705),
.B(n_750),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_717),
.B(n_565),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_745),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_753),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_669),
.B(n_565),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_760),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_706),
.B(n_450),
.Y(n_906)
);

O2A1O1Ixp5_ASAP7_75t_L g907 ( 
.A1(n_750),
.A2(n_456),
.B(n_454),
.C(n_453),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_671),
.B(n_456),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_687),
.B(n_456),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_687),
.A2(n_291),
.B1(n_252),
.B2(n_255),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_767),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_700),
.A2(n_291),
.B1(n_255),
.B2(n_268),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_720),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_625),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_708),
.B(n_718),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_708),
.B(n_454),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_727),
.B(n_453),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_642),
.B(n_107),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_751),
.A2(n_454),
.B(n_450),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_772),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_718),
.B(n_310),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_667),
.B(n_294),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_670),
.B(n_294),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_732),
.A2(n_370),
.B(n_289),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_733),
.A2(n_289),
.B(n_282),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_741),
.A2(n_282),
.B(n_268),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_625),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_740),
.B(n_237),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_737),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_713),
.B(n_4),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_714),
.B(n_237),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_749),
.B(n_777),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_697),
.A2(n_237),
.B(n_5),
.C(n_6),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_716),
.B(n_237),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_721),
.B(n_4),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_772),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_662),
.A2(n_150),
.B(n_146),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_694),
.A2(n_141),
.B1(n_135),
.B2(n_130),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_764),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_690),
.B(n_6),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_742),
.B(n_8),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_609),
.B(n_10),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_697),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_769),
.B(n_11),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_703),
.A2(n_127),
.B(n_121),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_755),
.B(n_93),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_720),
.B(n_11),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_692),
.B(n_13),
.C(n_14),
.Y(n_948)
);

AND2x2_ASAP7_75t_SL g949 ( 
.A(n_711),
.B(n_676),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_737),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_668),
.A2(n_80),
.B(n_76),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_755),
.B(n_71),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_723),
.A2(n_68),
.B(n_65),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_725),
.A2(n_62),
.B(n_60),
.Y(n_954)
);

AOI21x1_ASAP7_75t_L g955 ( 
.A1(n_641),
.A2(n_14),
.B(n_17),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_720),
.B(n_17),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_720),
.B(n_23),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_672),
.A2(n_23),
.B(n_24),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_729),
.B(n_25),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_641),
.A2(n_27),
.B(n_29),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_775),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_675),
.A2(n_31),
.B(n_33),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_654),
.A2(n_34),
.B(n_36),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_729),
.B(n_707),
.Y(n_964)
);

BUFx4f_ASAP7_75t_L g965 ( 
.A(n_737),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_754),
.B(n_34),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_702),
.B(n_39),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_731),
.B(n_55),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_729),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_755),
.B(n_41),
.Y(n_970)
);

AOI33xp33_ASAP7_75t_L g971 ( 
.A1(n_651),
.A2(n_43),
.A3(n_44),
.B1(n_45),
.B2(n_47),
.B3(n_51),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_917),
.B(n_761),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_902),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_854),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_840),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_967),
.A2(n_734),
.B(n_739),
.C(n_722),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_863),
.Y(n_978)
);

AOI21xp33_ASAP7_75t_L g979 ( 
.A1(n_966),
.A2(n_684),
.B(n_688),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_903),
.Y(n_980)
);

AO32x1_ASAP7_75t_L g981 ( 
.A1(n_968),
.A2(n_698),
.A3(n_633),
.B1(n_711),
.B2(n_778),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_905),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_964),
.A2(n_682),
.B(n_685),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_966),
.A2(n_619),
.B(n_695),
.C(n_696),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_868),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_846),
.A2(n_768),
.B(n_757),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_939),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_845),
.A2(n_654),
.B(n_681),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_791),
.A2(n_681),
.B(n_770),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_SL g990 ( 
.A(n_800),
.B(n_647),
.C(n_774),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_SL g991 ( 
.A1(n_946),
.A2(n_684),
.B(n_774),
.C(n_771),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_861),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_852),
.B(n_749),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_961),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_906),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_798),
.B(n_689),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_805),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_858),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_967),
.A2(n_689),
.B(n_688),
.C(n_771),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_SL g1000 ( 
.A1(n_949),
.A2(n_679),
.B1(n_777),
.B2(n_755),
.Y(n_1000)
);

NOR2x1p5_ASAP7_75t_SL g1001 ( 
.A(n_816),
.B(n_876),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_872),
.B(n_729),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_881),
.B(n_779),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_841),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_798),
.B(n_763),
.C(n_773),
.Y(n_1005)
);

CKINVDCx8_ASAP7_75t_R g1006 ( 
.A(n_839),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_805),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_826),
.B(n_763),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_787),
.A2(n_768),
.B1(n_47),
.B2(n_52),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_805),
.Y(n_1010)
);

CKINVDCx8_ASAP7_75t_R g1011 ( 
.A(n_830),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_795),
.A2(n_768),
.B1(n_44),
.B2(n_53),
.Y(n_1012)
);

AO32x2_ASAP7_75t_L g1013 ( 
.A1(n_910),
.A2(n_53),
.A3(n_912),
.B1(n_893),
.B2(n_882),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_793),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_796),
.A2(n_799),
.B(n_785),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_805),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_898),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_943),
.A2(n_944),
.B(n_795),
.C(n_873),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_813),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_886),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_809),
.A2(n_820),
.B(n_788),
.Y(n_1021)
);

AO21x1_ASAP7_75t_L g1022 ( 
.A1(n_945),
.A2(n_954),
.B(n_782),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_949),
.B(n_892),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_855),
.B(n_856),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_802),
.A2(n_859),
.B(n_789),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_965),
.B(n_943),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_929),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_786),
.B(n_822),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_L g1029 ( 
.A1(n_900),
.A2(n_877),
.B(n_801),
.C(n_806),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_793),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_821),
.A2(n_818),
.B(n_901),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_950),
.B(n_861),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_906),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_L g1034 ( 
.A(n_928),
.B(n_931),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_959),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_950),
.B(n_883),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_818),
.A2(n_901),
.B(n_874),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_827),
.B(n_873),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_783),
.A2(n_874),
.B(n_860),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_L g1040 ( 
.A(n_932),
.B(n_918),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_L g1041 ( 
.A(n_932),
.B(n_918),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_808),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_880),
.A2(n_915),
.B1(n_942),
.B2(n_914),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_871),
.Y(n_1044)
);

AO21x1_ASAP7_75t_L g1045 ( 
.A1(n_970),
.A2(n_960),
.B(n_963),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_828),
.A2(n_927),
.B1(n_914),
.B2(n_862),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_SL g1047 ( 
.A1(n_808),
.A2(n_870),
.B1(n_894),
.B2(n_824),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_965),
.B(n_927),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_808),
.Y(n_1049)
);

AO21x2_ASAP7_75t_L g1050 ( 
.A1(n_784),
.A2(n_814),
.B(n_843),
.Y(n_1050)
);

AOI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_828),
.A2(n_934),
.B(n_940),
.Y(n_1051)
);

NAND2xp33_ASAP7_75t_R g1052 ( 
.A(n_892),
.B(n_959),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_970),
.A2(n_921),
.B(n_922),
.C(n_923),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_815),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_930),
.B(n_935),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_930),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_925),
.A2(n_926),
.B(n_941),
.C(n_832),
.Y(n_1057)
);

OR2x2_ASAP7_75t_L g1058 ( 
.A(n_834),
.B(n_947),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_891),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_956),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_896),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_935),
.B(n_897),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_878),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_884),
.B(n_911),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_869),
.A2(n_797),
.B(n_803),
.Y(n_1065)
);

AND3x1_ASAP7_75t_SL g1066 ( 
.A(n_971),
.B(n_948),
.C(n_933),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_L g1067 ( 
.A(n_813),
.B(n_841),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_957),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_924),
.A2(n_836),
.B(n_958),
.C(n_962),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_920),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_936),
.B(n_813),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_813),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_841),
.B(n_885),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_783),
.A2(n_864),
.B(n_907),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_790),
.A2(n_792),
.B(n_794),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_781),
.B(n_823),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_946),
.A2(n_952),
.B(n_888),
.C(n_938),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_810),
.B(n_781),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_952),
.A2(n_889),
.B(n_853),
.C(n_907),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_823),
.B(n_969),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_811),
.A2(n_831),
.B1(n_829),
.B2(n_812),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_841),
.Y(n_1082)
);

AOI21xp33_ASAP7_75t_L g1083 ( 
.A1(n_833),
.A2(n_838),
.B(n_850),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_842),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_842),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_842),
.B(n_885),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_913),
.B(n_969),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_908),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_825),
.A2(n_817),
.B(n_879),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_842),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_909),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_851),
.A2(n_819),
.B(n_847),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_885),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_807),
.A2(n_919),
.B(n_887),
.C(n_895),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_916),
.A2(n_867),
.B(n_812),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_885),
.B(n_913),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_848),
.A2(n_849),
.B(n_865),
.C(n_857),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_890),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_890),
.A2(n_835),
.B1(n_837),
.B2(n_844),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_904),
.Y(n_1100)
);

OAI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_899),
.A2(n_875),
.B1(n_955),
.B2(n_937),
.C(n_951),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_953),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_866),
.B(n_864),
.Y(n_1103)
);

NOR2x1_ASAP7_75t_R g1104 ( 
.A(n_808),
.B(n_504),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_R g1105 ( 
.A(n_800),
.B(n_406),
.Y(n_1105)
);

INVx3_ASAP7_75t_SL g1106 ( 
.A(n_808),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_964),
.A2(n_607),
.B(n_632),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_826),
.B(n_660),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_781),
.B(n_823),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_966),
.A2(n_631),
.B1(n_629),
.B2(n_967),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_798),
.B(n_691),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_966),
.A2(n_967),
.B1(n_968),
.B2(n_631),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_966),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_854),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_868),
.B(n_473),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_932),
.B(n_780),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_840),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_854),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_854),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_826),
.B(n_660),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_949),
.B(n_636),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_854),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_917),
.B(n_626),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_917),
.B(n_626),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_964),
.A2(n_607),
.B(n_632),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1075),
.A2(n_1092),
.B(n_1095),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_997),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1124),
.B2(n_1123),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_977),
.A2(n_979),
.B(n_1018),
.C(n_1121),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_L g1132 ( 
.A1(n_1055),
.A2(n_1056),
.B1(n_1111),
.B2(n_972),
.C(n_1009),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_1006),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1024),
.B(n_1108),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1120),
.B(n_1038),
.Y(n_1135)
);

INVx3_ASAP7_75t_SL g1136 ( 
.A(n_1030),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1095),
.A2(n_1089),
.B(n_988),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_996),
.A2(n_1116),
.B1(n_1045),
.B2(n_1025),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1105),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1011),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1003),
.B(n_1059),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1061),
.B(n_1062),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1022),
.A2(n_1065),
.A3(n_1089),
.B(n_1015),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_SL g1145 ( 
.A(n_999),
.B(n_1012),
.C(n_1002),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_988),
.A2(n_1065),
.B(n_1074),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_999),
.B(n_1051),
.C(n_1005),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_980),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_SL g1149 ( 
.A1(n_1026),
.A2(n_1008),
.B(n_1094),
.C(n_1081),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1035),
.B(n_1036),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_1115),
.A2(n_984),
.B(n_1053),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1034),
.B(n_1060),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_1032),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_973),
.B(n_1076),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1076),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1113),
.B(n_995),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_997),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1077),
.A2(n_1053),
.B(n_984),
.C(n_1037),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1100),
.B(n_1046),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1113),
.B(n_1033),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1103),
.A2(n_1015),
.B(n_1029),
.Y(n_1161)
);

AOI31xp67_ASAP7_75t_L g1162 ( 
.A1(n_1101),
.A2(n_981),
.A3(n_1073),
.B(n_1086),
.Y(n_1162)
);

BUFx2_ASAP7_75t_R g1163 ( 
.A(n_1106),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1068),
.B(n_1028),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_978),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_SL g1166 ( 
.A1(n_1043),
.A2(n_1048),
.B1(n_1077),
.B2(n_1037),
.C(n_982),
.Y(n_1166)
);

INVxp67_ASAP7_75t_L g1167 ( 
.A(n_992),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1000),
.A2(n_1052),
.B1(n_1066),
.B2(n_1058),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1069),
.A2(n_1057),
.B(n_989),
.C(n_983),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_987),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_985),
.B(n_1027),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1014),
.A2(n_1047),
.B1(n_1020),
.B2(n_1017),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_994),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_990),
.A2(n_1041),
.B1(n_1040),
.B2(n_993),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1088),
.B(n_1091),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_983),
.B(n_1031),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1097),
.A2(n_1031),
.A3(n_1098),
.B(n_981),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1069),
.B(n_1057),
.C(n_991),
.Y(n_1178)
);

BUFx2_ASAP7_75t_R g1179 ( 
.A(n_1106),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_1039),
.B(n_1078),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1102),
.A2(n_1067),
.B(n_1050),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1050),
.A2(n_1079),
.B(n_1083),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1054),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1079),
.A2(n_976),
.B(n_1063),
.C(n_1042),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1023),
.B(n_1117),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_993),
.B(n_1049),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_975),
.A2(n_1122),
.B1(n_998),
.B2(n_1119),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_1072),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1044),
.B(n_1118),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1071),
.A2(n_1096),
.B(n_1114),
.C(n_1070),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1001),
.A2(n_1064),
.B(n_1099),
.C(n_1084),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1109),
.A2(n_1080),
.B(n_1087),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1098),
.A2(n_981),
.A3(n_1013),
.B(n_1019),
.Y(n_1193)
);

OAI22x1_ASAP7_75t_L g1194 ( 
.A1(n_1085),
.A2(n_1093),
.B1(n_1090),
.B2(n_1082),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1016),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1013),
.A2(n_1016),
.A3(n_1019),
.B(n_1004),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1004),
.Y(n_1197)
);

AO32x2_ASAP7_75t_L g1198 ( 
.A1(n_1013),
.A2(n_1109),
.A3(n_1010),
.B1(n_1007),
.B2(n_1104),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1013),
.A2(n_1022),
.A3(n_1045),
.B(n_1065),
.Y(n_1199)
);

INVx8_ASAP7_75t_L g1200 ( 
.A(n_1010),
.Y(n_1200)
);

CKINVDCx11_ASAP7_75t_R g1201 ( 
.A(n_1010),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1029),
.A2(n_1074),
.B(n_1021),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1115),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_973),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1022),
.A2(n_1045),
.A3(n_1065),
.B(n_1089),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1110),
.A2(n_966),
.B1(n_967),
.B2(n_1112),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1110),
.B(n_691),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1110),
.A2(n_966),
.B(n_1112),
.C(n_967),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_973),
.B(n_1076),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1124),
.B2(n_1123),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1112),
.A2(n_966),
.B(n_479),
.C(n_629),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1018),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_1018),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1110),
.A2(n_966),
.B1(n_967),
.B2(n_1112),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_977),
.A2(n_1110),
.B(n_979),
.C(n_1018),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_973),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_997),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1110),
.B(n_691),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1006),
.B(n_489),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_SL g1224 ( 
.A1(n_977),
.A2(n_1110),
.B(n_979),
.C(n_1018),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_992),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_1105),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1110),
.A2(n_966),
.B(n_1112),
.C(n_967),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1108),
.B(n_1120),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_974),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_974),
.Y(n_1234)
);

NOR2x1_ASAP7_75t_R g1235 ( 
.A(n_1030),
.B(n_504),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_974),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_974),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_992),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1110),
.A2(n_966),
.B(n_1112),
.C(n_967),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_973),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1124),
.B2(n_1123),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_SL g1247 ( 
.A1(n_1045),
.A2(n_963),
.B(n_960),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1110),
.B(n_719),
.Y(n_1248)
);

OAI21xp33_ASAP7_75t_L g1249 ( 
.A1(n_1110),
.A2(n_1112),
.B(n_966),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_SL g1250 ( 
.A1(n_979),
.A2(n_1121),
.B(n_1051),
.C(n_750),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1112),
.A2(n_966),
.B1(n_744),
.B2(n_479),
.C(n_651),
.Y(n_1253)
);

BUFx8_ASAP7_75t_L g1254 ( 
.A(n_973),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_974),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1076),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_986),
.A2(n_1075),
.B(n_1092),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1262)
);

AOI221x1_ASAP7_75t_L g1263 ( 
.A1(n_979),
.A2(n_966),
.B1(n_967),
.B2(n_944),
.C(n_629),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1021),
.Y(n_1264)
);

AO32x2_ASAP7_75t_L g1265 ( 
.A1(n_1009),
.A2(n_1043),
.A3(n_1081),
.B1(n_912),
.B2(n_910),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1110),
.A2(n_966),
.B1(n_1112),
.B2(n_967),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1124),
.B2(n_1123),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1254),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1171),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1141),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1208),
.A2(n_1217),
.B1(n_1253),
.B2(n_1215),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1189),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1148),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1266),
.A2(n_1217),
.B1(n_1208),
.B2(n_1243),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1183),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1165),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1173),
.Y(n_1278)
);

OAI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1139),
.A2(n_1209),
.B1(n_1222),
.B2(n_1168),
.Y(n_1279)
);

CKINVDCx11_ASAP7_75t_R g1280 ( 
.A(n_1133),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1216),
.A2(n_1168),
.B1(n_1139),
.B2(n_1135),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1207),
.B(n_1237),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1254),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1249),
.A2(n_1248),
.B1(n_1227),
.B2(n_1210),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1232),
.Y(n_1285)
);

INVx6_ASAP7_75t_L g1286 ( 
.A(n_1129),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1130),
.A2(n_1268),
.B1(n_1212),
.B2(n_1246),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1205),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1129),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1219),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1234),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1236),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1136),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_1186),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1226),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1241),
.Y(n_1296)
);

INVx6_ASAP7_75t_SL g1297 ( 
.A(n_1153),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1140),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1244),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1249),
.A2(n_1213),
.B1(n_1174),
.B2(n_1143),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1188),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1228),
.B(n_1150),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1174),
.A2(n_1152),
.B1(n_1142),
.B2(n_1132),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1256),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1187),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1145),
.A2(n_1267),
.B1(n_1261),
.B2(n_1258),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1247),
.A2(n_1147),
.B1(n_1172),
.B2(n_1178),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1187),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1164),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1175),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1134),
.B(n_1156),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1197),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1147),
.A2(n_1172),
.B1(n_1178),
.B2(n_1245),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1201),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1151),
.A2(n_1159),
.B1(n_1180),
.B2(n_1176),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1190),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1163),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1204),
.A2(n_1182),
.B1(n_1242),
.B2(n_1225),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1160),
.A2(n_1202),
.B1(n_1153),
.B2(n_1146),
.Y(n_1319)
);

BUFx4_ASAP7_75t_R g1320 ( 
.A(n_1179),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1202),
.A2(n_1263),
.B1(n_1167),
.B2(n_1194),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1223),
.A2(n_1198),
.B1(n_1224),
.B2(n_1218),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1126),
.A2(n_1203),
.B1(n_1264),
.B2(n_1220),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1196),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1154),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1158),
.A2(n_1169),
.B(n_1184),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1185),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1138),
.A2(n_1252),
.B1(n_1262),
.B2(n_1229),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1198),
.A2(n_1181),
.B1(n_1265),
.B2(n_1131),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1166),
.B(n_1257),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1193),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1235),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1235),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1211),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1200),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1230),
.A2(n_1233),
.B1(n_1259),
.B2(n_1231),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1198),
.A2(n_1265),
.B1(n_1161),
.B2(n_1137),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1157),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1191),
.A2(n_1257),
.B1(n_1155),
.B2(n_1195),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1265),
.A2(n_1255),
.B1(n_1250),
.B2(n_1128),
.Y(n_1340)
);

INVx8_ASAP7_75t_L g1341 ( 
.A(n_1157),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1221),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1192),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1149),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1162),
.A2(n_1199),
.B1(n_1177),
.B2(n_1193),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1127),
.A2(n_1214),
.B1(n_1251),
.B2(n_1240),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1199),
.B(n_1206),
.Y(n_1347)
);

INVx8_ASAP7_75t_L g1348 ( 
.A(n_1260),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1206),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_1193),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1144),
.A2(n_1110),
.B1(n_1112),
.B2(n_1266),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1144),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1238),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1239),
.A2(n_1110),
.B1(n_1112),
.B2(n_1266),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1266),
.B2(n_1217),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1266),
.B2(n_1217),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1254),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1228),
.B(n_1150),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1171),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1362)
);

BUFx4f_ASAP7_75t_SL g1363 ( 
.A(n_1133),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1170),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1254),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1171),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1266),
.B2(n_1217),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1133),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1170),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1254),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1266),
.B2(n_1217),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1170),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1209),
.A2(n_1222),
.B1(n_966),
.B2(n_1216),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1141),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_SL g1377 ( 
.A(n_1163),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1228),
.B(n_1150),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1266),
.A2(n_1110),
.B1(n_1112),
.B2(n_1208),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1249),
.A2(n_1253),
.B1(n_1266),
.B2(n_1217),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1170),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1133),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1323),
.A2(n_1336),
.B(n_1328),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1270),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1324),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1375),
.A2(n_1313),
.B1(n_1368),
.B2(n_1355),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1353),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1331),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1347),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1287),
.B(n_1349),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1287),
.B(n_1329),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1375),
.A2(n_1366),
.B1(n_1356),
.B2(n_1379),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1361),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1350),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1329),
.B(n_1315),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1367),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1344),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1360),
.A2(n_1371),
.B1(n_1362),
.B2(n_1357),
.C(n_1373),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1345),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1315),
.B(n_1319),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1275),
.A2(n_1351),
.B1(n_1300),
.B2(n_1354),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1286),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1282),
.B(n_1306),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1316),
.B(n_1305),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1352),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1286),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1319),
.B(n_1308),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1348),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1323),
.A2(n_1336),
.B(n_1328),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1274),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1278),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1296),
.B(n_1285),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1291),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1326),
.A2(n_1272),
.B(n_1281),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1302),
.B(n_1359),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1273),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1292),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1348),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1378),
.B(n_1311),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1348),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1310),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1339),
.B(n_1284),
.Y(n_1424)
);

AO21x1_ASAP7_75t_L g1425 ( 
.A1(n_1272),
.A2(n_1281),
.B(n_1303),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1321),
.B(n_1318),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1304),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1363),
.B(n_1382),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1313),
.A2(n_1373),
.B1(n_1355),
.B2(n_1357),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1330),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1286),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1337),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1289),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1374),
.A2(n_1381),
.B(n_1340),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1289),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1337),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1346),
.A2(n_1321),
.B(n_1312),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1364),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1309),
.Y(n_1439)
);

NAND2xp33_ASAP7_75t_SL g1440 ( 
.A(n_1295),
.B(n_1317),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1370),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1288),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1340),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1307),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1279),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1318),
.B(n_1368),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1325),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1307),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1280),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1322),
.B(n_1380),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1322),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1346),
.A2(n_1380),
.B(n_1289),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1294),
.B(n_1301),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1377),
.A2(n_1327),
.B1(n_1297),
.B2(n_1290),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1290),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1341),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1338),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1294),
.B(n_1299),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1341),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1335),
.B(n_1342),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1334),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1277),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1277),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1297),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1405),
.B(n_1358),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1410),
.B(n_1365),
.Y(n_1466)
);

OA21x2_ASAP7_75t_L g1467 ( 
.A1(n_1437),
.A2(n_1376),
.B(n_1271),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1432),
.B(n_1365),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1432),
.B(n_1269),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1401),
.B(n_1436),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1436),
.B(n_1269),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1410),
.B(n_1283),
.Y(n_1472)
);

AND2x2_ASAP7_75t_SL g1473 ( 
.A(n_1391),
.B(n_1320),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1402),
.B(n_1269),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1387),
.A2(n_1298),
.B1(n_1320),
.B2(n_1377),
.C(n_1382),
.Y(n_1475)
);

AND2x2_ASAP7_75t_SL g1476 ( 
.A(n_1391),
.B(n_1372),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1429),
.A2(n_1372),
.B1(n_1333),
.B2(n_1332),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1412),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_SL g1480 ( 
.A1(n_1400),
.A2(n_1314),
.B(n_1293),
.C(n_1363),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1402),
.B(n_1276),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1416),
.A2(n_1369),
.B(n_1393),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1449),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1409),
.B(n_1396),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1383),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1424),
.A2(n_1403),
.B(n_1392),
.C(n_1450),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1425),
.A2(n_1444),
.B1(n_1448),
.B2(n_1450),
.C(n_1392),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1409),
.B(n_1396),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_SL g1489 ( 
.A(n_1434),
.B(n_1426),
.Y(n_1489)
);

O2A1O1Ixp33_ASAP7_75t_SL g1490 ( 
.A1(n_1444),
.A2(n_1448),
.B(n_1424),
.C(n_1446),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1430),
.B(n_1394),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1383),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1413),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1462),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1397),
.B(n_1415),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1399),
.A2(n_1446),
.B1(n_1407),
.B2(n_1451),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1415),
.B(n_1419),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1401),
.B(n_1389),
.Y(n_1498)
);

AOI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1425),
.A2(n_1445),
.B1(n_1451),
.B2(n_1421),
.C(n_1443),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1383),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1388),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_SL g1504 ( 
.A1(n_1407),
.A2(n_1453),
.B(n_1463),
.C(n_1426),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1462),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1427),
.Y(n_1506)
);

AND2x6_ASAP7_75t_L g1507 ( 
.A(n_1420),
.B(n_1422),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1452),
.A2(n_1406),
.B(n_1442),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1437),
.A2(n_1443),
.B(n_1452),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1414),
.B(n_1418),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1414),
.B(n_1390),
.Y(n_1511)
);

NAND4xp25_ASAP7_75t_L g1512 ( 
.A(n_1417),
.B(n_1399),
.C(n_1414),
.D(n_1441),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1399),
.B(n_1428),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_SL g1514 ( 
.A(n_1454),
.B(n_1462),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1422),
.B(n_1398),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1460),
.B(n_1455),
.Y(n_1516)
);

AO32x2_ASAP7_75t_L g1517 ( 
.A1(n_1404),
.A2(n_1435),
.A3(n_1408),
.B1(n_1431),
.B2(n_1433),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1398),
.B(n_1395),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1507),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1507),
.B(n_1515),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1512),
.B(n_1447),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1517),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1485),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1485),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1507),
.B(n_1515),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1492),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1498),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1482),
.A2(n_1384),
.B1(n_1411),
.B2(n_1406),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1500),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1474),
.B(n_1457),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1487),
.A2(n_1411),
.B1(n_1384),
.B2(n_1463),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1507),
.Y(n_1532)
);

NAND4xp25_ASAP7_75t_L g1533 ( 
.A(n_1499),
.B(n_1461),
.C(n_1440),
.D(n_1464),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1475),
.A2(n_1384),
.B1(n_1411),
.B2(n_1438),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1517),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1509),
.B(n_1511),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1511),
.B(n_1384),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1498),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1477),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1467),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1529),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1529),
.Y(n_1544)
);

OAI33xp33_ASAP7_75t_L g1545 ( 
.A1(n_1533),
.A2(n_1496),
.A3(n_1502),
.B1(n_1495),
.B2(n_1491),
.B3(n_1470),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1520),
.B(n_1484),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1523),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1523),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1523),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1524),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1520),
.B(n_1484),
.Y(n_1551)
);

CKINVDCx16_ASAP7_75t_R g1552 ( 
.A(n_1532),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1527),
.B(n_1470),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1532),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_SL g1555 ( 
.A(n_1532),
.B(n_1497),
.Y(n_1555)
);

OR2x2_ASAP7_75t_SL g1556 ( 
.A(n_1541),
.B(n_1467),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1527),
.B(n_1488),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1524),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1540),
.Y(n_1559)
);

OAI33xp33_ASAP7_75t_L g1560 ( 
.A1(n_1533),
.A2(n_1465),
.A3(n_1493),
.B1(n_1479),
.B2(n_1506),
.B3(n_1386),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1533),
.A2(n_1473),
.B1(n_1478),
.B2(n_1481),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1531),
.A2(n_1486),
.B1(n_1473),
.B2(n_1478),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1532),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1481),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1520),
.B(n_1525),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1488),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1531),
.A2(n_1486),
.B1(n_1480),
.B2(n_1514),
.C(n_1508),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1534),
.A2(n_1478),
.B1(n_1490),
.B2(n_1480),
.C(n_1504),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1539),
.B(n_1510),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1519),
.B(n_1518),
.Y(n_1571)
);

NOR3xp33_ASAP7_75t_L g1572 ( 
.A(n_1521),
.B(n_1490),
.C(n_1474),
.Y(n_1572)
);

OAI222xp33_ASAP7_75t_L g1573 ( 
.A1(n_1528),
.A2(n_1468),
.B1(n_1471),
.B2(n_1469),
.C1(n_1494),
.C2(n_1516),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1522),
.B(n_1501),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1526),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1547),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1553),
.B(n_1539),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1566),
.B(n_1519),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1547),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1543),
.B(n_1522),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1575),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1542),
.B(n_1522),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.B(n_1535),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1542),
.B(n_1535),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1566),
.B(n_1519),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1574),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1501),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1567),
.B(n_1535),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1545),
.B(n_1513),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1548),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1574),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1549),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1546),
.B(n_1519),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1550),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1546),
.B(n_1537),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1551),
.B(n_1537),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1557),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1579),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1579),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1596),
.B(n_1554),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1601),
.B(n_1557),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1580),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1581),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1596),
.B(n_1563),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1581),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1591),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1580),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1601),
.B(n_1590),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1580),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1589),
.B(n_1555),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1539),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1570),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1588),
.A2(n_1562),
.B1(n_1568),
.B2(n_1564),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1602),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1603),
.B(n_1570),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1596),
.B(n_1578),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1538),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1589),
.B(n_1555),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1578),
.B(n_1563),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1602),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1588),
.B(n_1562),
.C(n_1561),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1576),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1577),
.B(n_1599),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1589),
.B(n_1571),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1576),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1583),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1587),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1583),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1594),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1592),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1592),
.B(n_1565),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1582),
.B(n_1571),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1595),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1615),
.B(n_1619),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1595),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1650)
);

AND3x2_ASAP7_75t_L g1651 ( 
.A(n_1642),
.B(n_1572),
.C(n_1569),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1587),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1619),
.B(n_1572),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1621),
.B(n_1569),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1608),
.B(n_1598),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1598),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1613),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1633),
.B(n_1597),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1637),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1640),
.B(n_1604),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1640),
.B(n_1587),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1637),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1621),
.B(n_1598),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1607),
.B(n_1578),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1620),
.B(n_1597),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1613),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1632),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1607),
.B(n_1586),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1631),
.B(n_1600),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1642),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1634),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1632),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1639),
.A2(n_1568),
.B(n_1593),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1643),
.Y(n_1676)
);

AND2x2_ASAP7_75t_SL g1677 ( 
.A(n_1618),
.B(n_1476),
.Y(n_1677)
);

INVx4_ASAP7_75t_L g1678 ( 
.A(n_1611),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1635),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1605),
.A2(n_1528),
.B(n_1534),
.Y(n_1681)
);

CKINVDCx14_ASAP7_75t_R g1682 ( 
.A(n_1672),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1680),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1648),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1675),
.A2(n_1593),
.B(n_1610),
.C(n_1612),
.Y(n_1687)
);

OAI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1681),
.A2(n_1573),
.A3(n_1593),
.B(n_1626),
.Y(n_1688)
);

NOR4xp25_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1622),
.C(n_1605),
.D(n_1617),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1651),
.B(n_1483),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1677),
.B(n_1618),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1681),
.A2(n_1664),
.B(n_1670),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1677),
.A2(n_1556),
.B1(n_1476),
.B2(n_1618),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1677),
.A2(n_1626),
.B(n_1610),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1483),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1678),
.Y(n_1696)
);

NOR4xp25_ASAP7_75t_L g1697 ( 
.A(n_1657),
.B(n_1622),
.C(n_1628),
.D(n_1606),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1678),
.Y(n_1698)
);

AOI32xp33_ASAP7_75t_L g1699 ( 
.A1(n_1648),
.A2(n_1626),
.A3(n_1627),
.B1(n_1624),
.B2(n_1645),
.Y(n_1699)
);

INVxp33_ASAP7_75t_L g1700 ( 
.A(n_1650),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_1624),
.Y(n_1702)
);

NOR2xp67_ASAP7_75t_L g1703 ( 
.A(n_1678),
.B(n_1627),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1655),
.B(n_1623),
.Y(n_1704)
);

OAI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1660),
.A2(n_1623),
.B(n_1521),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1659),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1652),
.A2(n_1556),
.B1(n_1586),
.B2(n_1645),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1684),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1701),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1682),
.A2(n_1652),
.B(n_1660),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1706),
.Y(n_1711)
);

OAI322xp33_ASAP7_75t_L g1712 ( 
.A1(n_1682),
.A2(n_1667),
.A3(n_1657),
.B1(n_1668),
.B2(n_1676),
.C1(n_1674),
.C2(n_1679),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1690),
.A2(n_1652),
.B(n_1667),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1690),
.A2(n_1652),
.B(n_1659),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1689),
.A2(n_1652),
.B(n_1661),
.Y(n_1715)
);

XOR2x2_ASAP7_75t_L g1716 ( 
.A(n_1692),
.B(n_1505),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1687),
.B(n_1674),
.C(n_1668),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1697),
.A2(n_1679),
.B(n_1676),
.C(n_1656),
.Y(n_1718)
);

NOR4xp25_ASAP7_75t_L g1719 ( 
.A(n_1685),
.B(n_1663),
.C(n_1662),
.D(n_1673),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1706),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1688),
.A2(n_1661),
.B(n_1494),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1695),
.Y(n_1722)
);

OAI33xp33_ASAP7_75t_L g1723 ( 
.A1(n_1696),
.A2(n_1662),
.A3(n_1663),
.B1(n_1612),
.B2(n_1628),
.B3(n_1606),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1686),
.B(n_1700),
.Y(n_1724)
);

OAI21xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1691),
.A2(n_1669),
.B(n_1665),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1702),
.B(n_1665),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1725),
.A2(n_1691),
.B1(n_1695),
.B2(n_1703),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1715),
.A2(n_1694),
.B1(n_1693),
.B2(n_1707),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1720),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1717),
.B(n_1713),
.C(n_1721),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1719),
.B(n_1696),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1724),
.Y(n_1733)
);

OAI211xp5_ASAP7_75t_SL g1734 ( 
.A1(n_1722),
.A2(n_1699),
.B(n_1705),
.C(n_1698),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1710),
.A2(n_1698),
.B1(n_1671),
.B2(n_1673),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1726),
.A2(n_1683),
.B1(n_1661),
.B2(n_1671),
.Y(n_1736)
);

NOR2xp67_ASAP7_75t_L g1737 ( 
.A(n_1733),
.B(n_1714),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1727),
.B(n_1713),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1736),
.B(n_1716),
.Y(n_1739)
);

NAND2xp33_ASAP7_75t_R g1740 ( 
.A(n_1732),
.B(n_1714),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1729),
.Y(n_1741)
);

NAND4xp25_ASAP7_75t_SL g1742 ( 
.A(n_1731),
.B(n_1718),
.C(n_1712),
.D(n_1704),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1730),
.C(n_1708),
.D(n_1709),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1735),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1728),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1742),
.A2(n_1723),
.B1(n_1661),
.B2(n_1617),
.C(n_1614),
.Y(n_1746)
);

AOI322xp5_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1582),
.A3(n_1584),
.B1(n_1585),
.B2(n_1669),
.C1(n_1609),
.C2(n_1616),
.Y(n_1747)
);

AOI221x1_ASAP7_75t_L g1748 ( 
.A1(n_1743),
.A2(n_1635),
.B1(n_1646),
.B2(n_1638),
.C(n_1636),
.Y(n_1748)
);

AOI222xp33_ASAP7_75t_L g1749 ( 
.A1(n_1737),
.A2(n_1560),
.B1(n_1609),
.B2(n_1614),
.C1(n_1616),
.C2(n_1573),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1738),
.A2(n_1609),
.B1(n_1614),
.B2(n_1616),
.C(n_1658),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1746),
.B(n_1744),
.Y(n_1751)
);

AOI31xp33_ASAP7_75t_L g1752 ( 
.A1(n_1750),
.A2(n_1740),
.A3(n_1741),
.B(n_1739),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1749),
.B(n_1740),
.C(n_1658),
.Y(n_1753)
);

OAI321xp33_ASAP7_75t_L g1754 ( 
.A1(n_1747),
.A2(n_1649),
.A3(n_1666),
.B1(n_1461),
.B2(n_1639),
.C(n_1625),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1748),
.A2(n_1649),
.B1(n_1666),
.B2(n_1629),
.C(n_1641),
.Y(n_1755)
);

AOI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1746),
.A2(n_1464),
.B(n_1505),
.C(n_1504),
.Y(n_1756)
);

NOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1752),
.B(n_1464),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1645),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1755),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1754),
.B(n_1464),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1753),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_L g1762 ( 
.A(n_1761),
.B(n_1756),
.C(n_1468),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1758),
.B(n_1625),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1757),
.B(n_1634),
.Y(n_1764)
);

AOI31xp33_ASAP7_75t_L g1765 ( 
.A1(n_1763),
.A2(n_1759),
.A3(n_1760),
.B(n_1435),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1764),
.B1(n_1762),
.B2(n_1646),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1629),
.B1(n_1641),
.B2(n_1638),
.Y(n_1767)
);

OAI22x1_ASAP7_75t_L g1768 ( 
.A1(n_1766),
.A2(n_1636),
.B1(n_1641),
.B2(n_1629),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1767),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1769),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1770),
.A2(n_1644),
.B(n_1594),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1771),
.Y(n_1773)
);

OA22x2_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1772),
.B1(n_1644),
.B2(n_1594),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1774),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1472),
.B1(n_1466),
.B2(n_1469),
.Y(n_1776)
);

AOI211xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1456),
.B(n_1459),
.C(n_1431),
.Y(n_1777)
);


endmodule