module fake_netlist_1_6231_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
INVxp67_ASAP7_75t_SL g12 ( .A(n_6), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx8_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NOR3xp33_ASAP7_75t_L g16 ( .A(n_10), .B(n_2), .C(n_3), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_17), .B(n_12), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_18), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g21 ( .A(n_20), .B(n_14), .Y(n_21) );
OAI21xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_13), .B(n_5), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_7), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
CKINVDCx20_ASAP7_75t_R g25 ( .A(n_24), .Y(n_25) );
OR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_9), .Y(n_26) );
endmodule