module fake_jpeg_20651_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

NAND2x1_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.C(n_18),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_8),
.C(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_29),
.B1(n_32),
.B2(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_16),
.B(n_28),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_37),
.B(n_40),
.C(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_41),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_48),
.B1(n_50),
.B2(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_43),
.B1(n_47),
.B2(n_7),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_5),
.C(n_6),
.Y(n_54)
);


endmodule