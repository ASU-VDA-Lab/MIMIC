module fake_jpeg_16224_n_45 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_28)
);

AOI221xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_23),
.C(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_36),
.C(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_7),
.C(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_13),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_14),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_41),
.Y(n_45)
);


endmodule