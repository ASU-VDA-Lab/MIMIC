module fake_jpeg_831_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx8_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_SL g8 ( 
.A(n_4),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp33_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_19),
.B(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_17),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_11),
.B1(n_9),
.B2(n_12),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_17),
.C(n_13),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_20),
.C(n_15),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_21),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_22),
.B1(n_20),
.B2(n_14),
.Y(n_28)
);

OAI221xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_30),
.B1(n_27),
.B2(n_15),
.C(n_14),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_23),
.C(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_9),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_29),
.C(n_12),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_3),
.Y(n_35)
);

AOI321xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_7),
.C(n_22),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_1),
.Y(n_37)
);


endmodule