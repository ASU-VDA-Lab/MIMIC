module fake_jpeg_19005_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_44),
.Y(n_64)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_30),
.B1(n_26),
.B2(n_28),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_30),
.B1(n_26),
.B2(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_31),
.Y(n_73)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_79),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_87),
.Y(n_113)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_64),
.B(n_27),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_90),
.B1(n_96),
.B2(n_36),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_39),
.B1(n_47),
.B2(n_49),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_75),
.B1(n_69),
.B2(n_82),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_44),
.C(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_44),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_45),
.B1(n_39),
.B2(n_47),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_97),
.B1(n_55),
.B2(n_60),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_37),
.B(n_36),
.C(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_34),
.B1(n_35),
.B2(n_25),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_55),
.B(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_59),
.Y(n_109)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_20),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_145)
);

NOR2x1p5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_38),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_127),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_123),
.B1(n_91),
.B2(n_37),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_72),
.B1(n_75),
.B2(n_99),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_133),
.B1(n_61),
.B2(n_53),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_35),
.B1(n_21),
.B2(n_25),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_21),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_48),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_48),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_132),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_38),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_93),
.B(n_63),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_20),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_93),
.C(n_89),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_105),
.C(n_110),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_20),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_139),
.B1(n_153),
.B2(n_157),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_80),
.B1(n_100),
.B2(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_150),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_23),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_117),
.B1(n_133),
.B2(n_118),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_109),
.B(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_118),
.B1(n_111),
.B2(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_158),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_23),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_115),
.Y(n_169)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_63),
.B1(n_76),
.B2(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_108),
.A2(n_74),
.B1(n_12),
.B2(n_14),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_61),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_107),
.B1(n_129),
.B2(n_102),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_163),
.A2(n_164),
.B1(n_175),
.B2(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_130),
.B1(n_127),
.B2(n_133),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_110),
.B1(n_131),
.B2(n_117),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_166),
.A2(n_29),
.B1(n_17),
.B2(n_33),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_185),
.B(n_154),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_192),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_155),
.B1(n_143),
.B2(n_147),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_172),
.A2(n_179),
.B1(n_7),
.B2(n_8),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_122),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_111),
.B1(n_124),
.B2(n_116),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_124),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_124),
.B1(n_116),
.B2(n_11),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_61),
.C(n_53),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_187),
.C(n_161),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_156),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_142),
.A2(n_53),
.B(n_29),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_135),
.A2(n_9),
.B1(n_11),
.B2(n_8),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_145),
.B1(n_156),
.B2(n_140),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_17),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_194),
.B(n_195),
.Y(n_235)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_198),
.Y(n_237)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx6p67_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_171),
.B(n_134),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g242 ( 
.A(n_200),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_160),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_214),
.B(n_224),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_163),
.B(n_20),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_216),
.B(n_218),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_144),
.C(n_32),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_210),
.C(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_192),
.B(n_165),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_32),
.Y(n_222)
);

OAI211xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_179),
.B(n_170),
.C(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_180),
.B(n_7),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_234),
.A2(n_202),
.B1(n_212),
.B2(n_211),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_164),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_247),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_162),
.C(n_189),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_162),
.B(n_17),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_221),
.B(n_193),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_33),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_198),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_32),
.C(n_24),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_24),
.C(n_18),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_218),
.A2(n_219),
.B1(n_216),
.B2(n_193),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_211),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_260),
.B1(n_234),
.B2(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_209),
.B(n_208),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_264),
.B(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_203),
.B1(n_213),
.B2(n_199),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_258),
.A2(n_265),
.B1(n_246),
.B2(n_229),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_197),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_240),
.B(n_6),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_270),
.B1(n_266),
.B2(n_250),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_199),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_228),
.B1(n_225),
.B2(n_243),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_199),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_0),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_267),
.C(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_287),
.C(n_289),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_232),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_259),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_236),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_33),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_247),
.C(n_249),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_242),
.C(n_230),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_251),
.C(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_297),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_258),
.C(n_260),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_284),
.C(n_285),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_255),
.C(n_268),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_1),
.Y(n_316)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_253),
.B1(n_262),
.B2(n_257),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_282),
.B1(n_281),
.B2(n_273),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_272),
.A2(n_270),
.B(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_5),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_287),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_306),
.A2(n_316),
.B(n_8),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_288),
.B(n_290),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_280),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_292),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_317),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_321),
.C(n_322),
.Y(n_333)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_303),
.B1(n_293),
.B2(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_323),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_312),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_325),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_296),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_18),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_309),
.CI(n_296),
.CON(n_330),
.SN(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_317),
.B(n_309),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_331),
.A2(n_4),
.B(n_2),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_333),
.A2(n_18),
.B1(n_24),
.B2(n_4),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_4),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_336),
.B(n_1),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_332),
.B1(n_329),
.B2(n_328),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_339),
.B(n_334),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_330),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_1),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_1),
.B(n_2),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_3),
.C(n_279),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_3),
.B(n_343),
.Y(n_346)
);


endmodule