module real_jpeg_23077_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_286;
wire n_288;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_1),
.A2(n_73),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_132),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_132),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_8),
.A2(n_64),
.B1(n_71),
.B2(n_73),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_191)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_10),
.A2(n_70),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_10),
.A2(n_59),
.B1(n_60),
.B2(n_85),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_85),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_85),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_11),
.B(n_133),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_80),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_42),
.C(n_56),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_11),
.B(n_153),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_182),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_28),
.C(n_47),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_11),
.A2(n_30),
.B(n_241),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_12),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_69),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_69),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_15),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_122)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_20),
.B(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_86),
.B2(n_112),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.C(n_66),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_23),
.A2(n_24),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_25),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_26),
.A2(n_30),
.B1(n_101),
.B2(n_121),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_27),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_30),
.A2(n_32),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_30),
.A2(n_161),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_30),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_30),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_31),
.Y(n_164)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_31),
.Y(n_242)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_35),
.A2(n_159),
.B1(n_253),
.B2(n_255),
.Y(n_252)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_36),
.B(n_182),
.Y(n_265)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_40),
.A2(n_49),
.B1(n_92),
.B2(n_124),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_42),
.B(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_50),
.B1(n_52),
.B2(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_45),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_45),
.A2(n_52),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_49),
.A2(n_124),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_49),
.A2(n_178),
.B(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_49),
.B(n_182),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_52),
.B(n_179),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_53),
.B(n_66),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_55),
.B1(n_65),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_54),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_54),
.A2(n_152),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_63),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_55),
.A2(n_127),
.B(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_60),
.B1(n_77),
.B2(n_78),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_59),
.A2(n_78),
.A3(n_134),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_60),
.B(n_77),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_60),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_74),
.B(n_81),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_75),
.B1(n_80),
.B2(n_131),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_71),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_75),
.A2(n_82),
.B(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_79),
.A2(n_110),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_97),
.B2(n_98),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_96),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_92),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_92),
.A2(n_229),
.B(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_117)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_125),
.C(n_130),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_123),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_151),
.B1(n_153),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_289),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_165),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_139),
.B(n_165),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_144),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_146),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_154),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_149),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_199),
.B(n_283),
.C(n_288),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_193),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.C(n_185),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_170),
.A2(n_171),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_184),
.B(n_185),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_192),
.A2(n_254),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_194),
.B(n_197),
.C(n_198),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_277),
.B(n_282),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_230),
.B(n_276),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_219),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_204),
.B(n_219),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.C(n_216),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_205),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_212),
.A2(n_216),
.B1(n_217),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_226),
.C(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_270),
.B(n_275),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_250),
.B(n_269),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_244),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_244),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_246),
.B1(n_248),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_248),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_258),
.B(n_268),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_256),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_263),
.B(n_267),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_281),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);


endmodule