module fake_jpeg_22814_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_46),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_50),
.B(n_26),
.C(n_27),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_28),
.B1(n_23),
.B2(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_28),
.B1(n_82),
.B2(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_59),
.A2(n_64),
.B1(n_71),
.B2(n_79),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_69),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_36),
.B1(n_39),
.B2(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_77),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_24),
.B(n_31),
.Y(n_103)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_50),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_99),
.B1(n_101),
.B2(n_108),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_50),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_37),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_18),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_66),
.B(n_18),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_2),
.B(n_3),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_51),
.C(n_18),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_22),
.C(n_34),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_28),
.B1(n_19),
.B2(n_37),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_1),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_120),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_37),
.B1(n_19),
.B2(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_111),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_65),
.A2(n_19),
.B1(n_31),
.B2(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_34),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_5),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_25),
.B1(n_21),
.B2(n_33),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_34),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_34),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_2),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_129),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_128),
.Y(n_160)
);

AO22x2_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_67),
.B1(n_83),
.B2(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_119),
.B1(n_98),
.B2(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_130),
.B(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_30),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_119),
.A2(n_67),
.B1(n_21),
.B2(n_30),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_87),
.B1(n_104),
.B2(n_110),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_22),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_137),
.B(n_140),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_139),
.B(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_159),
.B1(n_117),
.B2(n_131),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_103),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_148),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_150),
.Y(n_174)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_151),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_87),
.Y(n_152)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_120),
.B1(n_121),
.B2(n_100),
.Y(n_159)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_94),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_170),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_173),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_193),
.B1(n_191),
.B2(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_91),
.B1(n_121),
.B2(n_123),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_183),
.B1(n_186),
.B2(n_138),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_95),
.B(n_104),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_100),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_120),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_185),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_112),
.B1(n_95),
.B2(n_102),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_112),
.B(n_102),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_143),
.B(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_89),
.B1(n_7),
.B2(n_9),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_6),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_193),
.Y(n_210)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_136),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_127),
.B(n_139),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_194),
.A2(n_204),
.B(n_215),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_196),
.B1(n_200),
.B2(n_214),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_173),
.A2(n_127),
.B1(n_147),
.B2(n_156),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_129),
.B1(n_130),
.B2(n_158),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_202),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_203),
.A2(n_163),
.B1(n_166),
.B2(n_12),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_156),
.B(n_140),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_161),
.A2(n_149),
.B1(n_148),
.B2(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_185),
.A3(n_183),
.B1(n_181),
.B2(n_186),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_195),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_7),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_196),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_227),
.B(n_209),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_189),
.B1(n_163),
.B2(n_188),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_228),
.A2(n_247),
.B1(n_199),
.B2(n_208),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_222),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_232),
.B(n_235),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_169),
.C(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_201),
.C(n_11),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_194),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_192),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_206),
.C(n_202),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_169),
.B1(n_188),
.B2(n_164),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_203),
.B1(n_207),
.B2(n_219),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_235),
.B1(n_241),
.B2(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_166),
.B1(n_11),
.B2(n_13),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_251),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_260),
.B1(n_261),
.B2(n_246),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_258),
.C(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_253),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_228),
.B(n_211),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_254),
.A2(n_255),
.B(n_234),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_212),
.B(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_262),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_204),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_206),
.B1(n_218),
.B2(n_205),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_216),
.C(n_223),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.C(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_231),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_237),
.B(n_224),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_270),
.B(n_279),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_278),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_238),
.B1(n_241),
.B2(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_280),
.B1(n_283),
.B2(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_234),
.B(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_249),
.A2(n_230),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_259),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_229),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_289),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_242),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_291),
.B(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_295),
.C(n_297),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_282),
.C(n_271),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_258),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_253),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_283),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_273),
.B1(n_278),
.B2(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_269),
.B(n_272),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_297),
.B(n_288),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_275),
.B1(n_276),
.B2(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_298),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_309),
.A2(n_296),
.B1(n_287),
.B2(n_293),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_13),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_320),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_300),
.C(n_308),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_321),
.C(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_312),
.C(n_318),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_322),
.B(n_315),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_313),
.B(n_304),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_15),
.B(n_16),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_16),
.Y(n_332)
);


endmodule