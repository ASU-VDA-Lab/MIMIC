module fake_jpeg_21230_n_290 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_31),
.C(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_29),
.B(n_23),
.C(n_24),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_26),
.B(n_30),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_9),
.C(n_12),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_31),
.B1(n_25),
.B2(n_13),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_60),
.B1(n_28),
.B2(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_28),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_44),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_25),
.B1(n_13),
.B2(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_45),
.B1(n_41),
.B2(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_57),
.B1(n_60),
.B2(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_46),
.B1(n_38),
.B2(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_69),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_70),
.A2(n_81),
.B1(n_102),
.B2(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_76),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_19),
.B(n_30),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_73),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_14),
.A3(n_26),
.B1(n_19),
.B2(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_14),
.B1(n_20),
.B2(n_16),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_79),
.B(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_14),
.B1(n_20),
.B2(n_16),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_15),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_27),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_22),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_96),
.B1(n_0),
.B2(n_1),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_17),
.B1(n_15),
.B2(n_29),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_3),
.B(n_4),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_44),
.C(n_37),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_36),
.C(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_36),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_36),
.B1(n_44),
.B2(n_9),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_12),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_111),
.B1(n_112),
.B2(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_110),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_43),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_43),
.B1(n_22),
.B2(n_3),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_137),
.B(n_79),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_12),
.C(n_11),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_88),
.B1(n_77),
.B2(n_90),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_72),
.B1(n_71),
.B2(n_76),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_83),
.A2(n_4),
.B(n_5),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_119),
.B1(n_115),
.B2(n_126),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_95),
.B1(n_82),
.B2(n_66),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_158),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_64),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_149),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_116),
.B(n_133),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_148),
.B(n_157),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_70),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_116),
.B1(n_124),
.B2(n_128),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_159),
.B1(n_105),
.B2(n_109),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_75),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_93),
.Y(n_156)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_102),
.B1(n_78),
.B2(n_7),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_10),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_118),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_111),
.B1(n_106),
.B2(n_135),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_172),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_115),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_107),
.C(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_171),
.B(n_175),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_179),
.B1(n_187),
.B2(n_158),
.Y(n_198)
);

BUFx4f_ASAP7_75t_SL g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_176),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_110),
.C(n_108),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_139),
.C(n_153),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_109),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_162),
.B1(n_151),
.B2(n_154),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_188),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_144),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_194),
.C(n_205),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_211),
.B1(n_186),
.B2(n_185),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_179),
.B(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_154),
.A3(n_141),
.B1(n_147),
.B2(n_148),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_212),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_160),
.C(n_132),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_172),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_183),
.A2(n_159),
.B1(n_147),
.B2(n_121),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_222),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_174),
.B(n_167),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_226),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_224),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_169),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_182),
.C(n_184),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_205),
.C(n_207),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_201),
.B1(n_196),
.B2(n_163),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_174),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_230),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_197),
.C(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_247),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_190),
.B1(n_200),
.B2(n_212),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_243),
.B1(n_214),
.B2(n_228),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_229),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_190),
.B1(n_206),
.B2(n_208),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_225),
.B1(n_224),
.B2(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_119),
.C(n_196),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_231),
.A2(n_163),
.B1(n_180),
.B2(n_176),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_217),
.B1(n_216),
.B2(n_232),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_256),
.Y(n_262)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_222),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_215),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_126),
.B1(n_130),
.B2(n_104),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_248),
.C(n_235),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_239),
.B(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_243),
.B(n_245),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_247),
.C(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_254),
.C(n_233),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_263),
.B1(n_268),
.B2(n_250),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.C(n_265),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_249),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_265),
.B(n_6),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_251),
.B1(n_269),
.B2(n_238),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_104),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_276),
.A2(n_273),
.B1(n_275),
.B2(n_130),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_104),
.B1(n_7),
.B2(n_8),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_285),
.B1(n_280),
.B2(n_281),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_282),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.C(n_284),
.Y(n_288)
);

AOI31xp67_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_5),
.A3(n_7),
.B(n_8),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_5),
.Y(n_290)
);


endmodule