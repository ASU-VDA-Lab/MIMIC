module fake_jpeg_22478_n_307 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_43),
.Y(n_50)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_21),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_61),
.B1(n_46),
.B2(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_20),
.B1(n_19),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_69),
.B1(n_70),
.B2(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_74),
.B1(n_34),
.B2(n_33),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_36),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_31),
.B1(n_26),
.B2(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_46),
.Y(n_85)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_27),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_22),
.B1(n_23),
.B2(n_34),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_40),
.B1(n_37),
.B2(n_45),
.Y(n_75)
);

OA22x2_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_40),
.A2(n_43),
.B1(n_39),
.B2(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_35),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.C(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_32),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_43),
.C(n_44),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_83),
.B(n_112),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_28),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_99),
.B1(n_101),
.B2(n_117),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_62),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_97),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_34),
.B1(n_33),
.B2(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_102),
.Y(n_139)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_60),
.B(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_33),
.B1(n_30),
.B2(n_21),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_53),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_51),
.A2(n_30),
.B1(n_22),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_60),
.B1(n_74),
.B2(n_61),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_118),
.A2(n_144),
.B1(n_149),
.B2(n_107),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_53),
.B1(n_71),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_119),
.A2(n_150),
.B1(n_104),
.B2(n_116),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_67),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_131),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_50),
.B(n_77),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_82),
.B(n_75),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_50),
.B(n_65),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_105),
.B(n_75),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_106),
.B1(n_113),
.B2(n_96),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_64),
.B1(n_58),
.B2(n_75),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_70),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_76),
.B(n_75),
.C(n_78),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_75),
.B1(n_55),
.B2(n_71),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_152),
.B(n_171),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_141),
.B1(n_146),
.B2(n_150),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_178),
.B1(n_146),
.B2(n_118),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_81),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_163),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_162),
.B(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_105),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_0),
.Y(n_165)
);

AOI21x1_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_174),
.B(n_3),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_93),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_182),
.B1(n_121),
.B2(n_122),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_130),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_175),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_55),
.B1(n_90),
.B2(n_100),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_98),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_94),
.C(n_92),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_1),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_1),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_98),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_104),
.C(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_127),
.B(n_1),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_97),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2x1p5_ASAP7_75t_R g182 ( 
.A(n_149),
.B(n_3),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_187),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_193),
.B(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_126),
.B1(n_133),
.B2(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_145),
.B(n_125),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_119),
.B1(n_121),
.B2(n_128),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_207),
.B(n_165),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_122),
.B(n_123),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_138),
.B1(n_132),
.B2(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

AOI22x1_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_132),
.B1(n_135),
.B2(n_5),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_154),
.B(n_155),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_120),
.B1(n_5),
.B2(n_6),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_152),
.B1(n_174),
.B2(n_161),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_163),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_203),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_169),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_217),
.C(n_226),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_153),
.C(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

NAND5xp2_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_176),
.C(n_165),
.D(n_168),
.E(n_177),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_198),
.B(n_189),
.Y(n_248)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_180),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_181),
.C(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_232),
.C(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_4),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_229),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_233),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_17),
.C(n_8),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_4),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_207),
.C(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_188),
.B1(n_191),
.B2(n_184),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_231),
.B1(n_222),
.B2(n_219),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_201),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_240),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_222),
.B(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_200),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_250),
.B1(n_225),
.B2(n_219),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_184),
.B1(n_190),
.B2(n_205),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_249),
.B1(n_218),
.B2(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_217),
.C(n_226),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_221),
.C(n_216),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_198),
.B1(n_186),
.B2(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.C(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_261),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_212),
.C(n_224),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_260),
.B(n_262),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_237),
.B(n_251),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_235),
.A2(n_225),
.B1(n_227),
.B2(n_213),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_213),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_220),
.B1(n_216),
.B2(n_206),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_237),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_197),
.C(n_10),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_246),
.C(n_236),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_277),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_248),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_249),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_240),
.C(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_261),
.C(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_282),
.C(n_264),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_286),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_256),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_259),
.B(n_254),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_292),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_285),
.A2(n_274),
.B1(n_273),
.B2(n_258),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_290),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_14),
.C(n_15),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_281),
.A2(n_274),
.B1(n_262),
.B2(n_257),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_271),
.C(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_282),
.C(n_11),
.Y(n_295)
);

AOI31xp67_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_197),
.A3(n_245),
.B(n_12),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_12),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_299),
.C(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_300),
.B(n_302),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_293),
.A3(n_291),
.B1(n_16),
.B2(n_17),
.C1(n_15),
.C2(n_14),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_295),
.B(n_14),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_17),
.Y(n_307)
);


endmodule