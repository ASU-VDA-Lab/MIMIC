module fake_jpeg_16181_n_29 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

INVx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_18),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_11),
.C(n_10),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_18),
.B(n_11),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_9),
.B1(n_6),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_14),
.B1(n_12),
.B2(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_16),
.C(n_15),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_21),
.A2(n_22),
.B1(n_12),
.B2(n_1),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

AOI31xp67_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_2),
.A3(n_4),
.B(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_4),
.B1(n_5),
.B2(n_23),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_22),
.B(n_26),
.Y(n_29)
);


endmodule