module fake_ibex_20_n_1801 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_105, n_187, n_1, n_154, n_182, n_196, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_57, n_301, n_296, n_120, n_168, n_155, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_55, n_291, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1801);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_55;
input n_291;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1801;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_1782;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_1778;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_324;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1599;
wire n_712;
wire n_1400;
wire n_1539;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_344;
wire n_436;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_326;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_339;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_360;
wire n_1770;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_336;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1755;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_319;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx2_ASAP7_75t_L g315 ( 
.A(n_50),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_109),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_38),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_127),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_14),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_207),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_117),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_34),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_91),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_127),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_179),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_162),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_279),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_210),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_70),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_56),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_80),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_145),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_239),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_63),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_124),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_47),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_133),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_86),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_63),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_267),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_23),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_60),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_58),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_185),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_133),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_222),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_147),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_270),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_309),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_212),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_28),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_160),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_197),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g363 ( 
.A(n_148),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_66),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_271),
.B(n_199),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_247),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_45),
.B(n_32),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_194),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_242),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_57),
.B(n_45),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_57),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_38),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_62),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_293),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_47),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_273),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_64),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_167),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_72),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_287),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_230),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_84),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_250),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_150),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_53),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_276),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_48),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_13),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_129),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g392 ( 
.A(n_204),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_89),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_296),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_166),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_70),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_111),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_155),
.B(n_181),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_178),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_251),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_219),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_78),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_189),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_265),
.B(n_235),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_95),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_13),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_196),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_255),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_225),
.B(n_254),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_62),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_19),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_191),
.Y(n_412)
);

BUFx8_ASAP7_75t_SL g413 ( 
.A(n_126),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_137),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_217),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_83),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_131),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_310),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_123),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_139),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_232),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_31),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_277),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_244),
.B(n_143),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_311),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_195),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_186),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_17),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_307),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_153),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_165),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_266),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_93),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_182),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_123),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_215),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_248),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_313),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_253),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_231),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_154),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_252),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_301),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_240),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_29),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_180),
.B(n_205),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_245),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_100),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_268),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_216),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_183),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_49),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_224),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_314),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_43),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_297),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_234),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_141),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_211),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_289),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_46),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_128),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_274),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_5),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_159),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_236),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_229),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_294),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_258),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_227),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_228),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_203),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_202),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_33),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_74),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_288),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_263),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_303),
.Y(n_478)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_187),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_176),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_243),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_308),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_122),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_4),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_142),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_171),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_65),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_124),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_43),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_169),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_115),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_305),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_52),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_53),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_113),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_298),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_161),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_291),
.B(n_104),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_249),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_264),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_72),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_172),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_221),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_95),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_142),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_295),
.B(n_81),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_102),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_233),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_84),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_156),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_119),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_281),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_104),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_256),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_93),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_79),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_201),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_105),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_90),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_290),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_67),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_23),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_220),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_3),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_44),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_168),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_163),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_116),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_12),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_75),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_113),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_42),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_173),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_226),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_164),
.Y(n_535)
);

INVx4_ASAP7_75t_R g536 ( 
.A(n_121),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_7),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_77),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_135),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_260),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_51),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_261),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_333),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_392),
.B(n_0),
.Y(n_544)
);

BUFx12f_ASAP7_75t_L g545 ( 
.A(n_333),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_487),
.B(n_0),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g547 ( 
.A1(n_323),
.A2(n_146),
.B(n_144),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_333),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_363),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_363),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_363),
.Y(n_552)
);

OAI22x1_ASAP7_75t_L g553 ( 
.A1(n_334),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_363),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_363),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_321),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_421),
.B(n_1),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_331),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_2),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_331),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_4),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_363),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_315),
.B(n_319),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_315),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_319),
.Y(n_567)
);

CKINVDCx6p67_ASAP7_75t_R g568 ( 
.A(n_425),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_328),
.B(n_5),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_331),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_331),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_410),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_392),
.B(n_6),
.Y(n_574)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_355),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_363),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_321),
.B(n_6),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_353),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_477),
.Y(n_580)
);

BUFx12f_ASAP7_75t_L g581 ( 
.A(n_527),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_323),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_358),
.B(n_149),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_435),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_358),
.Y(n_585)
);

OAI22x1_ASAP7_75t_L g586 ( 
.A1(n_334),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_355),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_449),
.Y(n_589)
);

NOR2x1_ASAP7_75t_L g590 ( 
.A(n_485),
.B(n_151),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_385),
.B(n_152),
.Y(n_591)
);

OAI22x1_ASAP7_75t_R g592 ( 
.A1(n_364),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_353),
.B(n_525),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_385),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_526),
.B(n_10),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_336),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_525),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_355),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

CKINVDCx11_ASAP7_75t_R g601 ( 
.A(n_364),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_336),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_436),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_375),
.B(n_470),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_355),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_436),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_316),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_318),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_369),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_369),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_369),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_413),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_322),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_354),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_453),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_354),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_371),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_317),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_369),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_394),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_394),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_394),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_394),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_329),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_368),
.Y(n_625)
);

INVx6_ASAP7_75t_L g626 ( 
.A(n_423),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_473),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_423),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_368),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_356),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_335),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_362),
.B(n_15),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_379),
.A2(n_158),
.B(n_157),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_326),
.B(n_15),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_423),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_366),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_335),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_379),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_479),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_423),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_454),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_470),
.B(n_18),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_371),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_519),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_546),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_549),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g648 ( 
.A(n_631),
.B(n_519),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_550),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_568),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_546),
.Y(n_651)
);

NOR2x1p5_ASAP7_75t_L g652 ( 
.A(n_631),
.B(n_522),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_593),
.B(n_579),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_546),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_550),
.Y(n_655)
);

CKINVDCx6p67_ASAP7_75t_R g656 ( 
.A(n_568),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_615),
.A2(n_522),
.B1(n_387),
.B2(n_406),
.Y(n_657)
);

AND3x2_ASAP7_75t_L g658 ( 
.A(n_644),
.B(n_420),
.C(n_411),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_552),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_644),
.B(n_458),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_552),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_548),
.B(n_437),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_560),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_548),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_548),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_R g668 ( 
.A1(n_558),
.A2(n_521),
.B1(n_396),
.B2(n_324),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

BUFx6f_ASAP7_75t_SL g670 ( 
.A(n_562),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_604),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_579),
.B(n_479),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_563),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_575),
.B(n_490),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_575),
.B(n_374),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_575),
.B(n_320),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_575),
.B(n_376),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_598),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_580),
.B(n_377),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_580),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_580),
.B(n_327),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_577),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_580),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_582),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_642),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_604),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_559),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_559),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_559),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_544),
.B(n_351),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_583),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_562),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_589),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_612),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_559),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_639),
.A2(n_387),
.B1(n_406),
.B2(n_383),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_642),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_562),
.Y(n_698)
);

AOI21x1_ASAP7_75t_L g699 ( 
.A1(n_633),
.A2(n_590),
.B(n_607),
.Y(n_699)
);

AND3x2_ASAP7_75t_L g700 ( 
.A(n_637),
.B(n_413),
.C(n_340),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_570),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_551),
.Y(n_704)
);

CKINVDCx6p67_ASAP7_75t_R g705 ( 
.A(n_543),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_SL g706 ( 
.A1(n_595),
.A2(n_341),
.B1(n_343),
.B2(n_337),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_612),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_578),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_544),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_543),
.B(n_381),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_570),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_545),
.B(n_564),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_582),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_574),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_574),
.B(n_351),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_545),
.B(n_384),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_565),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_591),
.B(n_454),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_564),
.B(n_386),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_570),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_572),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_581),
.B(n_403),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_578),
.B(n_351),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_572),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_SL g725 ( 
.A(n_591),
.B(n_347),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_569),
.B(n_344),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_556),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_581),
.B(n_408),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_572),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_572),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_608),
.B(n_332),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_572),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_565),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_613),
.B(n_338),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_576),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_613),
.B(n_624),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_565),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_585),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_630),
.B(n_636),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_576),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_630),
.B(n_346),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_556),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_576),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_605),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_636),
.B(n_367),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_596),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

AO21x2_ASAP7_75t_L g750 ( 
.A1(n_633),
.A2(n_424),
.B(n_330),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_605),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_605),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_609),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_602),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_609),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_614),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_618),
.B(n_342),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_601),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_614),
.Y(n_759)
);

INVxp33_ASAP7_75t_L g760 ( 
.A(n_634),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_609),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_609),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_611),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_594),
.Y(n_764)
);

INVxp33_ASAP7_75t_SL g765 ( 
.A(n_553),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_603),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_611),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_611),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_573),
.B(n_588),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_616),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_611),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_616),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_573),
.B(n_350),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_619),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_619),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_603),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_547),
.A2(n_520),
.B(n_441),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_625),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_606),
.B(n_352),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_619),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_627),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_629),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_619),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_619),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_629),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_622),
.Y(n_786)
);

BUFx2_ASAP7_75t_L g787 ( 
.A(n_627),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_573),
.B(n_397),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_638),
.B(n_357),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_638),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_588),
.B(n_434),
.Y(n_791)
);

AO21x2_ASAP7_75t_L g792 ( 
.A1(n_557),
.A2(n_442),
.B(n_439),
.Y(n_792)
);

OA22x2_ASAP7_75t_L g793 ( 
.A1(n_553),
.A2(n_345),
.B1(n_349),
.B2(n_325),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_561),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_588),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_597),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_622),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_597),
.B(n_360),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_622),
.Y(n_799)
);

AND2x6_ASAP7_75t_L g800 ( 
.A(n_632),
.B(n_473),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_566),
.B(n_361),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_561),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_622),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_769),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_657),
.B(n_696),
.C(n_706),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_693),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_795),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_691),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_678),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_760),
.B(n_690),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_660),
.B(n_600),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_769),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_715),
.B(n_600),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_715),
.B(n_788),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_788),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_676),
.B(n_567),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_681),
.B(n_567),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_737),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_790),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_795),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_790),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_787),
.B(n_571),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_712),
.B(n_586),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_717),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_723),
.B(n_397),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_734),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_738),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_678),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_584),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_714),
.B(n_584),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_702),
.Y(n_831)
);

INVx4_ASAP7_75t_L g832 ( 
.A(n_670),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_703),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_672),
.B(n_339),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_781),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_725),
.B(n_390),
.C(n_373),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_742),
.B(n_399),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_704),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_685),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_693),
.B(n_400),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_723),
.B(n_685),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_693),
.B(n_444),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_697),
.B(n_401),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_773),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_697),
.B(n_407),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_671),
.A2(n_382),
.B1(n_388),
.B2(n_347),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_739),
.B(n_708),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_793),
.A2(n_586),
.B1(n_380),
.B2(n_389),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_731),
.B(n_447),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_708),
.Y(n_850)
);

AOI22x1_ASAP7_75t_SL g851 ( 
.A1(n_650),
.A2(n_484),
.B1(n_537),
.B2(n_383),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_726),
.B(n_412),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_726),
.B(n_402),
.C(n_391),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_735),
.B(n_456),
.Y(n_854)
);

INVxp67_ASAP7_75t_SL g855 ( 
.A(n_664),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_662),
.B(n_476),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_660),
.B(n_397),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_675),
.B(n_426),
.Y(n_858)
);

AND3x1_ASAP7_75t_L g859 ( 
.A(n_722),
.B(n_592),
.C(n_393),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_757),
.B(n_478),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_683),
.B(n_427),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_677),
.B(n_429),
.Y(n_862)
);

NOR2x1p5_ASAP7_75t_L g863 ( 
.A(n_705),
.B(n_405),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_796),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_683),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_800),
.B(n_646),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_679),
.B(n_430),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_653),
.B(n_348),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_674),
.B(n_431),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_705),
.B(n_417),
.Y(n_870)
);

NOR2xp67_ASAP7_75t_L g871 ( 
.A(n_650),
.B(n_409),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_651),
.B(n_432),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_683),
.B(n_438),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_686),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_654),
.B(n_443),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_766),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_684),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_656),
.B(n_422),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_713),
.Y(n_879)
);

NAND2x1p5_ASAP7_75t_L g880 ( 
.A(n_664),
.B(n_378),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_698),
.A2(n_382),
.B1(n_395),
.B2(n_388),
.Y(n_881)
);

BUFx6f_ASAP7_75t_SL g882 ( 
.A(n_758),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_798),
.B(n_451),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_665),
.Y(n_884)
);

NOR2x1_ASAP7_75t_L g885 ( 
.A(n_648),
.B(n_395),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_776),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_801),
.B(n_480),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_789),
.B(n_481),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_793),
.A2(n_416),
.B1(n_419),
.B2(n_414),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_692),
.A2(n_433),
.B(n_445),
.C(n_428),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_749),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_749),
.Y(n_892)
);

OAI221xp5_ASAP7_75t_L g893 ( 
.A1(n_728),
.A2(n_448),
.B1(n_489),
.B2(n_488),
.C(n_483),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_710),
.B(n_457),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_716),
.B(n_459),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_754),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_740),
.B(n_460),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_670),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_719),
.B(n_455),
.C(n_452),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_692),
.B(n_776),
.Y(n_901)
);

INVx1_ASAP7_75t_SL g902 ( 
.A(n_656),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_692),
.B(n_466),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_666),
.B(n_468),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_756),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_652),
.B(n_461),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_680),
.B(n_469),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_680),
.B(n_800),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_800),
.B(n_471),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_759),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_800),
.B(n_472),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_770),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_694),
.B(n_707),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_747),
.B(n_496),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_779),
.B(n_486),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_747),
.B(n_497),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_747),
.B(n_492),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_SL g918 ( 
.A1(n_765),
.A2(n_537),
.B1(n_484),
.B2(n_727),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_792),
.B(n_500),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_746),
.B(n_503),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_793),
.A2(n_504),
.B1(n_505),
.B2(n_493),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_764),
.B(n_510),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_668),
.A2(n_415),
.B1(n_450),
.B2(n_418),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_764),
.B(n_514),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_792),
.B(n_512),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_694),
.B(n_462),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_792),
.B(n_517),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_748),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_772),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_791),
.B(n_474),
.C(n_464),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_778),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_658),
.B(n_535),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_707),
.B(n_475),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_673),
.B(n_540),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_673),
.B(n_542),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_645),
.B(n_523),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_L g937 ( 
.A(n_668),
.B(n_495),
.C(n_494),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_782),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_785),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_699),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_718),
.B(n_359),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_758),
.B(n_501),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_647),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_727),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_699),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_700),
.B(n_513),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_649),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_655),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_794),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_765),
.A2(n_509),
.B1(n_511),
.B2(n_507),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_659),
.B(n_482),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_659),
.B(n_502),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_661),
.B(n_508),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_663),
.A2(n_516),
.B(n_532),
.C(n_531),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_743),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_667),
.B(n_541),
.Y(n_956)
);

OAI22xp33_ASAP7_75t_L g957 ( 
.A1(n_743),
.A2(n_418),
.B1(n_450),
.B2(n_415),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_669),
.B(n_515),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_682),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_682),
.B(n_524),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_777),
.B(n_372),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_750),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_750),
.B(n_528),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_794),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_750),
.B(n_441),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_802),
.B(n_529),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_SL g967 ( 
.A(n_802),
.B(n_463),
.Y(n_967)
);

BUFx5_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_687),
.B(n_370),
.Y(n_969)
);

AO221x1_ASAP7_75t_L g970 ( 
.A1(n_786),
.A2(n_465),
.B1(n_463),
.B2(n_518),
.C(n_372),
.Y(n_970)
);

INVx8_ASAP7_75t_L g971 ( 
.A(n_786),
.Y(n_971)
);

OAI221xp5_ASAP7_75t_L g972 ( 
.A1(n_688),
.A2(n_538),
.B1(n_530),
.B2(n_506),
.C(n_498),
.Y(n_972)
);

BUFx8_ASAP7_75t_L g973 ( 
.A(n_786),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_803),
.B(n_534),
.C(n_520),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_689),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_689),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_799),
.B(n_533),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_961),
.A2(n_547),
.B(n_534),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_940),
.A2(n_547),
.B(n_695),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_919),
.A2(n_398),
.B(n_404),
.C(n_365),
.Y(n_980)
);

AOI33xp33_ASAP7_75t_L g981 ( 
.A1(n_950),
.A2(n_536),
.A3(n_784),
.B1(n_783),
.B2(n_780),
.B3(n_775),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_814),
.A2(n_643),
.B(n_617),
.C(n_533),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_945),
.A2(n_547),
.B(n_695),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_866),
.A2(n_711),
.B(n_701),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_828),
.B(n_518),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_881),
.B(n_19),
.Y(n_986)
);

BUFx4f_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_809),
.B(n_446),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_810),
.B(n_20),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_857),
.B(n_20),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_832),
.Y(n_991)
);

OR2x2_ASAP7_75t_SL g992 ( 
.A(n_957),
.B(n_467),
.Y(n_992)
);

BUFx3_ASAP7_75t_L g993 ( 
.A(n_973),
.Y(n_993)
);

O2A1O1Ixp5_ASAP7_75t_L g994 ( 
.A1(n_856),
.A2(n_797),
.B(n_721),
.C(n_724),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_844),
.B(n_21),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_919),
.A2(n_729),
.B(n_720),
.Y(n_996)
);

AOI33xp33_ASAP7_75t_L g997 ( 
.A1(n_950),
.A2(n_797),
.A3(n_784),
.B1(n_783),
.B2(n_780),
.B3(n_775),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_825),
.A2(n_626),
.B1(n_499),
.B2(n_467),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_855),
.A2(n_732),
.B(n_730),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_938),
.A2(n_626),
.B1(n_499),
.B2(n_467),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

AO21x1_ASAP7_75t_L g1002 ( 
.A1(n_925),
.A2(n_736),
.B(n_733),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_839),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_925),
.A2(n_741),
.B(n_736),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_930),
.A2(n_626),
.B1(n_499),
.B2(n_587),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_815),
.B(n_21),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_823),
.B(n_22),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_829),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_830),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_882),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_963),
.A2(n_745),
.B(n_744),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_973),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_957),
.B(n_751),
.C(n_745),
.Y(n_1013)
);

CKINVDCx14_ASAP7_75t_R g1014 ( 
.A(n_918),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_842),
.B(n_24),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_938),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_899),
.B(n_896),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_842),
.B(n_25),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_874),
.B(n_25),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_927),
.A2(n_753),
.B(n_752),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_901),
.A2(n_755),
.B(n_753),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_850),
.B(n_26),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_841),
.B(n_26),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_896),
.B(n_561),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_967),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_811),
.B(n_27),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_813),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_870),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_908),
.A2(n_762),
.B(n_761),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_852),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_816),
.A2(n_763),
.B(n_762),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_819),
.B(n_29),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_821),
.B(n_30),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_817),
.A2(n_768),
.B(n_767),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_30),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_903),
.A2(n_774),
.B(n_771),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_964),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_930),
.A2(n_587),
.B1(n_599),
.B2(n_561),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_808),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_880),
.B(n_31),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_900),
.A2(n_599),
.B1(n_610),
.B2(n_587),
.Y(n_1041)
);

AO21x1_ASAP7_75t_L g1042 ( 
.A1(n_974),
.A2(n_774),
.B(n_628),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_880),
.B(n_32),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_807),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_807),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_948),
.A2(n_599),
.B(n_587),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_944),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_882),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_920),
.A2(n_620),
.B(n_610),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_914),
.B(n_35),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_916),
.B(n_36),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_926),
.B(n_37),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_922),
.A2(n_620),
.B(n_610),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_924),
.A2(n_621),
.B(n_620),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_822),
.B(n_37),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_909),
.A2(n_621),
.B(n_623),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_911),
.A2(n_621),
.B(n_623),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_824),
.B(n_39),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_851),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_826),
.B(n_39),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_827),
.B(n_40),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_804),
.B(n_812),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_856),
.B(n_40),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_831),
.Y(n_1064)
);

AO21x2_ASAP7_75t_L g1065 ( 
.A1(n_970),
.A2(n_640),
.B(n_635),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_902),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_872),
.A2(n_640),
.B(n_635),
.Y(n_1067)
);

BUFx4f_ASAP7_75t_L g1068 ( 
.A(n_942),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_917),
.B(n_41),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_917),
.B(n_41),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_875),
.A2(n_641),
.B(n_640),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_820),
.Y(n_1072)
);

OAI321xp33_ASAP7_75t_L g1073 ( 
.A1(n_893),
.A2(n_641),
.A3(n_42),
.B1(n_44),
.B2(n_46),
.C(n_48),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_923),
.B(n_49),
.Y(n_1074)
);

CKINVDCx10_ASAP7_75t_R g1075 ( 
.A(n_859),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_889),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_974),
.A2(n_54),
.B(n_55),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_933),
.B(n_56),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_906),
.B(n_58),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_L g1080 ( 
.A(n_937),
.B(n_805),
.C(n_955),
.Y(n_1080)
);

AOI211xp5_ASAP7_75t_L g1081 ( 
.A1(n_937),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_878),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_805),
.B(n_68),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_849),
.B(n_69),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_849),
.B(n_69),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_854),
.B(n_71),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_860),
.B(n_73),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_860),
.B(n_73),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_837),
.A2(n_175),
.B(n_170),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_913),
.B(n_74),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_887),
.B(n_75),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_887),
.B(n_76),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_877),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_1093)
);

OAI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_958),
.A2(n_79),
.B(n_80),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_863),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_879),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_871),
.B(n_85),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_833),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_928),
.B(n_87),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_865),
.B(n_87),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_915),
.B(n_88),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_836),
.B(n_89),
.Y(n_1102)
);

AO21x1_ASAP7_75t_L g1103 ( 
.A1(n_934),
.A2(n_90),
.B(n_91),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_834),
.B(n_92),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_915),
.B(n_92),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_888),
.B(n_94),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_888),
.B(n_94),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_977),
.A2(n_206),
.B(n_292),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_883),
.B(n_96),
.Y(n_1109)
);

CKINVDCx10_ASAP7_75t_R g1110 ( 
.A(n_969),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_868),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_840),
.B(n_98),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_949),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_869),
.B(n_99),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_949),
.B(n_100),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_885),
.B(n_101),
.C(n_102),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_932),
.B(n_929),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_921),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_838),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_946),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_949),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_931),
.B(n_939),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_949),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_891),
.Y(n_1124)
);

AND2x6_ASAP7_75t_L g1125 ( 
.A(n_892),
.B(n_184),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_897),
.B(n_103),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_921),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_966),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_932),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_905),
.B(n_110),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_907),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_910),
.B(n_110),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_894),
.B(n_111),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_848),
.B(n_112),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_848),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_912),
.B(n_114),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_895),
.B(n_884),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_969),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_843),
.B(n_117),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_941),
.A2(n_218),
.B(n_286),
.C(n_285),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_941),
.A2(n_213),
.B(n_284),
.C(n_283),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_845),
.B(n_118),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_934),
.A2(n_209),
.B(n_282),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_972),
.B(n_118),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_835),
.A2(n_208),
.B(n_280),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_935),
.A2(n_214),
.B(n_278),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_861),
.B(n_120),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_943),
.A2(n_959),
.B(n_947),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_935),
.A2(n_223),
.B(n_259),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_960),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_951),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_952),
.B(n_956),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_956),
.B(n_125),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1008),
.B(n_953),
.Y(n_1154)
);

OAI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_986),
.A2(n_969),
.B1(n_858),
.B2(n_862),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1009),
.B(n_898),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1123),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1064),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_1047),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_1001),
.B(n_864),
.Y(n_1160)
);

AND2x6_ASAP7_75t_SL g1161 ( 
.A(n_1010),
.B(n_904),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_993),
.B(n_873),
.Y(n_1162)
);

BUFx12f_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1004),
.A2(n_994),
.B(n_1148),
.Y(n_1164)
);

AOI21xp33_ASAP7_75t_L g1165 ( 
.A1(n_982),
.A2(n_876),
.B(n_886),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_983),
.A2(n_867),
.B(n_936),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1004),
.A2(n_1020),
.B(n_999),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1151),
.B(n_128),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1002),
.A2(n_976),
.A3(n_975),
.B(n_968),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1027),
.B(n_971),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1028),
.B(n_129),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1123),
.Y(n_1172)
);

AO221x2_ASAP7_75t_L g1173 ( 
.A1(n_1076),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.C(n_134),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1098),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1012),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1082),
.B(n_130),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1016),
.B(n_132),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1119),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1117),
.B(n_134),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1012),
.B(n_136),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1062),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_991),
.B(n_136),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_SL g1183 ( 
.A(n_991),
.B(n_1003),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1031),
.A2(n_137),
.B(n_138),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1124),
.B(n_138),
.Y(n_1185)
);

OAI22x1_ASAP7_75t_L g1186 ( 
.A1(n_1025),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_990),
.B(n_1150),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1031),
.A2(n_140),
.B(n_143),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1048),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1108),
.A2(n_188),
.B(n_190),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_SL g1191 ( 
.A1(n_1143),
.A2(n_192),
.B(n_193),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_1066),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1076),
.A2(n_198),
.B(n_200),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1074),
.B(n_237),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_SL g1195 ( 
.A(n_1112),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1120),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_987),
.B(n_1068),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1014),
.A2(n_238),
.B1(n_241),
.B2(n_246),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1113),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1125),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1006),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1078),
.B(n_1052),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1058),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1120),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_987),
.B(n_257),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1110),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1060),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_1095),
.B(n_1115),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1083),
.B(n_1128),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1034),
.A2(n_1141),
.B(n_1140),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1068),
.B(n_1134),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1056),
.A2(n_1057),
.B(n_1036),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1029),
.A2(n_1122),
.B(n_1021),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1137),
.B(n_1131),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1019),
.B(n_1112),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1137),
.B(n_1017),
.Y(n_1216)
);

INVx3_ASAP7_75t_L g1217 ( 
.A(n_1113),
.Y(n_1217)
);

AOI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1063),
.A2(n_1018),
.B(n_1015),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1079),
.B(n_1097),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_984),
.A2(n_1071),
.B(n_1067),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1061),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1099),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_980),
.A2(n_1103),
.A3(n_1077),
.B(n_1153),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1138),
.B(n_988),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1104),
.A2(n_1147),
.B1(n_1144),
.B2(n_1139),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1089),
.A2(n_1046),
.B(n_1145),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1116),
.B(n_1142),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1065),
.A2(n_1146),
.B(n_1149),
.Y(n_1228)
);

BUFx4_ASAP7_75t_SL g1229 ( 
.A(n_1059),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1022),
.B(n_1023),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1026),
.B(n_1035),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1121),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1069),
.A2(n_1070),
.B(n_1093),
.C(n_1096),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1040),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1032),
.B(n_1033),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1075),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1121),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1126),
.A2(n_1136),
.B1(n_1132),
.B2(n_1130),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1037),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_995),
.B(n_1055),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_985),
.B(n_1043),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1049),
.A2(n_1053),
.B(n_1054),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1039),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1037),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1084),
.A2(n_1092),
.B(n_1085),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1087),
.B(n_1088),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1086),
.A2(n_1091),
.B(n_1107),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1101),
.B(n_1105),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1106),
.B(n_1090),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_SL g1251 ( 
.A1(n_1118),
.A2(n_1129),
.B(n_1135),
.Y(n_1251)
);

AOI21x1_ASAP7_75t_SL g1252 ( 
.A1(n_981),
.A2(n_997),
.B(n_1065),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1005),
.A2(n_1013),
.B(n_1109),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1118),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1081),
.B(n_1007),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1114),
.B(n_1100),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1111),
.B(n_998),
.C(n_1102),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1133),
.A2(n_1073),
.B(n_1038),
.C(n_1041),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1044),
.B(n_1072),
.Y(n_1259)
);

AND3x2_ASAP7_75t_L g1260 ( 
.A(n_1073),
.B(n_1125),
.C(n_1127),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1044),
.Y(n_1261)
);

AOI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1000),
.A2(n_1024),
.B(n_1045),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_R g1263 ( 
.A(n_1125),
.B(n_1039),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1123),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_993),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1064),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1064),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1047),
.B(n_881),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1064),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1012),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1008),
.B(n_818),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1064),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1001),
.B(n_810),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1081),
.B(n_743),
.C(n_727),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_979),
.A2(n_983),
.B(n_978),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_979),
.A2(n_983),
.B(n_978),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_993),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_SL g1282 ( 
.A(n_993),
.B(n_806),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1001),
.B(n_810),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_979),
.A2(n_983),
.B(n_978),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_992),
.A2(n_1008),
.B1(n_1009),
.B2(n_818),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_993),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1002),
.A2(n_965),
.A3(n_1011),
.B(n_1042),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1064),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1047),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1064),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_992),
.A2(n_1008),
.B1(n_1009),
.B2(n_818),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1082),
.B(n_828),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1008),
.B(n_818),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_987),
.B(n_806),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1304)
);

OAI21xp33_ASAP7_75t_L g1305 ( 
.A1(n_1152),
.A2(n_828),
.B(n_671),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1080),
.A2(n_881),
.B1(n_846),
.B2(n_809),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1008),
.B(n_818),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_993),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1008),
.B(n_818),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_993),
.B(n_881),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_993),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1001),
.B(n_810),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_993),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1008),
.B(n_818),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1064),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1064),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1008),
.B(n_818),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1001),
.B(n_810),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1094),
.A2(n_954),
.B1(n_890),
.B2(n_980),
.C(n_965),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_SL g1322 ( 
.A(n_1081),
.B(n_743),
.C(n_727),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_996),
.A2(n_965),
.B(n_962),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_993),
.B(n_1012),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1047),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1064),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1064),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1082),
.B(n_828),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1047),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1008),
.B(n_818),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1331)
);

INVx5_ASAP7_75t_L g1332 ( 
.A(n_1012),
.Y(n_1332)
);

AND2x2_ASAP7_75t_SL g1333 ( 
.A(n_1012),
.B(n_846),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_993),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_987),
.B(n_806),
.Y(n_1335)
);

BUFx2_ASAP7_75t_L g1336 ( 
.A(n_1047),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_992),
.A2(n_1008),
.B1(n_1009),
.B2(n_818),
.Y(n_1337)
);

BUFx2_ASAP7_75t_SL g1338 ( 
.A(n_993),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1082),
.B(n_828),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1030),
.A2(n_1150),
.B(n_989),
.C(n_1104),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1001),
.B(n_810),
.Y(n_1342)
);

INVx3_ASAP7_75t_SL g1343 ( 
.A(n_1048),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1064),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1300),
.B(n_1331),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1200),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1163),
.B(n_1281),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1269),
.A2(n_1296),
.B(n_1283),
.Y(n_1349)
);

NOR2x1_ASAP7_75t_SL g1350 ( 
.A(n_1208),
.B(n_1200),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1300),
.B(n_1331),
.Y(n_1351)
);

O2A1O1Ixp33_ASAP7_75t_L g1352 ( 
.A1(n_1306),
.A2(n_1341),
.B(n_1340),
.C(n_1155),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1265),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1157),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1344),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1344),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1206),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1290),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1274),
.B(n_1302),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_SL g1360 ( 
.A1(n_1288),
.A2(n_1337),
.B(n_1299),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1209),
.B(n_1276),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1181),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1334),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1294),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1193),
.A2(n_1251),
.B(n_1233),
.C(n_1218),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1309),
.B(n_1311),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_SL g1367 ( 
.A(n_1200),
.B(n_1338),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1167),
.A2(n_1252),
.B(n_1226),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1172),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1272),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1324),
.Y(n_1371)
);

INVx4_ASAP7_75t_L g1372 ( 
.A(n_1200),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1182),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_SL g1374 ( 
.A(n_1281),
.B(n_1196),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1295),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1284),
.B(n_1314),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1320),
.B(n_1342),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1336),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1210),
.A2(n_1228),
.B(n_1266),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_1316),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1317),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1228),
.A2(n_1277),
.B(n_1273),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1319),
.B(n_1330),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1211),
.B(n_1305),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1318),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1258),
.A2(n_1250),
.B(n_1156),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1183),
.B(n_1208),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1326),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1273),
.A2(n_1286),
.B(n_1277),
.Y(n_1390)
);

NOR2x1_ASAP7_75t_SL g1391 ( 
.A(n_1208),
.B(n_1288),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1182),
.Y(n_1392)
);

CKINVDCx11_ASAP7_75t_R g1393 ( 
.A(n_1343),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1327),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1270),
.B(n_1159),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1308),
.B(n_1171),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1190),
.A2(n_1164),
.B(n_1220),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1168),
.B(n_1325),
.Y(n_1398)
);

INVx6_ASAP7_75t_SL g1399 ( 
.A(n_1312),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1329),
.B(n_1189),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1158),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1264),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1264),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1174),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1243),
.A2(n_1212),
.B(n_1213),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1282),
.B(n_1178),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1310),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1287),
.A2(n_1291),
.B(n_1289),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1173),
.A2(n_1254),
.B1(n_1278),
.B2(n_1322),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1291),
.A2(n_1298),
.B(n_1297),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1227),
.B(n_1215),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1267),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1301),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1297),
.A2(n_1304),
.B(n_1298),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1204),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1192),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1304),
.A2(n_1323),
.B(n_1307),
.Y(n_1417)
);

OR2x6_ASAP7_75t_L g1418 ( 
.A(n_1180),
.B(n_1312),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1328),
.B(n_1339),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1187),
.B(n_1236),
.Y(n_1420)
);

AOI22x1_ASAP7_75t_L g1421 ( 
.A1(n_1191),
.A2(n_1255),
.B1(n_1166),
.B2(n_1205),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1312),
.Y(n_1422)
);

NAND2x1p5_ASAP7_75t_L g1423 ( 
.A(n_1272),
.B(n_1332),
.Y(n_1423)
);

BUFx4_ASAP7_75t_SL g1424 ( 
.A(n_1161),
.Y(n_1424)
);

NOR2xp67_ASAP7_75t_SL g1425 ( 
.A(n_1197),
.B(n_1193),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1268),
.B(n_1271),
.Y(n_1426)
);

NOR2xp67_ASAP7_75t_L g1427 ( 
.A(n_1272),
.B(n_1332),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1247),
.A2(n_1249),
.B(n_1239),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1275),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1246),
.A2(n_1248),
.B(n_1257),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1244),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1246),
.A2(n_1248),
.B(n_1257),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1293),
.Y(n_1433)
);

AO21x1_ASAP7_75t_L g1434 ( 
.A1(n_1184),
.A2(n_1188),
.B(n_1251),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1333),
.B(n_1176),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1313),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1272),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1315),
.Y(n_1438)
);

INVx6_ASAP7_75t_L g1439 ( 
.A(n_1332),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1332),
.B(n_1244),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1253),
.A2(n_1188),
.B(n_1239),
.Y(n_1441)
);

AOI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1205),
.A2(n_1253),
.B1(n_1219),
.B2(n_1242),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1345),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1195),
.Y(n_1444)
);

CKINVDCx14_ASAP7_75t_R g1445 ( 
.A(n_1237),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1185),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1180),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1202),
.B(n_1201),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1177),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1225),
.B(n_1321),
.C(n_1173),
.Y(n_1450)
);

BUFx4f_ASAP7_75t_L g1451 ( 
.A(n_1162),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1162),
.Y(n_1452)
);

CKINVDCx16_ASAP7_75t_R g1453 ( 
.A(n_1195),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1160),
.B(n_1203),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1154),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1232),
.A2(n_1238),
.B(n_1259),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1179),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1214),
.B(n_1234),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1186),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1229),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1165),
.A2(n_1230),
.B(n_1231),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1241),
.A2(n_1263),
.B(n_1235),
.Y(n_1462)
);

AOI22x1_ASAP7_75t_L g1463 ( 
.A1(n_1207),
.A2(n_1222),
.B1(n_1221),
.B2(n_1256),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1175),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1169),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1175),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1169),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1170),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1216),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1194),
.A2(n_1260),
.B1(n_1198),
.B2(n_1224),
.Y(n_1470)
);

BUFx10_ASAP7_75t_L g1471 ( 
.A(n_1245),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1232),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1262),
.A2(n_1261),
.B(n_1199),
.Y(n_1473)
);

INVx5_ASAP7_75t_SL g1474 ( 
.A(n_1238),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1240),
.A2(n_1217),
.B1(n_1262),
.B2(n_1303),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1335),
.A2(n_1240),
.B(n_1223),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1223),
.B(n_1292),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1292),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1294),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1279),
.A2(n_1285),
.B(n_1280),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1274),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1344),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1274),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1300),
.B(n_1331),
.Y(n_1484)
);

BUFx4f_ASAP7_75t_SL g1485 ( 
.A(n_1163),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1485),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1362),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1485),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1388),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1388),
.B(n_1350),
.Y(n_1490)
);

BUFx10_ASAP7_75t_L g1491 ( 
.A(n_1388),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1401),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1405),
.A2(n_1368),
.B(n_1397),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1380),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1420),
.B(n_1355),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1480),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1425),
.B(n_1367),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1404),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1396),
.A2(n_1434),
.B1(n_1377),
.B2(n_1399),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1418),
.B(n_1423),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1420),
.A2(n_1361),
.B1(n_1366),
.B2(n_1359),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1412),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1429),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1433),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1481),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1423),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1443),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1428),
.A2(n_1365),
.B(n_1387),
.Y(n_1508)
);

CKINVDCx16_ASAP7_75t_R g1509 ( 
.A(n_1357),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1426),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1356),
.B(n_1482),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1376),
.B(n_1377),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1393),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1393),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1483),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1375),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1381),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1389),
.Y(n_1518)
);

OAI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1418),
.A2(n_1392),
.B1(n_1483),
.B2(n_1399),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1353),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1452),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1454),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1371),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1371),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1452),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1386),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_SL g1527 ( 
.A1(n_1391),
.A2(n_1360),
.B(n_1456),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1418),
.B(n_1427),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1447),
.A2(n_1422),
.B1(n_1373),
.B2(n_1442),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_SL g1530 ( 
.A1(n_1373),
.A2(n_1459),
.B1(n_1463),
.B2(n_1416),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1399),
.A2(n_1450),
.B1(n_1411),
.B2(n_1361),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1394),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1373),
.A2(n_1351),
.B1(n_1406),
.B2(n_1441),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1448),
.Y(n_1534)
);

NAND2x1_ASAP7_75t_L g1535 ( 
.A(n_1347),
.B(n_1372),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1383),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1351),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1359),
.A2(n_1366),
.B1(n_1411),
.B2(n_1435),
.Y(n_1538)
);

NAND2x1_ASAP7_75t_L g1539 ( 
.A(n_1347),
.B(n_1372),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1351),
.B(n_1419),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1346),
.B(n_1484),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1472),
.B(n_1369),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1455),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1458),
.B(n_1398),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1406),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1406),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1413),
.B(n_1468),
.Y(n_1547)
);

AO21x1_ASAP7_75t_SL g1548 ( 
.A1(n_1470),
.A2(n_1409),
.B(n_1475),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1354),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1366),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1383),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1395),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1384),
.A2(n_1446),
.B1(n_1453),
.B2(n_1349),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1353),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1364),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1441),
.A2(n_1378),
.B1(n_1474),
.B2(n_1451),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1451),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1385),
.B(n_1479),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1407),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1464),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1444),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1466),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1474),
.A2(n_1472),
.B1(n_1462),
.B2(n_1374),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1515),
.B(n_1365),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1496),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_SL g1566 ( 
.A1(n_1556),
.A2(n_1470),
.B(n_1409),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1491),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1494),
.B(n_1477),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1501),
.A2(n_1352),
.B1(n_1432),
.B2(n_1430),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1570)
);

BUFx4f_ASAP7_75t_SL g1571 ( 
.A(n_1513),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1526),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1494),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1512),
.B(n_1478),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1505),
.A2(n_1475),
.B1(n_1449),
.B2(n_1474),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1550),
.B(n_1414),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1505),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1548),
.Y(n_1579)
);

INVx5_ASAP7_75t_SL g1580 ( 
.A(n_1500),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1538),
.A2(n_1457),
.B1(n_1372),
.B2(n_1347),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1499),
.B(n_1414),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1520),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1499),
.B(n_1543),
.Y(n_1584)
);

NOR2xp67_ASAP7_75t_L g1585 ( 
.A(n_1490),
.B(n_1369),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1520),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1491),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1390),
.Y(n_1588)
);

NAND2x1_ASAP7_75t_L g1589 ( 
.A(n_1527),
.B(n_1402),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1492),
.B(n_1390),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1531),
.A2(n_1469),
.B1(n_1461),
.B2(n_1476),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1490),
.B(n_1465),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1498),
.B(n_1390),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1502),
.B(n_1408),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1503),
.B(n_1408),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1490),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1504),
.B(n_1408),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1511),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1507),
.B(n_1410),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1544),
.B(n_1487),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1542),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1542),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1537),
.A2(n_1489),
.B1(n_1500),
.B2(n_1528),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1531),
.A2(n_1558),
.B1(n_1519),
.B2(n_1540),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1516),
.B(n_1417),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1566),
.A2(n_1495),
.B1(n_1500),
.B2(n_1534),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1565),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1572),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1555),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1570),
.B(n_1467),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1580),
.A2(n_1537),
.B1(n_1528),
.B2(n_1506),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_1382),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1588),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1382),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1379),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1591),
.B(n_1417),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1578),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1606),
.A2(n_1519),
.B1(n_1497),
.B2(n_1533),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1601),
.B(n_1522),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1594),
.B(n_1417),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1510),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1578),
.Y(n_1625)
);

BUFx12f_ASAP7_75t_L g1626 ( 
.A(n_1567),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1493),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1598),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1574),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1493),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1603),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1576),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1571),
.B(n_1509),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1600),
.Y(n_1635)
);

NOR3xp33_ASAP7_75t_L g1636 ( 
.A(n_1566),
.B(n_1547),
.C(n_1559),
.Y(n_1636)
);

AND2x4_ASAP7_75t_SL g1637 ( 
.A(n_1593),
.B(n_1528),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1584),
.A2(n_1497),
.B1(n_1461),
.B2(n_1537),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1605),
.A2(n_1563),
.B1(n_1530),
.B2(n_1506),
.Y(n_1639)
);

AND2x4_ASAP7_75t_SL g1640 ( 
.A(n_1567),
.B(n_1587),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1610),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1610),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1615),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1628),
.B(n_1582),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1609),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1615),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1632),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1627),
.B(n_1600),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1627),
.B(n_1577),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1611),
.B(n_1599),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1654)
);

AOI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1636),
.A2(n_1569),
.B1(n_1599),
.B2(n_1575),
.C(n_1579),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1633),
.B(n_1607),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1634),
.B(n_1513),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1625),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1577),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.B(n_1607),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1608),
.A2(n_1579),
.B(n_1604),
.C(n_1603),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1646),
.B(n_1619),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1642),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1642),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1647),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1643),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1646),
.B(n_1620),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1629),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1648),
.B(n_1614),
.Y(n_1670)
);

OR2x2_ASAP7_75t_SL g1671 ( 
.A(n_1658),
.B(n_1586),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1625),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1641),
.B(n_1618),
.Y(n_1673)
);

NAND4xp75_ASAP7_75t_L g1674 ( 
.A(n_1655),
.B(n_1608),
.C(n_1585),
.D(n_1587),
.Y(n_1674)
);

NOR5xp2_ASAP7_75t_L g1675 ( 
.A(n_1662),
.B(n_1602),
.C(n_1590),
.D(n_1424),
.E(n_1549),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1644),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1644),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1649),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1649),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1651),
.B(n_1623),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1656),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1612),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1664),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1664),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1665),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1665),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1682),
.B(n_1660),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1686),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1671),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1675),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1685),
.A2(n_1639),
.B1(n_1621),
.B2(n_1654),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1682),
.B(n_1684),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1684),
.B(n_1660),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1666),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1645),
.Y(n_1700)
);

AOI32xp33_ASAP7_75t_L g1701 ( 
.A1(n_1671),
.A2(n_1605),
.A3(n_1613),
.B1(n_1637),
.B2(n_1640),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1674),
.A2(n_1597),
.B1(n_1580),
.B2(n_1622),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1663),
.B(n_1672),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1669),
.B(n_1652),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1683),
.B(n_1657),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1670),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1676),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1670),
.B(n_1652),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1668),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1707),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1701),
.A2(n_1460),
.B(n_1486),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1688),
.Y(n_1713)
);

OAI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1694),
.A2(n_1631),
.B1(n_1597),
.B2(n_1626),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1688),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1701),
.B(n_1638),
.C(n_1686),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1689),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1695),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1690),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1710),
.Y(n_1721)
);

OAI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1696),
.A2(n_1687),
.B(n_1661),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1702),
.A2(n_1525),
.B(n_1521),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1690),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1692),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1721),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1712),
.A2(n_1698),
.B1(n_1697),
.B2(n_1692),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1711),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1718),
.A2(n_1514),
.B(n_1488),
.C(n_1706),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1718),
.A2(n_1708),
.B1(n_1703),
.B2(n_1691),
.C(n_1693),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1723),
.B(n_1514),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1715),
.B(n_1698),
.Y(n_1733)
);

OAI332xp33_ASAP7_75t_L g1734 ( 
.A1(n_1714),
.A2(n_1700),
.A3(n_1705),
.B1(n_1569),
.B2(n_1445),
.B3(n_1654),
.C1(n_1661),
.C2(n_1575),
.Y(n_1734)
);

XNOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1714),
.B(n_1460),
.Y(n_1735)
);

NOR3xp33_ASAP7_75t_L g1736 ( 
.A(n_1716),
.B(n_1674),
.C(n_1348),
.Y(n_1736)
);

OAI322xp33_ASAP7_75t_L g1737 ( 
.A1(n_1717),
.A2(n_1693),
.A3(n_1691),
.B1(n_1673),
.B2(n_1704),
.C1(n_1699),
.C2(n_1709),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1724),
.A2(n_1698),
.B(n_1708),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1719),
.A2(n_1445),
.B(n_1698),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1720),
.B(n_1709),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1736),
.B(n_1415),
.C(n_1436),
.Y(n_1741)
);

NOR4xp25_ASAP7_75t_SL g1742 ( 
.A(n_1730),
.B(n_1486),
.C(n_1415),
.D(n_1545),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1732),
.A2(n_1708),
.B(n_1640),
.C(n_1604),
.Y(n_1743)
);

OAI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1725),
.A2(n_1704),
.B(n_1699),
.Y(n_1744)
);

NOR4xp25_ASAP7_75t_SL g1745 ( 
.A(n_1728),
.B(n_1546),
.C(n_1678),
.D(n_1681),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1726),
.B(n_1357),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1733),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1739),
.B(n_1659),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1735),
.Y(n_1749)
);

O2A1O1Ixp5_ASAP7_75t_L g1750 ( 
.A1(n_1739),
.A2(n_1704),
.B(n_1699),
.C(n_1589),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1727),
.A2(n_1581),
.B1(n_1680),
.B2(n_1679),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1729),
.A2(n_1400),
.B(n_1561),
.C(n_1363),
.Y(n_1752)
);

OAI221xp5_ASAP7_75t_R g1753 ( 
.A1(n_1734),
.A2(n_1592),
.B1(n_1529),
.B2(n_1580),
.C(n_1444),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1747),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1751),
.B(n_1740),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1746),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_L g1759 ( 
.A(n_1741),
.B(n_1737),
.C(n_1358),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1667),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1750),
.Y(n_1761)
);

NAND5xp2_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1557),
.C(n_1444),
.D(n_1440),
.E(n_1541),
.Y(n_1762)
);

OA22x2_ASAP7_75t_SL g1763 ( 
.A1(n_1753),
.A2(n_1581),
.B1(n_1580),
.B2(n_1626),
.Y(n_1763)
);

AOI31xp33_ASAP7_75t_L g1764 ( 
.A1(n_1752),
.A2(n_1438),
.A3(n_1551),
.B(n_1536),
.Y(n_1764)
);

NOR2xp67_ASAP7_75t_L g1765 ( 
.A(n_1744),
.B(n_1677),
.Y(n_1765)
);

NOR4xp75_ASAP7_75t_L g1766 ( 
.A(n_1755),
.B(n_1758),
.C(n_1756),
.D(n_1763),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1754),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1757),
.Y(n_1768)
);

NAND4xp75_ASAP7_75t_L g1769 ( 
.A(n_1761),
.B(n_1742),
.C(n_1743),
.D(n_1585),
.Y(n_1769)
);

NOR3xp33_ASAP7_75t_L g1770 ( 
.A(n_1764),
.B(n_1370),
.C(n_1437),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_L g1771 ( 
.A(n_1762),
.B(n_1370),
.C(n_1523),
.Y(n_1771)
);

NOR3x2_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1439),
.C(n_1471),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1760),
.B(n_1759),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1765),
.B(n_1369),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1757),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1757),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1757),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1757),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1767),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1768),
.Y(n_1780)
);

BUFx12f_ASAP7_75t_L g1781 ( 
.A(n_1766),
.Y(n_1781)
);

NOR2xp67_ASAP7_75t_L g1782 ( 
.A(n_1775),
.B(n_1567),
.Y(n_1782)
);

NOR4xp75_ASAP7_75t_L g1783 ( 
.A(n_1769),
.B(n_1524),
.C(n_1539),
.D(n_1535),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1776),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1779),
.B(n_1777),
.Y(n_1785)
);

NAND4xp75_ASAP7_75t_L g1786 ( 
.A(n_1780),
.B(n_1778),
.C(n_1773),
.D(n_1774),
.Y(n_1786)
);

XNOR2xp5_ASAP7_75t_L g1787 ( 
.A(n_1783),
.B(n_1772),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1784),
.Y(n_1788)
);

NAND4xp75_ASAP7_75t_L g1789 ( 
.A(n_1781),
.B(n_1782),
.C(n_1770),
.D(n_1771),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1785),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1787),
.A2(n_1781),
.B1(n_1771),
.B2(n_1580),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1791),
.A2(n_1790),
.B(n_1788),
.Y(n_1792)
);

OA21x2_ASAP7_75t_L g1793 ( 
.A1(n_1790),
.A2(n_1789),
.B(n_1786),
.Y(n_1793)
);

AOI21xp33_ASAP7_75t_SL g1794 ( 
.A1(n_1793),
.A2(n_1440),
.B(n_1587),
.Y(n_1794)
);

AO22x2_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1437),
.B1(n_1517),
.B2(n_1518),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1795),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1794),
.A2(n_1562),
.B(n_1560),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1797),
.B1(n_1431),
.B2(n_1604),
.C(n_1603),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1589),
.B(n_1431),
.Y(n_1799)
);

OA21x2_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1421),
.B(n_1473),
.Y(n_1800)
);

AOI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1431),
.B(n_1403),
.Y(n_1801)
);


endmodule