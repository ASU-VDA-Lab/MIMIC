module fake_netlist_5_1876_n_816 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_816);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_816;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_718;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_813;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_793;
wire n_478;
wire n_726;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_795;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_401;
wire n_187;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_23),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_4),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_49),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_107),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_7),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_59),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_4),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_17),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_119),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_53),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_0),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_77),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_99),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_66),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_83),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_58),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_85),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_75),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_61),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_93),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_26),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_131),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_39),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_72),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_37),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_45),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_95),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_103),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_63),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_9),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_35),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_15),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_51),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_92),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_24),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_147),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_113),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_171),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_173),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_165),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_175),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_0),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_R g245 ( 
.A(n_168),
.B(n_1),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_178),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_189),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_R g249 ( 
.A(n_166),
.B(n_197),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_176),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_217),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_197),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_222),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_204),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_168),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_179),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_191),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_191),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_238),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_216),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_230),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_211),
.B(n_212),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_180),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_203),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_249),
.B(n_212),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_224),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_248),
.B(n_182),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_247),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_187),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_227),
.B(n_213),
.Y(n_306)
);

INVx6_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_263),
.A2(n_213),
.B1(n_221),
.B2(n_220),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_265),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_237),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_190),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_274),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_192),
.Y(n_322)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_259),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_250),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_250),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

AND2x6_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_25),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_193),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_194),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_198),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_199),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_272),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_282),
.B(n_295),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_271),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_271),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_27),
.Y(n_346)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_282),
.B(n_202),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_296),
.B(n_208),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_293),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_254),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_279),
.B(n_209),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_272),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_254),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_316),
.B(n_210),
.Y(n_360)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_282),
.Y(n_361)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_28),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_277),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_215),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_273),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_308),
.A2(n_219),
.B1(n_223),
.B2(n_5),
.Y(n_368)
);

AND2x6_ASAP7_75t_SL g369 ( 
.A(n_298),
.B(n_2),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_279),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_282),
.B(n_30),
.Y(n_371)
);

AND2x4_ASAP7_75t_SL g372 ( 
.A(n_316),
.B(n_31),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_293),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_273),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_2),
.B(n_3),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_3),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_283),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_287),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_286),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_286),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_295),
.Y(n_384)
);

BUFx4f_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_297),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_325),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_351),
.A2(n_309),
.B1(n_304),
.B2(n_297),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_385),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_350),
.B(n_297),
.Y(n_392)
);

AO22x2_ASAP7_75t_L g393 ( 
.A1(n_368),
.A2(n_313),
.B1(n_310),
.B2(n_311),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_353),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_349),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_297),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

INVx3_ASAP7_75t_R g400 ( 
.A(n_333),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

NAND3xp33_ASAP7_75t_SL g403 ( 
.A(n_376),
.B(n_311),
.C(n_310),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

AO22x2_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_315),
.B1(n_304),
.B2(n_302),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_373),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

OAI221xp5_ASAP7_75t_L g412 ( 
.A1(n_381),
.A2(n_285),
.B1(n_284),
.B2(n_308),
.C(n_295),
.Y(n_412)
);

AO22x2_ASAP7_75t_L g413 ( 
.A1(n_357),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_319),
.B(n_280),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_285),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_335),
.B(n_346),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_293),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_319),
.B(n_305),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_374),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_385),
.Y(n_427)
);

XNOR2x2_ASAP7_75t_SL g428 ( 
.A(n_369),
.B(n_318),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_375),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_369),
.A2(n_315),
.B1(n_317),
.B2(n_275),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_381),
.A2(n_287),
.B1(n_377),
.B2(n_382),
.Y(n_431)
);

AO22x2_ASAP7_75t_L g432 ( 
.A1(n_322),
.A2(n_317),
.B1(n_293),
.B2(n_9),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_383),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_317),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_322),
.B(n_288),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_347),
.B(n_314),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_269),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_329),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_342),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_321),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g443 ( 
.A1(n_337),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g444 ( 
.A1(n_337),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

AND2x2_ASAP7_75t_SL g446 ( 
.A(n_372),
.B(n_287),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_348),
.B(n_287),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_348),
.B(n_276),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_332),
.Y(n_449)
);

OAI221xp5_ASAP7_75t_L g450 ( 
.A1(n_377),
.A2(n_276),
.B1(n_294),
.B2(n_270),
.C(n_269),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g451 ( 
.A1(n_339),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_380),
.Y(n_452)
);

OAI221xp5_ASAP7_75t_L g453 ( 
.A1(n_364),
.A2(n_270),
.B1(n_307),
.B2(n_17),
.C(n_18),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_360),
.A2(n_307),
.B1(n_98),
.B2(n_100),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_341),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_370),
.B(n_307),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_400),
.B(n_356),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_415),
.B(n_355),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_435),
.B(n_339),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_365),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_421),
.B(n_380),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_356),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_424),
.B(n_370),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_390),
.B(n_329),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_427),
.B(n_363),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_387),
.B(n_363),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_401),
.B(n_394),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_392),
.B(n_363),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_399),
.B(n_361),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_395),
.B(n_371),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_397),
.B(n_361),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_409),
.B(n_371),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_386),
.B(n_338),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_419),
.B(n_361),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_389),
.B(n_361),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_434),
.B(n_379),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_SL g478 ( 
.A(n_452),
.B(n_335),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_423),
.B(n_379),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_436),
.B(n_379),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_SL g481 ( 
.A(n_431),
.B(n_335),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_SL g482 ( 
.A(n_418),
.B(n_335),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_386),
.B(n_323),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_416),
.B(n_391),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_455),
.B(n_323),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_416),
.B(n_379),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_396),
.B(n_345),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_402),
.B(n_345),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_420),
.B(n_346),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_404),
.B(n_323),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_406),
.B(n_362),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_410),
.B(n_346),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_414),
.B(n_362),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_417),
.B(n_362),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_422),
.B(n_362),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_346),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_425),
.B(n_33),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_426),
.B(n_34),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_429),
.B(n_14),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_SL g500 ( 
.A(n_448),
.B(n_456),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_457),
.B(n_36),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_16),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_456),
.B(n_16),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_442),
.B(n_38),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_445),
.B(n_40),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_449),
.B(n_43),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_447),
.B(n_18),
.Y(n_507)
);

NAND2xp33_ASAP7_75t_SL g508 ( 
.A(n_388),
.B(n_19),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_454),
.B(n_44),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_19),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_388),
.B(n_47),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_438),
.B(n_48),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_484),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_468),
.B(n_413),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_483),
.A2(n_405),
.B(n_398),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_481),
.A2(n_412),
.B(n_450),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_503),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_496),
.A2(n_403),
.B(n_441),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_398),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_460),
.A2(n_463),
.B1(n_473),
.B2(n_471),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_405),
.B(n_411),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_487),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_413),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_461),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_461),
.B(n_411),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_485),
.A2(n_407),
.B(n_437),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_492),
.B(n_439),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_464),
.A2(n_453),
.B(n_432),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_474),
.B(n_408),
.Y(n_531)
);

AO31x2_ASAP7_75t_L g532 ( 
.A1(n_510),
.A2(n_432),
.A3(n_444),
.B(n_443),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_488),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_467),
.A2(n_469),
.B(n_494),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_470),
.B(n_408),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_493),
.A2(n_393),
.B(n_444),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_500),
.A2(n_393),
.B(n_443),
.C(n_451),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_482),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_489),
.A2(n_472),
.B(n_495),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_509),
.A2(n_451),
.B(n_430),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_490),
.A2(n_476),
.B(n_512),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_507),
.A2(n_430),
.B(n_428),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_466),
.B(n_465),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_501),
.A2(n_109),
.B(n_161),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_479),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_475),
.B(n_20),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_486),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_477),
.A2(n_106),
.B(n_159),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_105),
.B(n_158),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_498),
.A2(n_104),
.B(n_157),
.Y(n_553)
);

NOR2xp67_ASAP7_75t_SL g554 ( 
.A(n_480),
.B(n_20),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_458),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_504),
.B(n_505),
.Y(n_556)
);

OAI22x1_ASAP7_75t_L g557 ( 
.A1(n_462),
.A2(n_506),
.B1(n_22),
.B2(n_23),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_516),
.A2(n_21),
.B1(n_22),
.B2(n_50),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_521),
.A2(n_515),
.B(n_526),
.Y(n_559)
);

A2O1A1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_516),
.A2(n_21),
.B(n_52),
.C(n_54),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_513),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_524),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_517),
.A2(n_55),
.B1(n_57),
.B2(n_60),
.Y(n_565)
);

OAI221xp5_ASAP7_75t_L g566 ( 
.A1(n_542),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.C(n_67),
.Y(n_566)
);

AOI22x1_ASAP7_75t_L g567 ( 
.A1(n_557),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_542),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_568)
);

OR2x6_ASAP7_75t_L g569 ( 
.A(n_530),
.B(n_76),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_540),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_571)
);

AOI21x1_ASAP7_75t_L g572 ( 
.A1(n_539),
.A2(n_529),
.B(n_541),
.Y(n_572)
);

OAI22xp33_ASAP7_75t_L g573 ( 
.A1(n_548),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_535),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

CKINVDCx11_ASAP7_75t_R g576 ( 
.A(n_524),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_531),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_551),
.A2(n_555),
.B1(n_520),
.B2(n_514),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_537),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_518),
.A2(n_89),
.B(n_90),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_91),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_518),
.A2(n_96),
.B(n_97),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_527),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_544),
.A2(n_101),
.B(n_102),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_555),
.B(n_111),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_534),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_549),
.A2(n_114),
.B(n_115),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_545),
.B(n_117),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_554),
.B(n_118),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_525),
.B(n_121),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_550),
.B(n_122),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_519),
.B(n_124),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_536),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_536),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_598),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_590),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_586),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_532),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_559),
.A2(n_553),
.B(n_534),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_572),
.A2(n_523),
.B(n_544),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_578),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_562),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_584),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_599),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_561),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_591),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_564),
.B(n_552),
.Y(n_616)
);

AO21x2_ASAP7_75t_L g617 ( 
.A1(n_579),
.A2(n_538),
.B(n_532),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_581),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_585),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_562),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_558),
.B(n_532),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_576),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_587),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_579),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_596),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_596),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_567),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_558),
.B(n_556),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_583),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_571),
.A2(n_556),
.B1(n_126),
.B2(n_127),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_580),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_583),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_597),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_562),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_569),
.B(n_580),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_569),
.B(n_125),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_560),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_568),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_566),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_588),
.B(n_136),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_560),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_563),
.Y(n_651)
);

AOI21x1_ASAP7_75t_L g652 ( 
.A1(n_565),
.A2(n_138),
.B(n_139),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_593),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_638),
.B(n_593),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_615),
.B(n_568),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_606),
.B(n_595),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_600),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_R g658 ( 
.A(n_642),
.B(n_593),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_R g660 ( 
.A(n_616),
.B(n_571),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_R g661 ( 
.A(n_638),
.B(n_140),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_648),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_622),
.B(n_573),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_642),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_602),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_L g666 ( 
.A(n_640),
.B(n_573),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_650),
.B(n_637),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_650),
.B(n_141),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_606),
.B(n_594),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_R g670 ( 
.A(n_642),
.B(n_653),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_642),
.B(n_142),
.Y(n_671)
);

CKINVDCx11_ASAP7_75t_R g672 ( 
.A(n_640),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_R g673 ( 
.A(n_647),
.B(n_143),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_594),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_R g675 ( 
.A(n_647),
.B(n_653),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_603),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_566),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_646),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_607),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_631),
.B(n_146),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_R g681 ( 
.A(n_641),
.B(n_632),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_603),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_631),
.B(n_148),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_611),
.B(n_149),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_R g685 ( 
.A(n_641),
.B(n_150),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_R g686 ( 
.A(n_647),
.B(n_162),
.Y(n_686)
);

BUFx10_ASAP7_75t_L g687 ( 
.A(n_607),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_651),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_607),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_650),
.B(n_151),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_637),
.B(n_152),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_R g692 ( 
.A(n_641),
.B(n_153),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_607),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_611),
.B(n_156),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_633),
.B(n_154),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_666),
.A2(n_644),
.B1(n_641),
.B2(n_645),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_676),
.B(n_621),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_657),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_656),
.B(n_626),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_667),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_660),
.B(n_636),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_659),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_682),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_667),
.B(n_621),
.Y(n_704)
);

NAND2x1_ASAP7_75t_L g705 ( 
.A(n_669),
.B(n_629),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_663),
.A2(n_632),
.B1(n_634),
.B2(n_643),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_674),
.Y(n_707)
);

NAND2x1_ASAP7_75t_L g708 ( 
.A(n_677),
.B(n_629),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_688),
.B(n_617),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_684),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_675),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_662),
.B(n_626),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_608),
.Y(n_713)
);

BUFx12f_ASAP7_75t_L g714 ( 
.A(n_672),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_693),
.B(n_610),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_654),
.B(n_617),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_664),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_694),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_689),
.B(n_623),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_679),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_664),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_680),
.B(n_617),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_678),
.A2(n_649),
.B1(n_643),
.B2(n_635),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_679),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_683),
.B(n_623),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_695),
.B(n_625),
.Y(n_726)
);

AO21x2_ASAP7_75t_L g727 ( 
.A1(n_710),
.A2(n_624),
.B(n_625),
.Y(n_727)
);

OAI31xp33_ASAP7_75t_L g728 ( 
.A1(n_696),
.A2(n_706),
.A3(n_718),
.B(n_710),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_665),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_716),
.B(n_624),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_723),
.A2(n_649),
.B1(n_635),
.B2(n_630),
.Y(n_731)
);

AOI221xp5_ASAP7_75t_L g732 ( 
.A1(n_718),
.A2(n_613),
.B1(n_630),
.B2(n_608),
.C(n_612),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_704),
.B(n_610),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_707),
.B(n_613),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_698),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_701),
.A2(n_714),
.B1(n_605),
.B2(n_661),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_697),
.B(n_619),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_708),
.A2(n_671),
.B1(n_685),
.B2(n_692),
.C(n_658),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_698),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_702),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_702),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_714),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_703),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_743),
.B(n_707),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_730),
.B(n_716),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_730),
.B(n_697),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_737),
.B(n_722),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_733),
.B(n_713),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_729),
.B(n_739),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_740),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_734),
.B(n_703),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_735),
.B(n_709),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_735),
.B(n_722),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_728),
.A2(n_708),
.B(n_711),
.Y(n_754)
);

NOR2x1_ASAP7_75t_SL g755 ( 
.A(n_727),
.B(n_709),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_R g756 ( 
.A(n_754),
.B(n_673),
.Y(n_756)
);

AO221x2_ASAP7_75t_L g757 ( 
.A1(n_744),
.A2(n_738),
.B1(n_742),
.B2(n_712),
.C(n_724),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_748),
.B(n_739),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_749),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_747),
.B(n_742),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_751),
.B(n_740),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_745),
.B(n_742),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_747),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_760),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_761),
.Y(n_766)
);

XOR2x2_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_756),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_765),
.A2(n_757),
.B1(n_670),
.B2(n_736),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_766),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_764),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_770),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_769),
.B(n_758),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_767),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_771),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_773),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_771),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_775),
.A2(n_768),
.B(n_736),
.Y(n_778)
);

NAND4xp25_ASAP7_75t_SL g779 ( 
.A(n_776),
.B(n_731),
.C(n_759),
.D(n_732),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_777),
.B(n_720),
.C(n_668),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_774),
.A2(n_731),
.B1(n_752),
.B2(n_750),
.Y(n_781)
);

NOR2x1_ASAP7_75t_L g782 ( 
.A(n_774),
.B(n_690),
.Y(n_782)
);

AOI221xp5_ASAP7_75t_L g783 ( 
.A1(n_779),
.A2(n_686),
.B1(n_715),
.B2(n_699),
.C(n_720),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_SL g784 ( 
.A(n_778),
.B(n_705),
.C(n_636),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_782),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_780),
.A2(n_715),
.B1(n_681),
.B2(n_721),
.Y(n_786)
);

AOI221xp5_ASAP7_75t_L g787 ( 
.A1(n_781),
.A2(n_715),
.B1(n_753),
.B2(n_705),
.C(n_668),
.Y(n_787)
);

AOI221xp5_ASAP7_75t_L g788 ( 
.A1(n_779),
.A2(n_753),
.B1(n_690),
.B2(n_746),
.C(n_721),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_778),
.B(n_695),
.C(n_691),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_788),
.A2(n_717),
.B1(n_727),
.B2(n_741),
.Y(n_790)
);

NOR2x1_ASAP7_75t_SL g791 ( 
.A(n_785),
.B(n_607),
.Y(n_791)
);

NOR2x1_ASAP7_75t_L g792 ( 
.A(n_784),
.B(n_691),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_783),
.B(n_746),
.Y(n_793)
);

NAND4xp75_ASAP7_75t_L g794 ( 
.A(n_787),
.B(n_620),
.C(n_639),
.D(n_755),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_786),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_R g796 ( 
.A(n_795),
.B(n_155),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_793),
.B(n_791),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_R g798 ( 
.A(n_792),
.B(n_789),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_R g799 ( 
.A(n_794),
.B(n_652),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_796),
.B(n_620),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_797),
.Y(n_801)
);

NAND2x1_ASAP7_75t_L g802 ( 
.A(n_798),
.B(n_790),
.Y(n_802)
);

OAI21xp33_ASAP7_75t_L g803 ( 
.A1(n_799),
.A2(n_717),
.B(n_741),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_801),
.A2(n_717),
.B1(n_633),
.B2(n_719),
.Y(n_804)
);

INVxp67_ASAP7_75t_SL g805 ( 
.A(n_802),
.Y(n_805)
);

OR5x1_ASAP7_75t_L g806 ( 
.A(n_803),
.B(n_687),
.C(n_652),
.D(n_639),
.E(n_651),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_800),
.B(n_700),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_805),
.B(n_612),
.C(n_614),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_807),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_809),
.A2(n_804),
.B1(n_806),
.B2(n_628),
.Y(n_810)
);

AOI31xp33_ASAP7_75t_L g811 ( 
.A1(n_808),
.A2(n_628),
.A3(n_614),
.B(n_726),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_SL g812 ( 
.A(n_810),
.B(n_719),
.C(n_618),
.Y(n_812)
);

AOI222xp33_ASAP7_75t_L g813 ( 
.A1(n_812),
.A2(n_811),
.B1(n_619),
.B2(n_618),
.C1(n_627),
.C2(n_726),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_813),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_814),
.A2(n_627),
.B1(n_700),
.B2(n_725),
.C(n_601),
.Y(n_815)
);

AOI211xp5_ASAP7_75t_L g816 ( 
.A1(n_815),
.A2(n_725),
.B(n_700),
.C(n_604),
.Y(n_816)
);


endmodule