module fake_jpeg_25667_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_21),
.C(n_20),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_20),
.C(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_25),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_56),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_19),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_19),
.B(n_13),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_62),
.C(n_18),
.Y(n_81)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_61),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_64),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_10),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_13),
.B(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_24),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_80),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_83),
.Y(n_92)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_18),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_53),
.B(n_51),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_71),
.B(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_91),
.B1(n_72),
.B2(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_96),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_66),
.B1(n_61),
.B2(n_57),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_59),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.C(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_71),
.B1(n_72),
.B2(n_83),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_79),
.B1(n_17),
.B2(n_12),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_17),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_75),
.B1(n_50),
.B2(n_79),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_17),
.B(n_12),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_67),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_84),
.B(n_86),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_109),
.C(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_97),
.B1(n_95),
.B2(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_112),
.B(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_100),
.C(n_98),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_104),
.C(n_116),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_106),
.C(n_7),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_119),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_128),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_113),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_114),
.B1(n_118),
.B2(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_127),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_104),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_110),
.C(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_5),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_6),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_8),
.C(n_10),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_137),
.A2(n_134),
.B(n_8),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_138),
.Y(n_140)
);


endmodule