module fake_netlist_5_2536_n_1738 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1738);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1738;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_69),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_51),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_46),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_87),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

BUFx8_ASAP7_75t_SL g182 ( 
.A(n_152),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_67),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_12),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_29),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_53),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_100),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_41),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_38),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_123),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_14),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_32),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_21),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_75),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_17),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_108),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_44),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_43),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_97),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_71),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_85),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_159),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_51),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_144),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_56),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_13),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_117),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_25),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_72),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_47),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_127),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_98),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_50),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_4),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g242 ( 
.A(n_39),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_47),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_50),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_148),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_86),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_151),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_37),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_101),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_16),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_90),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_48),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_62),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_170),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_52),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_128),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_166),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_135),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_84),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_37),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_82),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_102),
.Y(n_268)
);

CKINVDCx11_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_1),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_27),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_119),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_83),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_150),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_171),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_79),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_21),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_34),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_55),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_48),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_22),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_136),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_88),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_130),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_163),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_18),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_160),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_99),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_11),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_3),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_113),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_115),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_161),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_26),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_20),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_120),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_114),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_61),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_65),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_57),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_140),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_27),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_165),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_1),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_121),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_174),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_110),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_19),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_57),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_169),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_41),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_167),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_23),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_125),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_14),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_96),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_104),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_20),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_58),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_173),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_24),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_168),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_147),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_155),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_129),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_70),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_122),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_134),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_22),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_33),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_126),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_153),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_77),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_52),
.Y(n_346)
);

BUFx2_ASAP7_75t_SL g347 ( 
.A(n_226),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_186),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_242),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_182),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_269),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_204),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_242),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_242),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_302),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_242),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_181),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_242),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_242),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_242),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_252),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_209),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_267),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_181),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_277),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_228),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_177),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_211),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_206),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_206),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_235),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_264),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_212),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_185),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_216),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_213),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_304),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_213),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_293),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_311),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_217),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_293),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_235),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g394 ( 
.A(n_220),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_235),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_240),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_240),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_241),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_184),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_235),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_241),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_222),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_326),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_263),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_178),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_224),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_236),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_185),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_238),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_333),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_188),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_284),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_190),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_239),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_202),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_214),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_223),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_244),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_251),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_235),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_227),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_234),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_210),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_192),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_192),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_254),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_235),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_258),
.Y(n_433)
);

INVx4_ASAP7_75t_R g434 ( 
.A(n_226),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_237),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_179),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_194),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_401),
.A2(n_259),
.B1(n_197),
.B2(n_205),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_363),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_370),
.B(n_181),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_364),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_221),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_413),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_187),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_430),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_370),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_349),
.A2(n_265),
.B(n_253),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_352),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_363),
.B(n_176),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_368),
.B(n_176),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_370),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_359),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_359),
.B(n_181),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_348),
.B(n_187),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_374),
.B(n_208),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_428),
.A2(n_340),
.B1(n_335),
.B2(n_330),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_371),
.B(n_183),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_349),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_356),
.B(n_194),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_367),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_348),
.B(n_221),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_376),
.B(n_208),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_353),
.Y(n_476)
);

CKINVDCx6p67_ASAP7_75t_R g477 ( 
.A(n_374),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_353),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_365),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_354),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_354),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_225),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_357),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_357),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_358),
.Y(n_486)
);

CKINVDCx8_ASAP7_75t_R g487 ( 
.A(n_364),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_417),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_358),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_360),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_373),
.B(n_225),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_360),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_361),
.B(n_230),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_361),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_362),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_362),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_347),
.B(n_183),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_380),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_380),
.B(n_230),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_347),
.B(n_189),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_393),
.B(n_181),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_393),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_416),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_381),
.B(n_189),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_397),
.B(n_231),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_377),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_460),
.B(n_247),
.C(n_231),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_465),
.B(n_381),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_382),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_384),
.Y(n_521)
);

OAI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_497),
.A2(n_407),
.B1(n_429),
.B2(n_415),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_465),
.A2(n_394),
.B1(n_386),
.B2(n_389),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_375),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

AO22x1_ASAP7_75t_L g526 ( 
.A1(n_446),
.A2(n_366),
.B1(n_281),
.B2(n_288),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_498),
.Y(n_528)
);

CKINVDCx6p67_ASAP7_75t_R g529 ( 
.A(n_477),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_465),
.B(n_390),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_501),
.B(n_246),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_477),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_498),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_470),
.A2(n_433),
.B1(n_424),
.B2(n_405),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_498),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_500),
.B(n_409),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_502),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_444),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_502),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_481),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_502),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_503),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_500),
.B(n_410),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_446),
.B(n_414),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_460),
.A2(n_474),
.B1(n_438),
.B2(n_448),
.Y(n_546)
);

CKINVDCx6p67_ASAP7_75t_R g547 ( 
.A(n_477),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_489),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_490),
.A2(n_191),
.B(n_180),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_479),
.B(n_419),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_514),
.B(n_423),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_490),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_452),
.A2(n_402),
.B1(n_408),
.B2(n_320),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_474),
.B(n_431),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

AO22x1_ASAP7_75t_L g560 ( 
.A1(n_446),
.A2(n_342),
.B1(n_318),
.B2(n_273),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_447),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_446),
.B(n_233),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_466),
.B(n_351),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_443),
.B(n_350),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_496),
.B(n_298),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_509),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_443),
.B(n_402),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_452),
.B(n_355),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_445),
.A2(n_372),
.B1(n_398),
.B2(n_406),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_451),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_444),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_509),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_L g580 ( 
.A(n_454),
.B(n_399),
.C(n_397),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_445),
.A2(n_203),
.B1(n_198),
.B2(n_325),
.Y(n_581)
);

AND3x2_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_287),
.C(n_247),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g583 ( 
.A1(n_499),
.A2(n_329),
.B(n_287),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_469),
.Y(n_584)
);

CKINVDCx6p67_ASAP7_75t_R g585 ( 
.A(n_471),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_516),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_488),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_476),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_487),
.B(n_473),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_468),
.B(n_400),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_516),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_476),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_468),
.B(n_404),
.C(n_400),
.Y(n_595)
);

AOI21x1_ASAP7_75t_L g596 ( 
.A1(n_499),
.A2(n_329),
.B(n_196),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_501),
.B(n_246),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_473),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_462),
.B(n_261),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_480),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_480),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_480),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_450),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_447),
.Y(n_605)
);

BUFx16f_ASAP7_75t_R g606 ( 
.A(n_439),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_485),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_450),
.A2(n_493),
.B1(n_499),
.B2(n_462),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_485),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_484),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_488),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_447),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_462),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_485),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_466),
.B(n_193),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_507),
.A2(n_266),
.B1(n_270),
.B2(n_271),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_482),
.B(n_262),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_482),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_486),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_447),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_486),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_447),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_450),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_492),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_478),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_440),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_482),
.B(n_193),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_439),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_491),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_493),
.A2(n_276),
.B1(n_257),
.B2(n_246),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_491),
.B(n_404),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_512),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_501),
.B(n_246),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_493),
.A2(n_203),
.B1(n_198),
.B2(n_309),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_449),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_440),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_495),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_458),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_493),
.B(n_309),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_458),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_507),
.B(n_411),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_512),
.B(n_316),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_512),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_511),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_475),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_544),
.B(n_505),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_635),
.B(n_505),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_635),
.B(n_505),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_528),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_653),
.B(n_316),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_538),
.B(n_505),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_528),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_608),
.B(n_246),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_517),
.B(n_257),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_538),
.B(n_505),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_517),
.B(n_257),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_568),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_614),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_651),
.A2(n_515),
.B1(n_511),
.B2(n_274),
.C(n_319),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_652),
.Y(n_669)
);

O2A1O1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_598),
.A2(n_515),
.B(n_411),
.C(n_412),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_653),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_576),
.B(n_505),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_614),
.B(n_195),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_576),
.B(n_510),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_524),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_652),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_628),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_575),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_591),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_517),
.B(n_257),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_654),
.B(n_257),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_651),
.B(n_412),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_524),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_572),
.B(n_321),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_321),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_620),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_530),
.A2(n_286),
.B1(n_292),
.B2(n_296),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_620),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_611),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_644),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_644),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_551),
.B(n_418),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_637),
.B(n_420),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_654),
.B(n_276),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_558),
.B(n_325),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_533),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_520),
.B(n_521),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_533),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_541),
.B(n_548),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_541),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_649),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_535),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_555),
.B(n_510),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_555),
.B(n_527),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_646),
.Y(n_707)
);

AND2x6_ASAP7_75t_SL g708 ( 
.A(n_553),
.B(n_420),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_524),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_562),
.B(n_510),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_519),
.A2(n_297),
.B1(n_299),
.B2(n_300),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_SL g713 ( 
.A(n_568),
.B(n_604),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_SL g714 ( 
.A(n_590),
.B(n_205),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_535),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_524),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_570),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_604),
.A2(n_421),
.B(n_422),
.C(n_426),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_536),
.B(n_331),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_636),
.B(n_235),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_646),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_537),
.Y(n_723)
);

AOI221xp5_ASAP7_75t_L g724 ( 
.A1(n_632),
.A2(n_310),
.B1(n_312),
.B2(n_313),
.C(n_317),
.Y(n_724)
);

BUFx8_ASAP7_75t_L g725 ( 
.A(n_606),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_582),
.Y(n_726)
);

AOI22x1_ASAP7_75t_L g727 ( 
.A1(n_627),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_563),
.B(n_510),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_522),
.B(n_331),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_648),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_629),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_625),
.A2(n_550),
.B1(n_617),
.B2(n_637),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_600),
.B(n_619),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_537),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_539),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_629),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_625),
.B(n_276),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_574),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_567),
.B(n_332),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_637),
.B(n_421),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_580),
.B(n_422),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_630),
.B(n_510),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_575),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_539),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_630),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_631),
.B(n_332),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_634),
.B(n_640),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_642),
.B(n_336),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_640),
.B(n_276),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_561),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_550),
.A2(n_276),
.B1(n_305),
.B2(n_291),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_518),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_523),
.B(n_426),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_542),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_571),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_645),
.B(n_513),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_534),
.B(n_427),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_560),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_581),
.A2(n_272),
.B1(n_275),
.B2(n_268),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_595),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_650),
.B(n_336),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_542),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_543),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_526),
.B(n_219),
.C(n_218),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_632),
.A2(n_435),
.B(n_427),
.C(n_564),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_585),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_573),
.B(n_579),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_557),
.B(n_513),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_573),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_579),
.B(n_513),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_584),
.B(n_504),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_584),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_647),
.B(n_337),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_543),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_531),
.B(n_215),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_588),
.A2(n_435),
.B(n_603),
.C(n_626),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_588),
.B(n_504),
.Y(n_778)
);

BUFx5_ASAP7_75t_L g779 ( 
.A(n_593),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_593),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_552),
.B(n_337),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_526),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_602),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_618),
.B(n_343),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_599),
.B(n_601),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_532),
.B(n_343),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_615),
.A2(n_314),
.B(n_250),
.C(n_323),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_549),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_549),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_546),
.A2(n_344),
.B1(n_278),
.B2(n_285),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_554),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_623),
.A2(n_248),
.B1(n_345),
.B2(n_339),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_560),
.B(n_229),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_SL g794 ( 
.A1(n_611),
.A2(n_312),
.B1(n_310),
.B2(n_313),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_599),
.B(n_463),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_601),
.B(n_463),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_554),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_SL g798 ( 
.A(n_532),
.B(n_317),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_565),
.B(n_464),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_585),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_529),
.Y(n_801)
);

AND2x6_ASAP7_75t_L g802 ( 
.A(n_666),
.B(n_607),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_685),
.B(n_587),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_669),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_666),
.B(n_525),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_690),
.Y(n_806)
);

NOR2x1p5_ASAP7_75t_L g807 ( 
.A(n_801),
.B(n_547),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_734),
.B(n_699),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_699),
.B(n_609),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_667),
.B(n_561),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_680),
.B(n_616),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_683),
.B(n_547),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_697),
.A2(n_550),
.B1(n_610),
.B2(n_638),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_669),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_694),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_667),
.B(n_561),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_676),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_679),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_697),
.A2(n_525),
.B1(n_610),
.B2(n_638),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_666),
.B(n_616),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_671),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_621),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_731),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_732),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_701),
.B(n_703),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_737),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_752),
.A2(n_587),
.B1(n_327),
.B2(n_328),
.Y(n_827)
);

BUFx12f_ASAP7_75t_L g828 ( 
.A(n_767),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_751),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_746),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_686),
.A2(n_525),
.B1(n_610),
.B2(n_638),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_659),
.B(n_378),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_742),
.Y(n_833)
);

NOR2x2_ASAP7_75t_L g834 ( 
.A(n_794),
.B(n_434),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_692),
.B(n_621),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_378),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_677),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_662),
.A2(n_338),
.B1(n_306),
.B2(n_307),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_677),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_678),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_744),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_798),
.B(n_583),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_691),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_693),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_702),
.B(n_556),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_693),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_583),
.B(n_596),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_707),
.Y(n_848)
);

BUFx8_ASAP7_75t_SL g849 ( 
.A(n_800),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_721),
.Y(n_850)
);

AND2x2_ASAP7_75t_SL g851 ( 
.A(n_749),
.B(n_786),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_751),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_742),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_662),
.B(n_559),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_751),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_738),
.B(n_569),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_695),
.B(n_379),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_738),
.B(n_569),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_751),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_712),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_712),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_722),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_735),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_730),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_770),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_773),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_744),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_695),
.Y(n_868)
);

BUFx5_ASAP7_75t_L g869 ( 
.A(n_780),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_782),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_741),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_741),
.B(n_379),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_759),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_706),
.B(n_577),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_577),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_783),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_655),
.B(n_578),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_687),
.B(n_689),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_736),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_800),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_801),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_736),
.Y(n_882)
);

CKINVDCx11_ASAP7_75t_R g883 ( 
.A(n_708),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_718),
.B(n_779),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_753),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_718),
.B(n_578),
.Y(n_886)
);

AO22x1_ASAP7_75t_L g887 ( 
.A1(n_784),
.A2(n_328),
.B1(n_322),
.B2(n_327),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_660),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_769),
.A2(n_612),
.B1(n_566),
.B2(n_633),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_779),
.B(n_664),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_779),
.B(n_586),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_745),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_779),
.B(n_586),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_745),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_759),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_740),
.B(n_566),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_673),
.B(n_589),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_781),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_656),
.A2(n_441),
.B(n_613),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_713),
.B(n_566),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_755),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_740),
.B(n_594),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_761),
.B(n_594),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_R g904 ( 
.A(n_714),
.B(n_675),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_684),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_733),
.A2(n_589),
.B1(n_592),
.B2(n_305),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_726),
.B(n_799),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_779),
.B(n_592),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_769),
.A2(n_643),
.B1(n_594),
.B2(n_633),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_725),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_752),
.A2(n_733),
.B1(n_790),
.B2(n_766),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_779),
.B(n_605),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_663),
.A2(n_596),
.B(n_613),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_754),
.A2(n_784),
.B1(n_793),
.B2(n_760),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_719),
.A2(n_643),
.B1(n_605),
.B2(n_624),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_672),
.B(n_674),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_709),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_717),
.B(n_232),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_716),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_763),
.Y(n_920)
);

AOI211xp5_ASAP7_75t_L g921 ( 
.A1(n_724),
.A2(n_330),
.B(n_322),
.C(n_290),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_719),
.B(n_605),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_781),
.B(n_613),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_763),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_793),
.A2(n_305),
.B1(n_475),
.B2(n_501),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_756),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_739),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_758),
.Y(n_928)
);

NOR2x1_ASAP7_75t_R g929 ( 
.A(n_725),
.B(n_243),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_776),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_657),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_774),
.A2(n_762),
.B1(n_747),
.B2(n_720),
.Y(n_932)
);

INVx8_ASAP7_75t_L g933 ( 
.A(n_670),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_665),
.B(n_622),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_658),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_765),
.B(n_385),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_774),
.A2(n_643),
.B1(n_624),
.B2(n_641),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_661),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_665),
.B(n_467),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_762),
.A2(n_305),
.B1(n_501),
.B2(n_641),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_747),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_797),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_710),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_700),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_668),
.A2(n_305),
.B1(n_501),
.B2(n_597),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_729),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_705),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_704),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_681),
.B(n_467),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_729),
.B(n_385),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_682),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_715),
.Y(n_953)
);

AO22x1_ASAP7_75t_L g954 ( 
.A1(n_792),
.A2(n_289),
.B1(n_283),
.B2(n_282),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_681),
.A2(n_305),
.B1(n_501),
.B2(n_597),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_723),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_764),
.Y(n_957)
);

NOR3xp33_ASAP7_75t_SL g958 ( 
.A(n_787),
.B(n_255),
.C(n_249),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_777),
.B(n_387),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_775),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_768),
.B(n_472),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_711),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_788),
.B(n_789),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_791),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_688),
.B(n_441),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_776),
.A2(n_305),
.B1(n_501),
.B2(n_472),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_748),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_898),
.B(n_245),
.C(n_256),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_808),
.B(n_696),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_871),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_L g971 ( 
.A(n_803),
.B(n_696),
.C(n_787),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_851),
.B(n_260),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_L g973 ( 
.A(n_914),
.B(n_727),
.C(n_777),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_808),
.B(n_743),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_916),
.A2(n_771),
.B(n_757),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_804),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_932),
.A2(n_750),
.B1(n_785),
.B2(n_757),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_806),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_802),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_814),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_828),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_942),
.B(n_795),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_825),
.B(n_815),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_863),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_802),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_832),
.B(n_796),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_916),
.A2(n_772),
.B(n_778),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_815),
.B(n_387),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_836),
.B(n_750),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_871),
.B(n_279),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_829),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_867),
.B(n_388),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_911),
.A2(n_501),
.B1(n_305),
.B2(n_457),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_890),
.A2(n_449),
.B(n_455),
.Y(n_994)
);

BUFx2_ASAP7_75t_SL g995 ( 
.A(n_880),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_890),
.A2(n_449),
.B(n_455),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_859),
.A2(n_449),
.B(n_455),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_812),
.B(n_388),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_947),
.B(n_280),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_859),
.A2(n_449),
.B(n_455),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_806),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_911),
.A2(n_294),
.B(n_301),
.C(n_303),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_859),
.A2(n_449),
.B(n_455),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_817),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_859),
.A2(n_455),
.B(n_453),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_928),
.A2(n_346),
.B(n_391),
.C(n_392),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_877),
.A2(n_455),
.B(n_453),
.Y(n_1007)
);

OA22x2_ASAP7_75t_L g1008 ( 
.A1(n_927),
.A2(n_396),
.B1(n_392),
.B2(n_391),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_873),
.B(n_895),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_878),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_841),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_870),
.B(n_0),
.Y(n_1012)
);

OR2x4_ASAP7_75t_L g1013 ( 
.A(n_917),
.B(n_396),
.Y(n_1013)
);

AND2x4_ASAP7_75t_SL g1014 ( 
.A(n_868),
.B(n_860),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_930),
.A2(n_456),
.B1(n_459),
.B2(n_461),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_877),
.A2(n_809),
.B(n_912),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_833),
.Y(n_1017)
);

INVx6_ASAP7_75t_L g1018 ( 
.A(n_881),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_865),
.Y(n_1019)
);

OAI21xp33_ASAP7_75t_SL g1020 ( 
.A1(n_809),
.A2(n_0),
.B(n_2),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_912),
.A2(n_453),
.B(n_461),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_818),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_918),
.B(n_3),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_829),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_894),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_853),
.B(n_456),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_849),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_930),
.A2(n_461),
.B1(n_459),
.B2(n_453),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_866),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_852),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_965),
.A2(n_172),
.B(n_162),
.C(n_158),
.Y(n_1031)
);

AO22x2_ASAP7_75t_L g1032 ( 
.A1(n_827),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_962),
.A2(n_461),
.B(n_459),
.C(n_13),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_904),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_852),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_951),
.A2(n_459),
.B1(n_10),
.B2(n_15),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_885),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_857),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_857),
.B(n_9),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_926),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_876),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_821),
.B(n_145),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_852),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_872),
.B(n_141),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_891),
.A2(n_442),
.B(n_457),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_821),
.B(n_138),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_921),
.A2(n_18),
.B(n_19),
.C(n_23),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_893),
.A2(n_442),
.B(n_457),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_811),
.B(n_457),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_887),
.B(n_24),
.C(n_26),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_811),
.B(n_457),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_827),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_967),
.A2(n_74),
.B1(n_112),
.B2(n_109),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_951),
.B(n_31),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_908),
.A2(n_822),
.B(n_820),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_907),
.B(n_107),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_926),
.A2(n_31),
.B(n_35),
.C(n_36),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_855),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_822),
.A2(n_442),
.B(n_105),
.Y(n_1059)
);

INVx3_ASAP7_75t_SL g1060 ( 
.A(n_834),
.Y(n_1060)
);

INVx3_ASAP7_75t_SL g1061 ( 
.A(n_910),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_855),
.Y(n_1062)
);

AOI21x1_ASAP7_75t_L g1063 ( 
.A1(n_847),
.A2(n_922),
.B(n_923),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_951),
.B(n_35),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_936),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_899),
.A2(n_80),
.B(n_103),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_875),
.A2(n_442),
.B(n_68),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_SL g1068 ( 
.A1(n_905),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_948),
.B(n_442),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_936),
.A2(n_45),
.B(n_54),
.C(n_55),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_855),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_917),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_823),
.B(n_824),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_826),
.B(n_59),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_933),
.A2(n_59),
.B1(n_92),
.B2(n_93),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_936),
.A2(n_94),
.B(n_95),
.C(n_903),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_933),
.B(n_860),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_917),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_875),
.A2(n_805),
.B(n_934),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_907),
.B(n_830),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_805),
.A2(n_934),
.B(n_884),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_924),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_874),
.A2(n_896),
.B(n_902),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_952),
.A2(n_838),
.B(n_933),
.C(n_813),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_883),
.A2(n_872),
.B1(n_906),
.B2(n_941),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_874),
.A2(n_854),
.B(n_913),
.Y(n_1086)
);

AO22x1_ASAP7_75t_L g1087 ( 
.A1(n_861),
.A2(n_967),
.B1(n_862),
.B2(n_864),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_931),
.B(n_888),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_848),
.A2(n_850),
.B1(n_959),
.B2(n_944),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_961),
.B(n_944),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_861),
.B(n_807),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_924),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_958),
.A2(n_959),
.B(n_961),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_954),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_854),
.A2(n_858),
.B(n_856),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_919),
.B(n_943),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_967),
.A2(n_819),
.B1(n_861),
.B2(n_937),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_839),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_856),
.A2(n_858),
.B(n_967),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_831),
.A2(n_900),
.B1(n_915),
.B2(n_950),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_886),
.B(n_950),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1023),
.A2(n_919),
.B(n_897),
.C(n_940),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_979),
.B(n_949),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_983),
.B(n_835),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1093),
.A2(n_835),
.B(n_953),
.C(n_956),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_986),
.B(n_845),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1018),
.Y(n_1107)
);

AO21x1_ASAP7_75t_L g1108 ( 
.A1(n_1100),
.A2(n_810),
.B(n_816),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_1097),
.A2(n_844),
.A3(n_837),
.B(n_846),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1079),
.A2(n_900),
.B(n_949),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1055),
.A2(n_996),
.B(n_994),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_998),
.B(n_938),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_972),
.B(n_964),
.Y(n_1113)
);

OA21x2_ASAP7_75t_L g1114 ( 
.A1(n_1081),
.A2(n_843),
.B(n_963),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_974),
.B(n_839),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_991),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1068),
.A2(n_925),
.B1(n_946),
.B2(n_955),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1090),
.B(n_840),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1086),
.A2(n_909),
.B(n_889),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_988),
.B(n_1010),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_969),
.B(n_939),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1080),
.B(n_957),
.Y(n_1122)
);

CKINVDCx6p67_ASAP7_75t_R g1123 ( 
.A(n_1061),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_987),
.A2(n_1099),
.B(n_1087),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1073),
.B(n_945),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_SL g1127 ( 
.A(n_979),
.B(n_949),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_1001),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_991),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1091),
.B(n_960),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1063),
.A2(n_920),
.B(n_901),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1021),
.A2(n_879),
.B(n_882),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1039),
.B(n_964),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_973),
.A2(n_892),
.B(n_966),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_1084),
.A2(n_973),
.B(n_971),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1095),
.A2(n_935),
.B(n_869),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1019),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_L g1138 ( 
.A(n_1037),
.B(n_935),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1029),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1088),
.B(n_869),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_970),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1009),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1094),
.B(n_869),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1093),
.A2(n_802),
.B(n_869),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1041),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_999),
.C(n_1047),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1038),
.B(n_842),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_975),
.A2(n_1007),
.B(n_1066),
.Y(n_1148)
);

AOI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_1052),
.A2(n_949),
.B(n_929),
.Y(n_1149)
);

AOI221x1_ASAP7_75t_L g1150 ( 
.A1(n_1032),
.A2(n_1033),
.B1(n_1050),
.B2(n_1057),
.C(n_1040),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_979),
.A2(n_985),
.B(n_989),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_1018),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1096),
.B(n_1034),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1031),
.A2(n_977),
.B(n_1067),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1015),
.A2(n_1028),
.A3(n_1051),
.B(n_1049),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_970),
.Y(n_1156)
);

AOI211x1_ASAP7_75t_L g1157 ( 
.A1(n_1036),
.A2(n_1074),
.B(n_982),
.C(n_1056),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1059),
.A2(n_1048),
.A3(n_1045),
.B(n_976),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1017),
.B(n_1022),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_985),
.Y(n_1160)
);

OAI22x1_ASAP7_75t_L g1161 ( 
.A1(n_1012),
.A2(n_1060),
.B1(n_1054),
.B2(n_1064),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_977),
.A2(n_993),
.B(n_1076),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_980),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1026),
.A2(n_1069),
.B(n_1000),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1089),
.B(n_1044),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1044),
.B(n_1098),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1032),
.A2(n_1042),
.B1(n_993),
.B2(n_1091),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_984),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1065),
.A2(n_1070),
.B(n_1020),
.C(n_990),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1085),
.A2(n_1075),
.B1(n_1068),
.B2(n_1077),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_997),
.A2(n_1003),
.B(n_1005),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1020),
.A2(n_968),
.B(n_1092),
.C(n_1025),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_991),
.Y(n_1173)
);

NOR4xp25_ASAP7_75t_L g1174 ( 
.A(n_1053),
.B(n_1082),
.C(n_1024),
.D(n_1062),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1078),
.B(n_1085),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1072),
.B(n_1077),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1008),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_992),
.B(n_1078),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1077),
.A2(n_992),
.B(n_1062),
.Y(n_1179)
);

BUFx8_ASAP7_75t_L g1180 ( 
.A(n_1078),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1011),
.B(n_1030),
.C(n_1058),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_995),
.B(n_1046),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1030),
.A2(n_1035),
.B(n_1043),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1014),
.B(n_1071),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_981),
.A2(n_1030),
.B(n_1035),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1043),
.A2(n_1058),
.B(n_1071),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1027),
.A2(n_1100),
.A3(n_1083),
.B(n_1097),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1027),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1023),
.A2(n_808),
.B(n_932),
.C(n_914),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1016),
.A2(n_808),
.B(n_1083),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1023),
.A2(n_808),
.B1(n_851),
.B2(n_914),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1084),
.A2(n_808),
.B(n_1097),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_983),
.B(n_808),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1004),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_978),
.B(n_815),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_983),
.B(n_898),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_983),
.B(n_808),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_983),
.B(n_808),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1023),
.B(n_898),
.C(n_914),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1083),
.A2(n_808),
.B(n_1016),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1023),
.A2(n_808),
.B(n_932),
.C(n_914),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1037),
.B(n_671),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_991),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_978),
.B(n_815),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1091),
.B(n_1096),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1055),
.A2(n_996),
.B(n_994),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1023),
.B(n_685),
.C(n_914),
.Y(n_1207)
);

INVx6_ASAP7_75t_L g1208 ( 
.A(n_1018),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1023),
.B(n_898),
.C(n_914),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_983),
.B(n_808),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_970),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1083),
.A2(n_808),
.B(n_1016),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1004),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_979),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_978),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_983),
.B(n_808),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1027),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1023),
.A2(n_898),
.B1(n_803),
.B2(n_632),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1100),
.A2(n_1083),
.A3(n_1097),
.B(n_1081),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_983),
.B(n_808),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1016),
.A2(n_808),
.B(n_1083),
.Y(n_1221)
);

AOI31xp67_ASAP7_75t_L g1222 ( 
.A1(n_977),
.A2(n_813),
.A3(n_922),
.B(n_665),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_986),
.A2(n_808),
.B1(n_914),
.B2(n_932),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1004),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_978),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1097),
.A2(n_1079),
.B(n_1016),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1027),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1037),
.B(n_671),
.Y(n_1228)
);

NOR2xp67_ASAP7_75t_L g1229 ( 
.A(n_1037),
.B(n_671),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1004),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1004),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1083),
.A2(n_808),
.B(n_1016),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1023),
.A2(n_808),
.B(n_932),
.C(n_914),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1100),
.A2(n_1083),
.A3(n_1097),
.B(n_1081),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_R g1235 ( 
.A(n_1034),
.B(n_532),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1097),
.A2(n_1079),
.B(n_1016),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1013),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1016),
.A2(n_808),
.B(n_1083),
.Y(n_1238)
);

OAI22x1_ASAP7_75t_L g1239 ( 
.A1(n_1023),
.A2(n_898),
.B1(n_803),
.B2(n_632),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1023),
.A2(n_1032),
.B1(n_971),
.B2(n_911),
.C(n_1093),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1191),
.A2(n_1207),
.B1(n_1193),
.B2(n_1220),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1207),
.A2(n_1201),
.B(n_1189),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1120),
.B(n_1112),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1123),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_R g1245 ( 
.A(n_1235),
.B(n_1208),
.Y(n_1245)
);

AO21x2_ASAP7_75t_L g1246 ( 
.A1(n_1125),
.A2(n_1221),
.B(n_1190),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1110),
.A2(n_1236),
.B(n_1226),
.Y(n_1247)
);

NAND2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1214),
.B(n_1160),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1221),
.A2(n_1238),
.B(n_1162),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1179),
.B(n_1176),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1233),
.A2(n_1191),
.B(n_1162),
.C(n_1223),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1108),
.A2(n_1240),
.A3(n_1232),
.B(n_1212),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1132),
.A2(n_1164),
.B(n_1200),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1197),
.A2(n_1198),
.B1(n_1210),
.B2(n_1216),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1199),
.A2(n_1209),
.B1(n_1170),
.B2(n_1223),
.Y(n_1255)
);

OA21x2_ASAP7_75t_L g1256 ( 
.A1(n_1238),
.A2(n_1119),
.B(n_1101),
.Y(n_1256)
);

OAI222xp33_ASAP7_75t_L g1257 ( 
.A1(n_1170),
.A2(n_1196),
.B1(n_1175),
.B2(n_1165),
.C1(n_1177),
.C2(n_1128),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1214),
.B(n_1160),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1195),
.B(n_1204),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1142),
.A2(n_1104),
.B1(n_1113),
.B2(n_1157),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1150),
.A2(n_1105),
.B(n_1134),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1114),
.A2(n_1151),
.B(n_1134),
.Y(n_1262)
);

NAND2x1p5_ASAP7_75t_L g1263 ( 
.A(n_1214),
.B(n_1176),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1179),
.B(n_1192),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1128),
.B(n_1215),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1208),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1194),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1213),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1146),
.A2(n_1169),
.B(n_1102),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1141),
.B(n_1156),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1172),
.A2(n_1115),
.B(n_1121),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_SL g1272 ( 
.A1(n_1127),
.A2(n_1115),
.B(n_1106),
.Y(n_1272)
);

OAI222xp33_ASAP7_75t_L g1273 ( 
.A1(n_1215),
.A2(n_1122),
.B1(n_1153),
.B2(n_1225),
.C1(n_1124),
.C2(n_1147),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1166),
.B(n_1133),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1143),
.A2(n_1140),
.B(n_1118),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1222),
.A2(n_1163),
.B(n_1126),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1154),
.A2(n_1103),
.B(n_1186),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1149),
.B(n_1159),
.C(n_1229),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1174),
.A2(n_1145),
.B(n_1224),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1218),
.A2(n_1239),
.B1(n_1135),
.B2(n_1117),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1211),
.A2(n_1185),
.B(n_1230),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1211),
.A2(n_1185),
.B(n_1137),
.Y(n_1282)
);

NOR3xp33_ASAP7_75t_L g1283 ( 
.A(n_1149),
.B(n_1182),
.C(n_1117),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1139),
.A2(n_1231),
.B(n_1138),
.C(n_1168),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1109),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1161),
.A2(n_1205),
.B1(n_1228),
.B2(n_1202),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1178),
.A2(n_1184),
.B(n_1158),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1227),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1205),
.B(n_1152),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1167),
.A2(n_1234),
.A3(n_1219),
.B(n_1109),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1130),
.B(n_1152),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1181),
.A2(n_1107),
.B1(n_1217),
.B2(n_1188),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1219),
.A2(n_1234),
.B(n_1109),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1130),
.B(n_1237),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1180),
.Y(n_1296)
);

AOI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1187),
.A2(n_1155),
.B(n_1183),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1155),
.A2(n_1187),
.B(n_1183),
.C(n_1180),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_1187),
.A3(n_1129),
.B(n_1173),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1116),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1116),
.A2(n_1129),
.B(n_1173),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1116),
.A2(n_1129),
.B(n_1173),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1203),
.A2(n_1206),
.B(n_1111),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1203),
.A2(n_1136),
.B(n_1111),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1207),
.A2(n_1199),
.B1(n_1209),
.B2(n_851),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1191),
.A2(n_898),
.B1(n_808),
.B2(n_914),
.Y(n_1306)
);

INVx8_ASAP7_75t_L g1307 ( 
.A(n_1214),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1225),
.Y(n_1308)
);

AOI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1207),
.A2(n_685),
.B1(n_1209),
.B2(n_1199),
.C(n_898),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1144),
.B(n_1077),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1214),
.B(n_979),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1131),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1207),
.A2(n_1199),
.B1(n_1209),
.B2(n_851),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1131),
.Y(n_1314)
);

AOI222xp33_ASAP7_75t_L g1315 ( 
.A1(n_1199),
.A2(n_1068),
.B1(n_851),
.B2(n_439),
.C1(n_1209),
.C2(n_1207),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1214),
.B(n_979),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1179),
.B(n_1077),
.Y(n_1317)
);

OAI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1207),
.A2(n_914),
.B1(n_898),
.B2(n_685),
.C(n_1191),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1195),
.B(n_1204),
.Y(n_1319)
);

BUFx12f_ASAP7_75t_L g1320 ( 
.A(n_1237),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1207),
.A2(n_685),
.B(n_1189),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1214),
.Y(n_1322)
);

CKINVDCx8_ASAP7_75t_R g1323 ( 
.A(n_1188),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1208),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1208),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1148),
.A2(n_1206),
.B(n_1111),
.Y(n_1326)
);

NAND2x1p5_ASAP7_75t_L g1327 ( 
.A(n_1214),
.B(n_979),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1131),
.A2(n_1110),
.B(n_1171),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1148),
.A2(n_1206),
.B(n_1111),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1237),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1148),
.A2(n_1206),
.B(n_1111),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1148),
.A2(n_1206),
.B(n_1111),
.Y(n_1332)
);

AOI222xp33_ASAP7_75t_L g1333 ( 
.A1(n_1199),
.A2(n_1068),
.B1(n_851),
.B2(n_439),
.C1(n_1209),
.C2(n_1207),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1124),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1125),
.A2(n_1221),
.B(n_1190),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1109),
.Y(n_1336)
);

AO21x1_ASAP7_75t_L g1337 ( 
.A1(n_1223),
.A2(n_1023),
.B(n_1191),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1148),
.A2(n_1206),
.B(n_1111),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1120),
.B(n_1112),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1207),
.A2(n_1199),
.B1(n_1209),
.B2(n_851),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1188),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1195),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1207),
.A2(n_1199),
.B1(n_1209),
.B2(n_851),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1108),
.A2(n_1240),
.A3(n_1125),
.B(n_1212),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1189),
.A2(n_808),
.B(n_1233),
.C(n_1201),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1111),
.A2(n_1206),
.B(n_1238),
.Y(n_1346)
);

AND2x6_ASAP7_75t_L g1347 ( 
.A(n_1160),
.B(n_1177),
.Y(n_1347)
);

OAI221xp5_ASAP7_75t_L g1348 ( 
.A1(n_1207),
.A2(n_914),
.B1(n_898),
.B2(n_685),
.C(n_1191),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1144),
.B(n_1077),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1214),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1120),
.B(n_1112),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1179),
.B(n_1077),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1342),
.B(n_1254),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1269),
.A2(n_1306),
.B(n_1318),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1254),
.B(n_1259),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1285),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1348),
.A2(n_1321),
.B(n_1309),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1243),
.B(n_1339),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1255),
.A2(n_1280),
.B1(n_1313),
.B2(n_1305),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1351),
.B(n_1274),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1315),
.A2(n_1333),
.B(n_1257),
.C(n_1251),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1274),
.B(n_1283),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1289),
.B(n_1280),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1242),
.B(n_1308),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1241),
.B(n_1260),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1279),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_L g1367 ( 
.A(n_1278),
.B(n_1266),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1251),
.A2(n_1345),
.B(n_1337),
.C(n_1255),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1279),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1345),
.A2(n_1311),
.B(n_1316),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1324),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1266),
.B(n_1334),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1285),
.Y(n_1373)
);

AOI221x1_ASAP7_75t_SL g1374 ( 
.A1(n_1293),
.A2(n_1265),
.B1(n_1295),
.B2(n_1289),
.C(n_1267),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1324),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1305),
.A2(n_1313),
.B1(n_1340),
.B2(n_1343),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1265),
.B(n_1340),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1268),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1343),
.A2(n_1286),
.B1(n_1293),
.B2(n_1292),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1262),
.A2(n_1253),
.B(n_1247),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1311),
.A2(n_1316),
.B(n_1327),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1341),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1279),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1287),
.B(n_1264),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1317),
.B(n_1352),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1264),
.A2(n_1295),
.B1(n_1284),
.B2(n_1296),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1281),
.B(n_1282),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1299),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1245),
.Y(n_1389)
);

O2A1O1Ixp5_ASAP7_75t_L g1390 ( 
.A1(n_1297),
.A2(n_1290),
.B(n_1328),
.C(n_1273),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1298),
.A2(n_1272),
.B(n_1261),
.C(n_1336),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1310),
.A2(n_1349),
.B1(n_1263),
.B2(n_1261),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1287),
.B(n_1271),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1300),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1299),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_1248),
.B1(n_1258),
.B2(n_1271),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1248),
.A2(n_1258),
.B1(n_1270),
.B2(n_1325),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1302),
.B(n_1301),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1347),
.B(n_1249),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1245),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1281),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1270),
.A2(n_1330),
.B1(n_1320),
.B2(n_1350),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1320),
.A2(n_1330),
.B1(n_1350),
.B2(n_1322),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1256),
.A2(n_1307),
.B1(n_1275),
.B2(n_1276),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1282),
.B(n_1347),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1301),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_SL g1408 ( 
.A1(n_1344),
.A2(n_1252),
.B(n_1291),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1347),
.B(n_1256),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1275),
.B(n_1291),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1246),
.A2(n_1335),
.B(n_1314),
.C(n_1312),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1307),
.A2(n_1276),
.B1(n_1294),
.B2(n_1312),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1252),
.A2(n_1291),
.B(n_1294),
.C(n_1277),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1288),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1303),
.A2(n_1346),
.B(n_1288),
.C(n_1277),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1326),
.A2(n_1329),
.B(n_1331),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1329),
.A2(n_1331),
.B(n_1332),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1304),
.A2(n_1209),
.B(n_1199),
.C(n_1201),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1338),
.B(n_1243),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1285),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1324),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1243),
.B(n_1339),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1342),
.B(n_1254),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1243),
.B(n_1339),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1243),
.B(n_1339),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1269),
.A2(n_1207),
.B(n_1023),
.C(n_803),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_SL g1428 ( 
.A1(n_1280),
.A2(n_898),
.B1(n_851),
.B2(n_1068),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1259),
.B(n_1319),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1250),
.B(n_1317),
.Y(n_1430)
);

O2A1O1Ixp5_ASAP7_75t_L g1431 ( 
.A1(n_1269),
.A2(n_1337),
.B(n_1321),
.C(n_1207),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1342),
.B(n_1254),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1255),
.A2(n_898),
.B1(n_851),
.B2(n_1191),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1255),
.A2(n_898),
.B1(n_851),
.B2(n_1191),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1419),
.B(n_1366),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1426),
.B(n_1376),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1355),
.B(n_1365),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1369),
.B(n_1383),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1387),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1356),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1373),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1420),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1382),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1353),
.B(n_1423),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1406),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1393),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1368),
.B(n_1361),
.Y(n_1447)
);

INVxp33_ASAP7_75t_L g1448 ( 
.A(n_1360),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1367),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1407),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1384),
.B(n_1405),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1400),
.B(n_1409),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1399),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1402),
.B(n_1413),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1412),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1413),
.B(n_1430),
.Y(n_1456)
);

INVx5_ASAP7_75t_L g1457 ( 
.A(n_1385),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1429),
.Y(n_1458)
);

INVxp67_ASAP7_75t_L g1459 ( 
.A(n_1364),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1388),
.B(n_1395),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1432),
.B(n_1362),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1378),
.B(n_1377),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1415),
.A2(n_1411),
.B(n_1391),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1359),
.A2(n_1434),
.B1(n_1433),
.B2(n_1428),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1390),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1390),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1392),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1416),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1363),
.Y(n_1469)
);

OR2x2_ASAP7_75t_SL g1470 ( 
.A(n_1357),
.B(n_1354),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1470),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1436),
.B(n_1379),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1446),
.B(n_1417),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1452),
.B(n_1368),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1450),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1469),
.B(n_1431),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1358),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1470),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1470),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1435),
.B(n_1456),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1436),
.A2(n_1361),
.B1(n_1422),
.B2(n_1425),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1435),
.B(n_1456),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1468),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.B(n_1424),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1451),
.B(n_1386),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1451),
.B(n_1394),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1438),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1396),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1455),
.B(n_1408),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1468),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1418),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1483),
.Y(n_1494)
);

AO21x1_ASAP7_75t_SL g1495 ( 
.A1(n_1493),
.A2(n_1467),
.B(n_1466),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1487),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1475),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1472),
.A2(n_1464),
.B1(n_1447),
.B2(n_1437),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1487),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1465),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1492),
.Y(n_1501)
);

NOR3xp33_ASAP7_75t_L g1502 ( 
.A(n_1472),
.B(n_1447),
.C(n_1464),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1481),
.A2(n_1437),
.B1(n_1461),
.B2(n_1458),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1475),
.Y(n_1504)
);

OAI211xp5_ASAP7_75t_L g1505 ( 
.A1(n_1481),
.A2(n_1444),
.B(n_1461),
.C(n_1465),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1471),
.B(n_1457),
.Y(n_1506)
);

OAI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1493),
.A2(n_1444),
.B1(n_1389),
.B2(n_1467),
.C(n_1466),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1491),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1453),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1471),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1488),
.A2(n_1474),
.B1(n_1485),
.B2(n_1489),
.C(n_1479),
.Y(n_1512)
);

AOI211xp5_ASAP7_75t_L g1513 ( 
.A1(n_1488),
.A2(n_1403),
.B(n_1404),
.C(n_1370),
.Y(n_1513)
);

OA222x2_ASAP7_75t_L g1514 ( 
.A1(n_1485),
.A2(n_1460),
.B1(n_1462),
.B2(n_1441),
.C1(n_1442),
.C2(n_1440),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1476),
.B(n_1440),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1454),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1486),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1471),
.A2(n_1458),
.B1(n_1463),
.B2(n_1448),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1474),
.A2(n_1448),
.B1(n_1462),
.B2(n_1449),
.Y(n_1519)
);

INVx3_ASAP7_75t_SL g1520 ( 
.A(n_1490),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1478),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1519),
.B(n_1478),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1497),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1497),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1504),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1515),
.B(n_1476),
.Y(n_1526)
);

INVx4_ASAP7_75t_L g1527 ( 
.A(n_1511),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1516),
.B(n_1482),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

NAND4xp25_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1476),
.C(n_1478),
.D(n_1479),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1500),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_L g1533 ( 
.A(n_1502),
.B(n_1490),
.C(n_1489),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1473),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1496),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1508),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1509),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1496),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1499),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1499),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1508),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1515),
.B(n_1484),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1506),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1482),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1506),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1508),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1506),
.B(n_1478),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1494),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1526),
.B(n_1517),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1535),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1537),
.B(n_1509),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1535),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1414),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1549),
.B(n_1501),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1531),
.B(n_1443),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1539),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_SL g1564 ( 
.A(n_1533),
.B(n_1512),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1533),
.B(n_1484),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1537),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1523),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1539),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1537),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.B(n_1517),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1549),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1540),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1523),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1542),
.B(n_1519),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1549),
.B(n_1520),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1522),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1527),
.B(n_1503),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1529),
.B(n_1544),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1520),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1527),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_SL g1586 ( 
.A(n_1527),
.B(n_1495),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1524),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1530),
.B(n_1509),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1520),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1530),
.A2(n_1498),
.B1(n_1505),
.B2(n_1479),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1525),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1532),
.A2(n_1512),
.B1(n_1498),
.B2(n_1507),
.C(n_1505),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1525),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1568),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1503),
.Y(n_1595)
);

NAND2xp33_ASAP7_75t_L g1596 ( 
.A(n_1590),
.B(n_1401),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1586),
.B(n_1543),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1566),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1565),
.B(n_1528),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1592),
.B(n_1527),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1581),
.B(n_1582),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1571),
.B(n_1530),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1593),
.Y(n_1604)
);

INVxp33_ASAP7_75t_L g1605 ( 
.A(n_1557),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1588),
.B(n_1530),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1584),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1579),
.B(n_1507),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1588),
.B(n_1530),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1586),
.B(n_1543),
.Y(n_1610)
);

AO22x1_ASAP7_75t_L g1611 ( 
.A1(n_1588),
.A2(n_1521),
.B1(n_1509),
.B2(n_1511),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1554),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1555),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1559),
.A2(n_1518),
.B(n_1513),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1556),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1516),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1556),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1552),
.B(n_1528),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1521),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1562),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1567),
.B(n_1477),
.Y(n_1623)
);

INVxp33_ASAP7_75t_L g1624 ( 
.A(n_1555),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1543),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1562),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1543),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1552),
.B(n_1534),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1572),
.B(n_1534),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1606),
.A2(n_1580),
.B(n_1589),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1607),
.B(n_1555),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1595),
.A2(n_1518),
.B1(n_1479),
.B2(n_1485),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1599),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1613),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1614),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1596),
.A2(n_1573),
.B1(n_1553),
.B2(n_1558),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1604),
.B(n_1585),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1601),
.A2(n_1463),
.B1(n_1591),
.B2(n_1578),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1607),
.B(n_1583),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1617),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1619),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1622),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1612),
.B(n_1560),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1573),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1596),
.A2(n_1605),
.B1(n_1594),
.B2(n_1612),
.C1(n_1615),
.C2(n_1624),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1560),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1583),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1626),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1609),
.B(n_1578),
.Y(n_1652)
);

AND3x1_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1513),
.C(n_1551),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1654)
);

AOI222xp33_ASAP7_75t_L g1655 ( 
.A1(n_1603),
.A2(n_1532),
.B1(n_1558),
.B2(n_1551),
.C1(n_1553),
.C2(n_1569),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1656),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1637),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1634),
.A2(n_1511),
.B1(n_1606),
.B2(n_1600),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1637),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1635),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1632),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1648),
.A2(n_1621),
.B(n_1597),
.C(n_1610),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1647),
.B(n_1620),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1654),
.B(n_1600),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1642),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1638),
.A2(n_1625),
.B1(n_1627),
.B2(n_1610),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1644),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1643),
.B(n_1628),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1654),
.B(n_1625),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1645),
.Y(n_1675)
);

OAI211xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1640),
.A2(n_1629),
.B(n_1628),
.C(n_1618),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1672),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1666),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1652),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1639),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1657),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1663),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1662),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1673),
.B(n_1630),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1665),
.Y(n_1686)
);

AND2x4_ASAP7_75t_SL g1687 ( 
.A(n_1661),
.B(n_1630),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1669),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1671),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1675),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1677),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_SL g1692 ( 
.A(n_1679),
.B(n_1670),
.C(n_1640),
.Y(n_1692)
);

OAI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1685),
.A2(n_1676),
.B(n_1664),
.C(n_1668),
.Y(n_1693)
);

NAND4xp25_ASAP7_75t_L g1694 ( 
.A(n_1683),
.B(n_1674),
.C(n_1655),
.D(n_1676),
.Y(n_1694)
);

O2A1O1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1688),
.A2(n_1659),
.B(n_1633),
.C(n_1630),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1688),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1678),
.B(n_1659),
.C(n_1633),
.Y(n_1697)
);

OAI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1683),
.A2(n_1631),
.B(n_1597),
.C(n_1649),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1680),
.B(n_1641),
.Y(n_1699)
);

O2A1O1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1680),
.A2(n_1646),
.B(n_1629),
.C(n_1545),
.Y(n_1700)
);

NAND5xp2_ASAP7_75t_SL g1701 ( 
.A(n_1687),
.B(n_1631),
.C(n_1611),
.D(n_1514),
.E(n_1510),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1681),
.A2(n_1545),
.B1(n_1521),
.B2(n_1511),
.C(n_1506),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1696),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1699),
.Y(n_1704)
);

OAI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1695),
.A2(n_1693),
.B(n_1692),
.C(n_1694),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1697),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1701),
.A2(n_1680),
.B1(n_1682),
.B2(n_1690),
.C(n_1691),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1698),
.A2(n_1687),
.B1(n_1690),
.B2(n_1702),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1703),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1704),
.B(n_1690),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1708),
.B(n_1684),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1706),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1705),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1707),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1703),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1710),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1710),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1709),
.Y(n_1718)
);

XNOR2xp5_ASAP7_75t_L g1719 ( 
.A(n_1714),
.B(n_1686),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1713),
.A2(n_1689),
.B1(n_1545),
.B2(n_1569),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1711),
.B(n_1623),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1718),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1712),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1717),
.B(n_1709),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1722),
.Y(n_1725)
);

OAI322xp33_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1720),
.A3(n_1724),
.B1(n_1715),
.B2(n_1719),
.C1(n_1718),
.C2(n_1721),
.Y(n_1726)
);

XNOR2xp5_ASAP7_75t_L g1727 ( 
.A(n_1726),
.B(n_1723),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1726),
.A2(n_1700),
.B1(n_1563),
.B2(n_1570),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1727),
.Y(n_1729)
);

XNOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_1728),
.B(n_1375),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1730),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1729),
.A2(n_1397),
.B1(n_1427),
.B2(n_1421),
.Y(n_1732)
);

AOI222xp33_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1570),
.B1(n_1563),
.B2(n_1574),
.C1(n_1561),
.C2(n_1575),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1733),
.B(n_1731),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1734),
.B(n_1371),
.Y(n_1735)
);

AOI322xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1521),
.A3(n_1536),
.B1(n_1548),
.B2(n_1541),
.C1(n_1546),
.C2(n_1547),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1736),
.A2(n_1372),
.B1(n_1550),
.B2(n_1547),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1398),
.B(n_1381),
.C(n_1534),
.Y(n_1738)
);


endmodule