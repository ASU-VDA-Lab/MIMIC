module fake_netlist_5_2511_n_1705 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1705);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1705;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_48),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_29),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_29),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_92),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_25),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_40),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_51),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_49),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_123),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_20),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_14),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_23),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_58),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_21),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_65),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_87),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_22),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_79),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_85),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_14),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_72),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_56),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_31),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_63),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_5),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_8),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_34),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_66),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_137),
.Y(n_211)
);

BUFx10_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_113),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_122),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_36),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_33),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_32),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_5),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_42),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_17),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_110),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_90),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_94),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_30),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_121),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_148),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_88),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_101),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_126),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_9),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_91),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_37),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_59),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_49),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_45),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_13),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_127),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_13),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_84),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_115),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_102),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_30),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_104),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_7),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_3),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_147),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_71),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_61),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_76),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_34),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_130),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_103),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_51),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_81),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_12),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_58),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_134),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_19),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_116),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_39),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_68),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_46),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_48),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_46),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_119),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_32),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_73),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_23),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_53),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_108),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_35),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_225),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_164),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_184),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_209),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_190),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_234),
.B(n_1),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_243),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_244),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_248),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_190),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_190),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_190),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_166),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_190),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_190),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_177),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_227),
.B(n_1),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_179),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_181),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_185),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_277),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_245),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_189),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_250),
.B(n_2),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_277),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_232),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_192),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_171),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_171),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_175),
.B(n_2),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_196),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_229),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_R g353 ( 
.A(n_201),
.B(n_211),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_213),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_215),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_216),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_229),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_222),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_226),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_247),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_232),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_256),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_253),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_210),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_256),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

BUFx6f_ASAP7_75t_SL g369 ( 
.A(n_212),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_254),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_258),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_259),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_265),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_273),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_274),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_275),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_204),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_269),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_278),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_286),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_204),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_198),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

CKINVDCx6p67_ASAP7_75t_R g387 ( 
.A(n_316),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_366),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_159),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_340),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_313),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_331),
.A2(n_269),
.B(n_165),
.Y(n_397)
);

CKINVDCx8_ASAP7_75t_R g398 ( 
.A(n_345),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_183),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_331),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_157),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_340),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_335),
.B(n_167),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_353),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_336),
.B(n_167),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_319),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_337),
.A2(n_165),
.B(n_156),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_310),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_339),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_342),
.B(n_290),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_342),
.B(n_159),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_319),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_321),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_344),
.Y(n_428)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_345),
.A2(n_297),
.B1(n_287),
.B2(n_252),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_322),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_314),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g433 ( 
.A(n_326),
.B(n_186),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_328),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_323),
.B(n_186),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_324),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_324),
.B(n_160),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_343),
.A2(n_252),
.B1(n_207),
.B2(n_307),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_330),
.B(n_188),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_325),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_325),
.B(n_348),
.Y(n_443)
);

BUFx8_ASAP7_75t_L g444 ( 
.A(n_369),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_349),
.B(n_292),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_352),
.B(n_160),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_327),
.B(n_212),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_395),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_394),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_401),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_172),
.C(n_169),
.Y(n_456)
);

OR2x6_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_169),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_441),
.B(n_332),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

OR2x6_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_172),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_397),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_401),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_394),
.B(n_364),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_401),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_394),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_365),
.B1(n_347),
.B2(n_351),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_397),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_396),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_443),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_441),
.B(n_355),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_413),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_416),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_405),
.B(n_360),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_410),
.B(n_372),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_384),
.B(n_364),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_402),
.Y(n_489)
);

AND2x2_ASAP7_75t_SL g490 ( 
.A(n_416),
.B(n_280),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_440),
.A2(n_207),
.B1(n_170),
.B2(n_194),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

NOR2x1p5_ASAP7_75t_L g493 ( 
.A(n_387),
.B(n_311),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_432),
.A2(n_219),
.B1(n_193),
.B2(n_180),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_373),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_433),
.B(n_375),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_387),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_384),
.B(n_367),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g502 ( 
.A(n_416),
.B(n_280),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_427),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_384),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_449),
.B(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_390),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_449),
.B(n_367),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_396),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_435),
.B(n_379),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_417),
.B(n_382),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_437),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_417),
.B(n_383),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_399),
.B(n_191),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_399),
.B(n_293),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_449),
.B(n_381),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_439),
.B(n_176),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_388),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_407),
.B(n_421),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_406),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_414),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_388),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_396),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_306),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_396),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_425),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_424),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_427),
.Y(n_545)
);

OAI22xp33_ASAP7_75t_L g546 ( 
.A1(n_419),
.A2(n_260),
.B1(n_173),
.B2(n_168),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_396),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_413),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_385),
.B(n_341),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_439),
.B(n_302),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_430),
.B(n_309),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_385),
.B(n_176),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_413),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_L g556 ( 
.A1(n_419),
.A2(n_240),
.B1(n_238),
.B2(n_237),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_439),
.B(n_178),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_416),
.B(n_182),
.C(n_178),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_389),
.B(n_354),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_387),
.Y(n_561)
);

OAI22xp33_ASAP7_75t_L g562 ( 
.A1(n_433),
.A2(n_206),
.B1(n_228),
.B2(n_220),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_389),
.B(n_356),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_413),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_416),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_415),
.B(n_182),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_415),
.B(n_203),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_388),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_392),
.A2(n_156),
.B1(n_170),
.B2(n_261),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_438),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_444),
.B(n_359),
.Y(n_575)
);

NAND3xp33_ASAP7_75t_L g576 ( 
.A(n_422),
.B(n_246),
.C(n_203),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_395),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_447),
.B(n_361),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_438),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_392),
.B(n_381),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_415),
.B(n_447),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_442),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_444),
.B(n_362),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_450),
.B(n_370),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_422),
.B(n_302),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_386),
.B(n_338),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_442),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_422),
.B(n_368),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_436),
.B(n_208),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_436),
.A2(n_200),
.B1(n_242),
.B2(n_261),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_436),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_387),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_395),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_436),
.A2(n_199),
.B1(n_200),
.B2(n_285),
.Y(n_601)
);

BUFx8_ASAP7_75t_L g602 ( 
.A(n_527),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_504),
.B(n_509),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_476),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_528),
.B(n_436),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_506),
.B(n_436),
.Y(n_606)
);

BUFx6f_ASAP7_75t_SL g607 ( 
.A(n_480),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_506),
.B(n_431),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_478),
.B(n_508),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_508),
.B(n_386),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_431),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_490),
.B(n_398),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_490),
.B(n_398),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_454),
.B(n_424),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_490),
.B(n_398),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_464),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_551),
.B(n_376),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_431),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_484),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_463),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_592),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_531),
.B(n_431),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_464),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_518),
.B(n_377),
.Y(n_627)
);

NOR2x1p5_ASAP7_75t_L g628 ( 
.A(n_561),
.B(n_187),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_479),
.B(n_431),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_520),
.B(n_431),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_485),
.B(n_378),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_487),
.B(n_424),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_495),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_502),
.B(n_431),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_581),
.A2(n_315),
.B1(n_317),
.B2(n_450),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_527),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_598),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_502),
.B(n_429),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_429),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_592),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_495),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_454),
.B(n_429),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_484),
.B(n_398),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_467),
.B(n_429),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_429),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_598),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_484),
.B(n_221),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_540),
.B(n_429),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_503),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_503),
.B(n_510),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_590),
.A2(n_430),
.B1(n_409),
.B2(n_412),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_457),
.A2(n_409),
.B1(n_412),
.B2(n_369),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_468),
.B(n_158),
.C(n_155),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_487),
.B(n_451),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_497),
.B(n_369),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_573),
.B(n_264),
.C(n_162),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

A2O1A1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_456),
.A2(n_223),
.B(n_307),
.C(n_304),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_529),
.B(n_221),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_553),
.A2(n_163),
.B1(n_161),
.B2(n_202),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_463),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_560),
.B(n_564),
.C(n_562),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_510),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_458),
.B(n_205),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_516),
.B(n_231),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_511),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_524),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_522),
.B(n_255),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_524),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_529),
.B(n_221),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_457),
.A2(n_409),
.B1(n_412),
.B2(n_262),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_552),
.B(n_221),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_395),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_595),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_517),
.Y(n_676)
);

XOR2xp5_ASAP7_75t_L g677 ( 
.A(n_553),
.B(n_505),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_486),
.B(n_514),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_523),
.B(n_395),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_457),
.A2(n_412),
.B1(n_409),
.B2(n_224),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_512),
.A2(n_409),
.B(n_412),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_529),
.A2(n_409),
.B1(n_412),
.B2(n_239),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_L g684 ( 
.A(n_552),
.B(n_221),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_567),
.B(n_236),
.Y(n_685)
);

O2A1O1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_557),
.A2(n_223),
.B(n_304),
.C(n_194),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_501),
.B(n_583),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_523),
.B(n_391),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_526),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_544),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_526),
.B(n_391),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_567),
.B(n_236),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_525),
.B(n_391),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_393),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_567),
.B(n_236),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_501),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_572),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_525),
.B(n_393),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_494),
.B(n_266),
.Y(n_700)
);

AO22x2_ASAP7_75t_L g701 ( 
.A1(n_456),
.A2(n_559),
.B1(n_576),
.B2(n_575),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_583),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_525),
.B(n_393),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_559),
.A2(n_214),
.B1(n_208),
.B2(n_224),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_461),
.B(n_400),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_572),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_469),
.B(n_400),
.Y(n_707)
);

AND2x6_ASAP7_75t_SL g708 ( 
.A(n_457),
.B(n_174),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_480),
.B(n_444),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_552),
.A2(n_591),
.B1(n_463),
.B2(n_469),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_471),
.B(n_403),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_471),
.B(n_403),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_472),
.A2(n_423),
.B(n_408),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_472),
.B(n_403),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_457),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_588),
.B(n_214),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_473),
.B(n_236),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_473),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_571),
.B(n_404),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_571),
.Y(n_721)
);

NOR2xp67_ASAP7_75t_L g722 ( 
.A(n_599),
.B(n_451),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_596),
.Y(n_723)
);

XNOR2x2_ASAP7_75t_SL g724 ( 
.A(n_576),
.B(n_174),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_460),
.B(n_404),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_569),
.Y(n_726)
);

INVxp33_ASAP7_75t_L g727 ( 
.A(n_554),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_455),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_460),
.B(n_404),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_570),
.A2(n_483),
.B(n_466),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_532),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_460),
.B(n_408),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_SL g733 ( 
.A(n_491),
.B(n_233),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_455),
.Y(n_734)
);

AND2x2_ASAP7_75t_SL g735 ( 
.A(n_498),
.B(n_235),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_460),
.B(n_271),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_SL g737 ( 
.A(n_474),
.B(n_236),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_474),
.B(n_444),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_460),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_459),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_546),
.B(n_272),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_459),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_556),
.B(n_279),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_552),
.B(n_408),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_552),
.B(n_591),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_411),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_474),
.B(n_444),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_597),
.A2(n_283),
.B1(n_288),
.B2(n_235),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_532),
.A2(n_582),
.B(n_533),
.C(n_534),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_462),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_591),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_533),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_534),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_466),
.A2(n_420),
.B(n_423),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_474),
.B(n_444),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_462),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_465),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_474),
.B(n_446),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_591),
.B(n_411),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_545),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_480),
.B(n_282),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_591),
.A2(n_241),
.B1(n_267),
.B2(n_270),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_535),
.A2(n_411),
.B(n_418),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_480),
.B(n_470),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_453),
.B(n_451),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_591),
.B(n_418),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_591),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_535),
.A2(n_251),
.B1(n_262),
.B2(n_239),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_536),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_493),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_499),
.A2(n_289),
.B1(n_291),
.B2(n_295),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_609),
.B(n_466),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_632),
.B(n_610),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_727),
.B(n_470),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_669),
.B(n_466),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_690),
.Y(n_776)
);

AOI21xp33_ASAP7_75t_L g777 ( 
.A1(n_627),
.A2(n_601),
.B(n_246),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_664),
.A2(n_249),
.B(n_241),
.C(n_299),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_604),
.B(n_483),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_604),
.B(n_483),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_643),
.A2(n_536),
.B(n_542),
.C(n_589),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_727),
.B(n_470),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_634),
.A2(n_481),
.B(n_470),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_704),
.A2(n_733),
.B1(n_719),
.B2(n_611),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_605),
.A2(n_548),
.B(n_530),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_710),
.A2(n_586),
.B1(n_493),
.B2(n_299),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_603),
.B(n_474),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

NAND2x1_ASAP7_75t_L g789 ( 
.A(n_623),
.B(n_483),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_607),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_641),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_647),
.A2(n_542),
.B(n_549),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_643),
.A2(n_549),
.B(n_550),
.C(n_589),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_638),
.A2(n_548),
.B(n_530),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_611),
.B(n_521),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_717),
.A2(n_550),
.B(n_563),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_641),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_613),
.B(n_521),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_717),
.A2(n_563),
.B(n_574),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_639),
.A2(n_530),
.B(n_548),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_662),
.A2(n_541),
.B1(n_521),
.B2(n_539),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_718),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_649),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_632),
.B(n_257),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

AO21x1_ASAP7_75t_L g806 ( 
.A1(n_647),
.A2(n_281),
.B(n_249),
.Y(n_806)
);

OAI21xp33_ASAP7_75t_L g807 ( 
.A1(n_700),
.A2(n_300),
.B(n_301),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_648),
.A2(n_530),
.B(n_548),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_617),
.B(n_539),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_640),
.B(n_481),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_614),
.A2(n_547),
.B1(n_541),
.B2(n_539),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_612),
.A2(n_537),
.B(n_481),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_702),
.A2(n_578),
.B(n_580),
.C(n_587),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_663),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_617),
.B(n_539),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_665),
.A2(n_251),
.B(n_270),
.C(n_288),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_635),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_706),
.B(n_267),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_687),
.B(n_482),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_726),
.B(n_541),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_741),
.A2(n_743),
.B(n_610),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_631),
.B(n_481),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_654),
.B(n_541),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_642),
.A2(n_537),
.B(n_482),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_736),
.A2(n_547),
.B(n_580),
.C(n_587),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_644),
.A2(n_645),
.B(n_630),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_L g827 ( 
.A1(n_620),
.A2(n_303),
.B(n_199),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_659),
.A2(n_582),
.B(n_584),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_702),
.A2(n_584),
.B(n_594),
.C(n_488),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_654),
.B(n_547),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_663),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_659),
.A2(n_507),
.B(n_594),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_676),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_679),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_676),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_671),
.A2(n_543),
.B(n_492),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_771),
.B(n_197),
.C(n_218),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_671),
.A2(n_543),
.B(n_492),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_619),
.A2(n_500),
.B(n_465),
.C(n_488),
.Y(n_839)
);

AO21x2_ASAP7_75t_L g840 ( 
.A1(n_685),
.A2(n_558),
.B(n_500),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_739),
.A2(n_586),
.B1(n_482),
.B2(n_555),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_624),
.B(n_537),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_619),
.B(n_257),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_685),
.A2(n_489),
.B(n_496),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_739),
.A2(n_586),
.B1(n_482),
.B2(n_555),
.Y(n_845)
);

INVx4_ASAP7_75t_L g846 ( 
.A(n_623),
.Y(n_846)
);

AOI22x1_ASAP7_75t_L g847 ( 
.A1(n_701),
.A2(n_565),
.B1(n_555),
.B2(n_537),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_705),
.A2(n_558),
.B(n_489),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_626),
.A2(n_515),
.B(n_496),
.C(n_568),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_706),
.B(n_565),
.Y(n_850)
);

AOI21x1_ASAP7_75t_L g851 ( 
.A1(n_707),
.A2(n_568),
.B(n_515),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_657),
.B(n_452),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_673),
.A2(n_482),
.B(n_577),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_689),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_673),
.A2(n_577),
.B(n_565),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_684),
.A2(n_577),
.B(n_565),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_711),
.A2(n_507),
.B(n_566),
.Y(n_857)
);

OAI321xp33_ASAP7_75t_L g858 ( 
.A1(n_651),
.A2(n_197),
.A3(n_242),
.B1(n_230),
.B2(n_218),
.C(n_294),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_723),
.B(n_566),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_679),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_614),
.A2(n_600),
.B1(n_453),
.B2(n_579),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_719),
.B(n_577),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_636),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_668),
.B(n_678),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_L g865 ( 
.A(n_653),
.B(n_298),
.C(n_230),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_718),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_760),
.B(n_453),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_684),
.A2(n_577),
.B(n_593),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_606),
.B(n_577),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_622),
.B(n_519),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_622),
.A2(n_600),
.B(n_579),
.C(n_519),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_745),
.A2(n_593),
.B(n_513),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_637),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_728),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_622),
.A2(n_696),
.B(n_692),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_767),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_692),
.A2(n_593),
.B(n_513),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_697),
.B(n_519),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_698),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_696),
.A2(n_600),
.B(n_579),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_608),
.A2(n_593),
.B(n_513),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_666),
.B(n_418),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_682),
.A2(n_593),
.B(n_513),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_623),
.A2(n_423),
.B1(n_420),
.B2(n_428),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_667),
.B(n_420),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_L g886 ( 
.A(n_761),
.B(n_298),
.C(n_284),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_621),
.A2(n_593),
.B(n_513),
.Y(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_661),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_661),
.Y(n_889)
);

INVx11_ASAP7_75t_L g890 ( 
.A(n_602),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_646),
.A2(n_452),
.B(n_284),
.C(n_294),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_763),
.A2(n_428),
.B(n_452),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_670),
.B(n_428),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_L g894 ( 
.A(n_615),
.B(n_285),
.C(n_374),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_661),
.B(n_212),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_733),
.B(n_374),
.C(n_368),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_607),
.B(n_212),
.Y(n_897)
);

BUFx4f_ASAP7_75t_L g898 ( 
.A(n_616),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_731),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_629),
.A2(n_513),
.B(n_475),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_675),
.B(n_448),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_616),
.B(n_296),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_693),
.B(n_448),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_656),
.A2(n_448),
.B(n_445),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_625),
.A2(n_475),
.B(n_448),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_767),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_712),
.A2(n_475),
.B(n_445),
.Y(n_907)
);

CKINVDCx10_ASAP7_75t_R g908 ( 
.A(n_607),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_655),
.B(n_445),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_SL g910 ( 
.A(n_628),
.B(n_445),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_683),
.A2(n_446),
.B1(n_475),
.B2(n_99),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_734),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_650),
.B(n_446),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_764),
.B(n_446),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_751),
.B(n_475),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_714),
.A2(n_475),
.B(n_446),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_735),
.B(n_446),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_615),
.A2(n_446),
.B1(n_296),
.B2(n_257),
.Y(n_918)
);

OAI321xp33_ASAP7_75t_L g919 ( 
.A1(n_748),
.A2(n_296),
.A3(n_257),
.B1(n_446),
.B2(n_8),
.C(n_11),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_618),
.B(n_446),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_722),
.B(n_296),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_735),
.B(n_4),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_730),
.A2(n_152),
.B(n_143),
.Y(n_923)
);

AO21x1_ASAP7_75t_L g924 ( 
.A1(n_618),
.A2(n_6),
.B(n_7),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_616),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_721),
.B(n_6),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_694),
.A2(n_141),
.B(n_140),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_701),
.A2(n_129),
.B1(n_100),
.B2(n_98),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_752),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_695),
.B(n_15),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_616),
.Y(n_931)
);

O2A1O1Ixp5_ASAP7_75t_L g932 ( 
.A1(n_699),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_753),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_658),
.A2(n_16),
.B(n_18),
.C(n_21),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_715),
.A2(n_96),
.B1(n_93),
.B2(n_82),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_769),
.Y(n_936)
);

BUFx5_ASAP7_75t_L g937 ( 
.A(n_751),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_716),
.B(n_24),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_701),
.A2(n_80),
.B1(n_75),
.B2(n_69),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_703),
.B(n_67),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_708),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_749),
.A2(n_24),
.B(n_27),
.C(n_28),
.Y(n_942)
);

NOR2x1p5_ASAP7_75t_SL g943 ( 
.A(n_734),
.B(n_64),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_720),
.A2(n_28),
.B(n_31),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_758),
.A2(n_33),
.B(n_36),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_701),
.B(n_37),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_744),
.A2(n_746),
.B(n_759),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_716),
.B(n_38),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_716),
.B(n_38),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_724),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_766),
.A2(n_39),
.B(n_40),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_725),
.B(n_41),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_729),
.B(n_41),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_831),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_888),
.B(n_747),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_SL g956 ( 
.A(n_821),
.B(n_658),
.C(n_686),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_SL g957 ( 
.A(n_807),
.B(n_660),
.C(n_677),
.Y(n_957)
);

NOR2x1_ASAP7_75t_L g958 ( 
.A(n_802),
.B(n_842),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_773),
.B(n_691),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_931),
.B(n_770),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_833),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_777),
.A2(n_732),
.B(n_652),
.C(n_681),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_888),
.B(n_709),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_888),
.B(n_602),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_774),
.B(n_688),
.Y(n_965)
);

BUFx2_ASAP7_75t_L g966 ( 
.A(n_879),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_835),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_922),
.A2(n_716),
.B(n_747),
.C(n_738),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_788),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_774),
.B(n_713),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_875),
.A2(n_754),
.B(n_674),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_888),
.A2(n_738),
.B(n_755),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_860),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_804),
.B(n_704),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_822),
.B(n_672),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_938),
.B(n_602),
.C(n_755),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_822),
.B(n_757),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_947),
.A2(n_758),
.B(n_680),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_776),
.B(n_704),
.Y(n_979)
);

OAI21x1_ASAP7_75t_SL g980 ( 
.A1(n_924),
.A2(n_768),
.B(n_762),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_782),
.B(n_742),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_846),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_854),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_931),
.B(n_852),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_817),
.A2(n_765),
.B1(n_704),
.B2(n_750),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_869),
.A2(n_756),
.B(n_750),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_914),
.A2(n_775),
.B(n_826),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_816),
.A2(n_742),
.B(n_740),
.C(n_47),
.Y(n_989)
);

BUFx8_ASAP7_75t_L g990 ( 
.A(n_925),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_782),
.B(n_737),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_864),
.B(n_43),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_778),
.A2(n_43),
.B(n_44),
.C(n_47),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_784),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_785),
.A2(n_60),
.B(n_53),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_879),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_L g997 ( 
.A1(n_909),
.A2(n_52),
.B(n_55),
.C(n_56),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_SL g998 ( 
.A(n_919),
.B(n_57),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_783),
.A2(n_59),
.B(n_60),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_823),
.B(n_830),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_834),
.B(n_863),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_SL g1002 ( 
.A1(n_940),
.A2(n_920),
.B(n_946),
.C(n_921),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_834),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_863),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_843),
.B(n_950),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_898),
.B(n_842),
.Y(n_1006)
);

AO32x1_ASAP7_75t_L g1007 ( 
.A1(n_786),
.A2(n_935),
.A3(n_884),
.B1(n_805),
.B2(n_797),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_865),
.A2(n_942),
.B(n_827),
.C(n_949),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_902),
.Y(n_1009)
);

OAI22x1_ASAP7_75t_L g1010 ( 
.A1(n_950),
.A2(n_948),
.B1(n_949),
.B2(n_938),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_889),
.B(n_876),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_772),
.B(n_873),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_784),
.A2(n_928),
.B1(n_939),
.B2(n_898),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_870),
.A2(n_808),
.B(n_800),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_859),
.B(n_791),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_803),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_876),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_818),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_R g1019 ( 
.A(n_790),
.B(n_941),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_876),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_794),
.A2(n_812),
.B(n_862),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_920),
.A2(n_857),
.B(n_851),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_866),
.B(n_867),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_814),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_852),
.B(n_866),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_948),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_866),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_858),
.A2(n_953),
.B(n_952),
.C(n_894),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_876),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_910),
.A2(n_865),
.B1(n_895),
.B2(n_810),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_899),
.A2(n_933),
.B(n_929),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_818),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_906),
.B(n_802),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_936),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_894),
.A2(n_886),
.B(n_930),
.C(n_810),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_940),
.A2(n_825),
.B(n_871),
.C(n_917),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_787),
.A2(n_850),
.B1(n_906),
.B2(n_819),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_906),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_824),
.A2(n_848),
.B(n_880),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_913),
.A2(n_792),
.B(n_828),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_820),
.B(n_850),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_818),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_941),
.B(n_897),
.Y(n_1043)
);

NOR2x1p5_ASAP7_75t_SL g1044 ( 
.A(n_937),
.B(n_796),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_906),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_896),
.Y(n_1046)
);

AO21x1_ASAP7_75t_L g1047 ( 
.A1(n_911),
.A2(n_923),
.B(n_951),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_918),
.B(n_837),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_901),
.B(n_903),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_837),
.B(n_885),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_801),
.A2(n_943),
.B(n_781),
.C(n_793),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_878),
.B(n_882),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_904),
.A2(n_806),
.B1(n_944),
.B2(n_893),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_874),
.B(n_912),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_900),
.A2(n_779),
.B(n_780),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_789),
.B(n_934),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_811),
.B(n_861),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_813),
.A2(n_829),
.B(n_839),
.C(n_849),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_795),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_890),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_937),
.B(n_798),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_891),
.B(n_945),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_841),
.A2(n_845),
.B1(n_809),
.B2(n_815),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_937),
.B(n_892),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_937),
.A2(n_840),
.B1(n_892),
.B2(n_927),
.Y(n_1065)
);

BUFx8_ASAP7_75t_SL g1066 ( 
.A(n_908),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_799),
.B(n_840),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_937),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_847),
.A2(n_937),
.B1(n_836),
.B2(n_838),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_907),
.B(n_832),
.Y(n_1070)
);

CKINVDCx11_ASAP7_75t_R g1071 ( 
.A(n_932),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_853),
.A2(n_855),
.B(n_856),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_844),
.B(n_905),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_872),
.A2(n_883),
.B(n_877),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_881),
.A2(n_868),
.B(n_887),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_916),
.A2(n_915),
.B(n_932),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_915),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_773),
.B(n_509),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_773),
.B(n_931),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_784),
.A2(n_950),
.B1(n_821),
.B2(n_609),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_821),
.A2(n_669),
.B(n_777),
.C(n_662),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_773),
.B(n_509),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_773),
.B(n_609),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_821),
.B(n_509),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_788),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_773),
.B(n_609),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_824),
.A2(n_851),
.B(n_848),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_888),
.A2(n_622),
.B(n_623),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_773),
.B(n_609),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_875),
.A2(n_947),
.B(n_920),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_821),
.A2(n_669),
.B(n_777),
.C(n_662),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1075),
.A2(n_1021),
.B(n_1014),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1034),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1029),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_988),
.A2(n_970),
.B(n_977),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_L g1097 ( 
.A1(n_972),
.A2(n_1022),
.B(n_1076),
.Y(n_1097)
);

AO32x2_ASAP7_75t_L g1098 ( 
.A1(n_1080),
.A2(n_1013),
.A3(n_994),
.B1(n_1071),
.B2(n_1010),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1025),
.B(n_985),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1039),
.A2(n_978),
.B(n_987),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1004),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1082),
.B(n_1078),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1090),
.A2(n_971),
.B(n_1055),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_954),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_961),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1090),
.A2(n_971),
.B(n_1088),
.Y(n_1108)
);

BUFx12f_ASAP7_75t_L g1109 ( 
.A(n_1060),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_1008),
.C(n_1084),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_973),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_996),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1089),
.B(n_1050),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1089),
.B(n_959),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_1048),
.A2(n_1028),
.B(n_1035),
.C(n_962),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_983),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_967),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_992),
.A2(n_1080),
.B1(n_998),
.B2(n_994),
.C(n_1005),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_970),
.A2(n_1052),
.B(n_1040),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1025),
.B(n_985),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_984),
.Y(n_1121)
);

AOI221x1_ASAP7_75t_L g1122 ( 
.A1(n_1013),
.A2(n_995),
.B1(n_999),
.B2(n_1051),
.C(n_991),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1047),
.A2(n_1067),
.A3(n_1070),
.B(n_1058),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1079),
.B(n_1026),
.Y(n_1124)
);

AOI221x1_ASAP7_75t_L g1125 ( 
.A1(n_991),
.A2(n_975),
.B1(n_965),
.B2(n_980),
.C(n_1062),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1041),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1064),
.A2(n_1061),
.B(n_1073),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1049),
.A2(n_1041),
.B(n_965),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_974),
.A2(n_959),
.B1(n_979),
.B2(n_1079),
.Y(n_1129)
);

CKINVDCx14_ASAP7_75t_R g1130 ( 
.A(n_1060),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1026),
.B(n_1009),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1065),
.A2(n_968),
.B(n_1036),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_990),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1006),
.A2(n_993),
.B(n_1003),
.C(n_1043),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_981),
.A2(n_1061),
.A3(n_1045),
.B(n_1000),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_1030),
.A2(n_956),
.B(n_1031),
.C(n_957),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1069),
.A2(n_955),
.B(n_1000),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1012),
.B(n_1015),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1015),
.B(n_1059),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1054),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1057),
.B(n_1024),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_955),
.A2(n_1002),
.B(n_1054),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_SL g1143 ( 
.A1(n_963),
.A2(n_1023),
.B(n_1033),
.C(n_964),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1063),
.A2(n_1053),
.B(n_958),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_989),
.A2(n_1037),
.B(n_986),
.C(n_1046),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1066),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1068),
.A2(n_1007),
.B(n_1056),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_976),
.A2(n_997),
.B(n_1044),
.C(n_969),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1057),
.B(n_1085),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1032),
.B(n_1042),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1011),
.B(n_1038),
.Y(n_1151)
);

AND3x4_ASAP7_75t_L g1152 ( 
.A(n_960),
.B(n_1019),
.C(n_990),
.Y(n_1152)
);

AO21x1_ASAP7_75t_L g1153 ( 
.A1(n_1077),
.A2(n_1011),
.B(n_1007),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1057),
.B(n_1016),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_1029),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1056),
.A2(n_982),
.B(n_1077),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_960),
.A2(n_1057),
.B1(n_1018),
.B2(n_1001),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1056),
.A2(n_1029),
.B1(n_1038),
.B2(n_1020),
.Y(n_1158)
);

AO21x2_ASAP7_75t_L g1159 ( 
.A1(n_1017),
.A2(n_1038),
.B(n_1027),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1017),
.A2(n_1027),
.B(n_983),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_983),
.A2(n_1081),
.B(n_1091),
.C(n_821),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1162)
);

CKINVDCx6p67_ASAP7_75t_R g1163 ( 
.A(n_1004),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1047),
.A2(n_1051),
.A3(n_1067),
.B(n_1076),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1165)
);

AO21x1_ASAP7_75t_L g1166 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1048),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1034),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1047),
.A2(n_1051),
.A3(n_1067),
.B(n_1076),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1171)
);

BUFx4f_ASAP7_75t_L g1172 ( 
.A(n_1029),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_1091),
.B(n_1081),
.C(n_662),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_L g1177 ( 
.A(n_1081),
.B(n_1091),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_992),
.A2(n_662),
.B1(n_821),
.B2(n_817),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1047),
.A2(n_1051),
.A3(n_1067),
.B(n_1076),
.Y(n_1180)
);

BUFx10_ASAP7_75t_L g1181 ( 
.A(n_1043),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1083),
.B(n_509),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1047),
.A2(n_1051),
.A3(n_1067),
.B(n_1076),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1047),
.A2(n_1051),
.A3(n_1067),
.B(n_1076),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_992),
.A2(n_662),
.B1(n_821),
.B2(n_817),
.Y(n_1191)
);

AOI31xp67_ASAP7_75t_L g1192 ( 
.A1(n_1065),
.A2(n_1063),
.A3(n_1030),
.B(n_909),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1025),
.B(n_985),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1025),
.B(n_985),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1029),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1081),
.A2(n_1091),
.B1(n_1013),
.B2(n_1010),
.C(n_662),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1029),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1083),
.B(n_509),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_966),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_1083),
.B(n_506),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_L g1208 ( 
.A(n_1081),
.B(n_1091),
.C(n_662),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1048),
.A2(n_1091),
.B(n_1081),
.C(n_662),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1080),
.A2(n_1083),
.B1(n_1089),
.B2(n_1086),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_983),
.Y(n_1212)
);

CKINVDCx8_ASAP7_75t_R g1213 ( 
.A(n_966),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1214)
);

AO21x1_ASAP7_75t_L g1215 ( 
.A1(n_1013),
.A2(n_968),
.B(n_1048),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1081),
.A2(n_1091),
.B(n_821),
.C(n_1008),
.Y(n_1220)
);

BUFx4f_ASAP7_75t_L g1221 ( 
.A(n_1029),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1003),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1087),
.A2(n_1074),
.B(n_1072),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1029),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_988),
.A2(n_888),
.B(n_970),
.Y(n_1226)
);

NOR2x1_ASAP7_75t_L g1227 ( 
.A(n_1027),
.B(n_509),
.Y(n_1227)
);

INVx6_ASAP7_75t_L g1228 ( 
.A(n_1155),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1177),
.A2(n_1118),
.B1(n_1208),
.B2(n_1191),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1113),
.B(n_1105),
.Y(n_1230)
);

CKINVDCx8_ASAP7_75t_R g1231 ( 
.A(n_1146),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1208),
.A2(n_1184),
.B1(n_1202),
.B2(n_1181),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_1131),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1109),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1172),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1179),
.A2(n_1191),
.B1(n_1215),
.B2(n_1166),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1179),
.A2(n_1198),
.B1(n_1225),
.B2(n_1187),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1181),
.A2(n_1187),
.B1(n_1216),
.B2(n_1105),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1106),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1140),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1094),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1157),
.A2(n_1110),
.B1(n_1136),
.B2(n_1162),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1102),
.A2(n_1206),
.B1(n_1211),
.B2(n_1107),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1104),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1107),
.A2(n_1225),
.B1(n_1216),
.B2(n_1114),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1204),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1112),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1169),
.A2(n_1218),
.B1(n_1195),
.B2(n_1220),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1150),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1133),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1111),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1117),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1211),
.A2(n_1114),
.B1(n_1129),
.B2(n_1206),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1121),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1101),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1172),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1132),
.A2(n_1124),
.B1(n_1098),
.B2(n_1158),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1130),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1163),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1141),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1221),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1203),
.A2(n_1210),
.B1(n_1138),
.B2(n_1213),
.Y(n_1263)
);

INVx6_ASAP7_75t_L g1264 ( 
.A(n_1155),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1129),
.A2(n_1138),
.B1(n_1132),
.B2(n_1126),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1098),
.A2(n_1158),
.B1(n_1222),
.B2(n_1149),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1155),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1116),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1141),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1128),
.A2(n_1139),
.B1(n_1154),
.B2(n_1149),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1139),
.B(n_1175),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1221),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1099),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1227),
.A2(n_1115),
.B1(n_1196),
.B2(n_1099),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1116),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1119),
.A2(n_1144),
.B1(n_1096),
.B2(n_1098),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1209),
.A2(n_1152),
.B1(n_1194),
.B2(n_1196),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1127),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1120),
.B(n_1161),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1151),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_1147),
.B1(n_1137),
.B2(n_1153),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1212),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1224),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_SL g1284 ( 
.A1(n_1156),
.A2(n_1145),
.B1(n_1122),
.B2(n_1108),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1212),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1151),
.Y(n_1286)
);

INVx3_ASAP7_75t_SL g1287 ( 
.A(n_1095),
.Y(n_1287)
);

AOI22x1_ASAP7_75t_SL g1288 ( 
.A1(n_1197),
.A2(n_1201),
.B1(n_1134),
.B2(n_1143),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1125),
.A2(n_1226),
.B1(n_1214),
.B2(n_1182),
.Y(n_1289)
);

BUFx12f_ASAP7_75t_L g1290 ( 
.A(n_1201),
.Y(n_1290)
);

BUFx2_ASAP7_75t_SL g1291 ( 
.A(n_1165),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1167),
.A2(n_1207),
.B1(n_1205),
.B2(n_1200),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1148),
.A2(n_1174),
.B1(n_1188),
.B2(n_1173),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1160),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1183),
.A2(n_1185),
.B1(n_1193),
.B2(n_1199),
.Y(n_1295)
);

INVx3_ASAP7_75t_SL g1296 ( 
.A(n_1159),
.Y(n_1296)
);

INVx3_ASAP7_75t_SL g1297 ( 
.A(n_1159),
.Y(n_1297)
);

BUFx8_ASAP7_75t_SL g1298 ( 
.A(n_1097),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1142),
.A2(n_1100),
.B1(n_1192),
.B2(n_1123),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1123),
.A2(n_1092),
.B1(n_1223),
.B2(n_1219),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1171),
.B(n_1178),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1135),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1093),
.A2(n_1123),
.B1(n_1217),
.B2(n_1190),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1176),
.A2(n_1164),
.B1(n_1170),
.B2(n_1180),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1164),
.A2(n_1170),
.B1(n_1180),
.B2(n_1186),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1189),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1146),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1222),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1155),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1113),
.B(n_1184),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1168),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1112),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1155),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1179),
.A2(n_1191),
.B1(n_817),
.B2(n_620),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1208),
.A2(n_620),
.B1(n_817),
.B2(n_627),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1177),
.A2(n_1118),
.B1(n_1208),
.B2(n_950),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1113),
.B(n_1184),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1213),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1179),
.A2(n_1191),
.B1(n_817),
.B2(n_897),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1109),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1177),
.A2(n_1118),
.B1(n_1208),
.B2(n_950),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1213),
.Y(n_1322)
);

CKINVDCx6p67_ASAP7_75t_R g1323 ( 
.A(n_1109),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1168),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1112),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1168),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_SL g1327 ( 
.A1(n_1179),
.A2(n_620),
.B(n_627),
.Y(n_1327)
);

INVx6_ASAP7_75t_L g1328 ( 
.A(n_1155),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1109),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1204),
.Y(n_1330)
);

BUFx2_ASAP7_75t_SL g1331 ( 
.A(n_1213),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1168),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1109),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1168),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_SL g1335 ( 
.A(n_1109),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1278),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1246),
.B(n_1271),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1327),
.B(n_1310),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1317),
.B(n_1315),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1293),
.A2(n_1295),
.B(n_1301),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1250),
.B(n_1314),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1306),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1249),
.A2(n_1243),
.B1(n_1263),
.B2(n_1229),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1302),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1230),
.B(n_1238),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1296),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1297),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1301),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1292),
.A2(n_1300),
.B(n_1299),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1308),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1261),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1298),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1241),
.Y(n_1353)
);

INVxp33_ASAP7_75t_L g1354 ( 
.A(n_1330),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1319),
.A2(n_1229),
.B1(n_1316),
.B2(n_1321),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1269),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1316),
.A2(n_1321),
.B1(n_1237),
.B2(n_1232),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1242),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1237),
.B(n_1270),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1284),
.A2(n_1244),
.B(n_1265),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1245),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1253),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1255),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1270),
.B(n_1254),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1292),
.A2(n_1300),
.B(n_1299),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1254),
.B(n_1266),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1273),
.B(n_1312),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1258),
.B(n_1265),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1281),
.A2(n_1276),
.B(n_1304),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1298),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1281),
.A2(n_1276),
.B(n_1304),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1305),
.B(n_1240),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1294),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1234),
.A2(n_1280),
.B(n_1279),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1294),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1325),
.B(n_1248),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1291),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1311),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1324),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1326),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1332),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1239),
.B(n_1334),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1228),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1289),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1274),
.A2(n_1303),
.B(n_1277),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1288),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1228),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1282),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1282),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1252),
.A2(n_1287),
.B(n_1286),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1228),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1264),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1331),
.A2(n_1251),
.B1(n_1318),
.B2(n_1322),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1272),
.A2(n_1247),
.B(n_1262),
.C(n_1236),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1247),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1264),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1233),
.B(n_1285),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1313),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1343),
.A2(n_1260),
.B1(n_1251),
.B2(n_1259),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1354),
.B(n_1322),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1372),
.B(n_1233),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1343),
.A2(n_1260),
.B1(n_1272),
.B2(n_1256),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1384),
.A2(n_1333),
.B1(n_1329),
.B2(n_1236),
.C(n_1262),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_SL g1404 ( 
.A1(n_1394),
.A2(n_1328),
.B(n_1275),
.C(n_1309),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1337),
.A2(n_1360),
.B(n_1345),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1337),
.B(n_1256),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1355),
.A2(n_1262),
.B(n_1236),
.C(n_1257),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1345),
.B(n_1318),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1355),
.A2(n_1236),
.B(n_1257),
.C(n_1262),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1357),
.A2(n_1267),
.B(n_1309),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1384),
.A2(n_1329),
.B1(n_1333),
.B2(n_1257),
.C(n_1307),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1360),
.A2(n_1328),
.B(n_1323),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1358),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1338),
.A2(n_1339),
.B1(n_1386),
.B2(n_1366),
.Y(n_1414)
);

AOI211x1_ASAP7_75t_SL g1415 ( 
.A1(n_1382),
.A2(n_1275),
.B(n_1268),
.C(n_1290),
.Y(n_1415)
);

A2O1A1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1366),
.A2(n_1320),
.B(n_1283),
.C(n_1335),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_SL g1417 ( 
.A1(n_1386),
.A2(n_1320),
.B(n_1283),
.C(n_1335),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1342),
.B(n_1320),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1341),
.B(n_1231),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1344),
.B(n_1235),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1364),
.A2(n_1359),
.B(n_1368),
.C(n_1385),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1376),
.B(n_1367),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1395),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1374),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1388),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1350),
.B(n_1361),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1379),
.Y(n_1427)
);

BUFx2_ASAP7_75t_R g1428 ( 
.A(n_1370),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1395),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1362),
.B(n_1363),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1397),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1362),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1374),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1359),
.A2(n_1364),
.B(n_1382),
.C(n_1377),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1379),
.B(n_1380),
.Y(n_1435)
);

INVx8_ASAP7_75t_L g1436 ( 
.A(n_1396),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1349),
.A2(n_1365),
.B(n_1369),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1385),
.A2(n_1371),
.B(n_1369),
.C(n_1340),
.Y(n_1439)
);

NAND2xp33_ASAP7_75t_L g1440 ( 
.A(n_1352),
.B(n_1373),
.Y(n_1440)
);

AOI221x1_ASAP7_75t_L g1441 ( 
.A1(n_1377),
.A2(n_1352),
.B1(n_1391),
.B2(n_1398),
.C(n_1392),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1381),
.B(n_1356),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1353),
.B(n_1369),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1373),
.A2(n_1375),
.B(n_1352),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1351),
.B(n_1378),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1342),
.B(n_1374),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1385),
.A2(n_1371),
.B(n_1352),
.C(n_1375),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1443),
.B(n_1371),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1413),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.B(n_1349),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1413),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1446),
.B(n_1348),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1432),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1432),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1446),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1365),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1446),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1434),
.B(n_1414),
.C(n_1421),
.Y(n_1458)
);

NOR2x1p5_ASAP7_75t_L g1459 ( 
.A(n_1418),
.B(n_1373),
.Y(n_1459)
);

OAI222xp33_ASAP7_75t_L g1460 ( 
.A1(n_1402),
.A2(n_1370),
.B1(n_1375),
.B2(n_1373),
.C1(n_1389),
.C2(n_1388),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1427),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1445),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1435),
.B(n_1356),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1424),
.B(n_1433),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1347),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1423),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1426),
.B(n_1347),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1430),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1424),
.B(n_1348),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1442),
.B(n_1346),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1429),
.B(n_1346),
.Y(n_1471)
);

BUFx2_ASAP7_75t_SL g1472 ( 
.A(n_1418),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1439),
.B(n_1336),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1471),
.Y(n_1474)
);

OAI21xp33_ASAP7_75t_L g1475 ( 
.A1(n_1458),
.A2(n_1421),
.B(n_1399),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1465),
.B(n_1401),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1449),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1461),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1459),
.B(n_1440),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1461),
.Y(n_1480)
);

AOI31xp33_ASAP7_75t_L g1481 ( 
.A1(n_1458),
.A2(n_1418),
.A3(n_1412),
.B(n_1411),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1468),
.B(n_1447),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1466),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1464),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1452),
.B(n_1424),
.Y(n_1485)
);

OAI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1455),
.A2(n_1447),
.B1(n_1416),
.B2(n_1444),
.C(n_1406),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1465),
.B(n_1433),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1462),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.Y(n_1489)
);

OAI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1457),
.A2(n_1416),
.B1(n_1408),
.B2(n_1420),
.C(n_1419),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1463),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1456),
.B(n_1422),
.C(n_1407),
.D(n_1409),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1453),
.Y(n_1495)
);

OAI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1457),
.A2(n_1393),
.B1(n_1409),
.B2(n_1407),
.C(n_1403),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1452),
.B(n_1431),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1453),
.Y(n_1498)
);

AOI211xp5_ASAP7_75t_L g1499 ( 
.A1(n_1460),
.A2(n_1404),
.B(n_1410),
.C(n_1417),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1469),
.Y(n_1501)
);

OAI31xp33_ASAP7_75t_L g1502 ( 
.A1(n_1460),
.A2(n_1404),
.A3(n_1375),
.B(n_1417),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1456),
.B(n_1441),
.C(n_1440),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1454),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1487),
.B(n_1467),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1477),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1425),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1479),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1477),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1482),
.B(n_1450),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1485),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1488),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1484),
.B(n_1464),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_1478),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1482),
.B(n_1450),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1491),
.B(n_1462),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1484),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1480),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1492),
.Y(n_1519)
);

NOR3xp33_ASAP7_75t_L g1520 ( 
.A(n_1475),
.B(n_1400),
.C(n_1389),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1490),
.B(n_1425),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1500),
.B(n_1450),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1487),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1495),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1479),
.B(n_1459),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1503),
.B(n_1467),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1448),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1498),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1473),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1514),
.B(n_1483),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1519),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1528),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1528),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1519),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1524),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1518),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1524),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1528),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1513),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1508),
.B(n_1530),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1518),
.B(n_1483),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1528),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1530),
.B(n_1501),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1506),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1530),
.B(n_1485),
.Y(n_1549)
);

NAND2x1_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1522),
.B(n_1485),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1522),
.B(n_1485),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1504),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1512),
.B(n_1526),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1526),
.B(n_1504),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1520),
.A2(n_1499),
.B1(n_1481),
.B2(n_1496),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1520),
.A2(n_1481),
.B1(n_1405),
.B2(n_1494),
.C(n_1503),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1522),
.B(n_1493),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1506),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1526),
.B(n_1489),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1523),
.B(n_1476),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1509),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1509),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1474),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1525),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1513),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1511),
.B(n_1513),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1505),
.B(n_1474),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1511),
.B(n_1493),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1550),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1556),
.B(n_1507),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1510),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1547),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1547),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1556),
.B(n_1507),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1557),
.B(n_1502),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1557),
.A2(n_1499),
.B1(n_1521),
.B2(n_1486),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1510),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1531),
.B(n_1521),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1550),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1543),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1548),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1531),
.B(n_1510),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1544),
.B(n_1428),
.Y(n_1587)
);

NAND2x1p5_ASAP7_75t_L g1588 ( 
.A(n_1566),
.B(n_1390),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1548),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1544),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1533),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1561),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1554),
.A2(n_1502),
.B(n_1494),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1560),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1561),
.B(n_1523),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1560),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1511),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1523),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1566),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1549),
.B(n_1511),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1546),
.A2(n_1472),
.B1(n_1497),
.B2(n_1342),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1546),
.B(n_1516),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1505),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1575),
.B(n_1549),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1574),
.B(n_1562),
.Y(n_1609)
);

AOI32xp33_ASAP7_75t_L g1610 ( 
.A1(n_1580),
.A2(n_1546),
.A3(n_1540),
.B1(n_1541),
.B2(n_1551),
.Y(n_1610)
);

NAND4xp75_ASAP7_75t_SL g1611 ( 
.A(n_1587),
.B(n_1540),
.C(n_1541),
.D(n_1569),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1583),
.B(n_1472),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1593),
.B(n_1555),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1576),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1578),
.A2(n_1555),
.B(n_1553),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1582),
.B(n_1562),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1573),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1603),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1583),
.A2(n_1562),
.B1(n_1541),
.B2(n_1540),
.C(n_1565),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1592),
.B(n_1516),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1577),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1592),
.B(n_1535),
.C(n_1532),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1573),
.A2(n_1552),
.B1(n_1571),
.B2(n_1569),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1577),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1585),
.Y(n_1629)
);

NAND3x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1601),
.C(n_1607),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1585),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1586),
.A2(n_1568),
.B1(n_1572),
.B2(n_1569),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1613),
.B(n_1584),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1621),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1614),
.A2(n_1573),
.B1(n_1598),
.B2(n_1584),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1608),
.B(n_1597),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1610),
.A2(n_1615),
.B(n_1617),
.C(n_1609),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_R g1639 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1620),
.A2(n_1603),
.B1(n_1619),
.B2(n_1623),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1630),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1608),
.B(n_1597),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1575),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1581),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1622),
.A2(n_1588),
.B(n_1596),
.C(n_1535),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1618),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1632),
.B(n_1581),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1626),
.A2(n_1536),
.B1(n_1538),
.B2(n_1532),
.C1(n_1604),
.C2(n_1589),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1618),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1616),
.B(n_1629),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1624),
.Y(n_1651)
);

AOI322xp5_ASAP7_75t_L g1652 ( 
.A1(n_1641),
.A2(n_1611),
.A3(n_1631),
.B1(n_1624),
.B2(n_1628),
.C1(n_1536),
.C2(n_1538),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1641),
.A2(n_1588),
.B1(n_1601),
.B2(n_1602),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1640),
.B(n_1628),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_SL g1655 ( 
.A(n_1645),
.B(n_1588),
.C(n_1605),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1639),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1637),
.A2(n_1604),
.B(n_1607),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1636),
.Y(n_1658)
);

AOI211xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1640),
.A2(n_1602),
.B(n_1600),
.C(n_1589),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_SL g1660 ( 
.A1(n_1634),
.A2(n_1602),
.B(n_1591),
.C(n_1594),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1646),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1649),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1643),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1658),
.B(n_1635),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1654),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1656),
.B(n_1637),
.Y(n_1666)
);

NAND5xp2_ASAP7_75t_L g1667 ( 
.A(n_1659),
.B(n_1648),
.C(n_1647),
.D(n_1633),
.E(n_1644),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1659),
.A2(n_1638),
.B1(n_1650),
.B2(n_1651),
.C(n_1642),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1655),
.A2(n_1600),
.B1(n_1602),
.B2(n_1599),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1661),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1663),
.B(n_1599),
.C(n_1594),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1662),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1652),
.B(n_1657),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1665),
.A2(n_1653),
.B1(n_1600),
.B2(n_1568),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1667),
.B(n_1660),
.C(n_1600),
.D(n_1591),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_L g1676 ( 
.A(n_1666),
.B(n_1567),
.C(n_1542),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1673),
.A2(n_1542),
.B1(n_1567),
.B2(n_1564),
.C(n_1563),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1563),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1675),
.A2(n_1669),
.B(n_1668),
.C(n_1671),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1678),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1674),
.A2(n_1664),
.B1(n_1670),
.B2(n_1672),
.Y(n_1681)
);

OAI211xp5_ASAP7_75t_L g1682 ( 
.A1(n_1677),
.A2(n_1567),
.B(n_1542),
.C(n_1565),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1676),
.B(n_1534),
.C(n_1533),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1675),
.B(n_1551),
.Y(n_1684)
);

NAND4xp75_ASAP7_75t_L g1685 ( 
.A(n_1680),
.B(n_1553),
.C(n_1564),
.D(n_1571),
.Y(n_1685)
);

NAND4xp75_ASAP7_75t_L g1686 ( 
.A(n_1684),
.B(n_1571),
.C(n_1551),
.D(n_1559),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1681),
.Y(n_1687)
);

NOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1679),
.B(n_1542),
.Y(n_1688)
);

NOR2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1683),
.B(n_1567),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1687),
.B(n_1682),
.C(n_1534),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1686),
.A2(n_1568),
.B1(n_1511),
.B2(n_1517),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1688),
.A2(n_1568),
.B1(n_1572),
.B2(n_1559),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1690),
.Y(n_1693)
);

OAI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1689),
.B1(n_1692),
.B2(n_1685),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1694),
.A2(n_1691),
.B1(n_1572),
.B2(n_1517),
.Y(n_1695)
);

AOI22x1_ASAP7_75t_L g1696 ( 
.A1(n_1694),
.A2(n_1534),
.B1(n_1533),
.B2(n_1558),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1539),
.Y(n_1697)
);

OAI22x1_ASAP7_75t_L g1698 ( 
.A1(n_1696),
.A2(n_1572),
.B1(n_1539),
.B2(n_1558),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1697),
.A2(n_1558),
.B1(n_1545),
.B2(n_1539),
.C(n_1517),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1698),
.A2(n_1572),
.B1(n_1545),
.B2(n_1390),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1700),
.B(n_1545),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1699),
.B(n_1383),
.C(n_1387),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

OAI221xp5_ASAP7_75t_R g1704 ( 
.A1(n_1703),
.A2(n_1436),
.B1(n_1552),
.B2(n_1559),
.C(n_1415),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1704),
.A2(n_1383),
.B(n_1387),
.C(n_1396),
.Y(n_1705)
);


endmodule