module fake_netlist_6_2992_n_548 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_548);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_548;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_525;
wire n_156;
wire n_491;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_456;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_477;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_546;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_16),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_31),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_21),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_33),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_99),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_43),
.B(n_121),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_72),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_108),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_50),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_39),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_73),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_103),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_26),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_41),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_112),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_70),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_65),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_143),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_55),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_32),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_69),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_88),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_6),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_46),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_111),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_67),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_78),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_77),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_76),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_101),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_107),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_94),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_44),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_47),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_58),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_141),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_85),
.B(n_59),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_126),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_28),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_0),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_0),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

BUFx8_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_159),
.Y(n_252)
);

CKINVDCx6p67_ASAP7_75t_R g253 ( 
.A(n_172),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_174),
.A2(n_71),
.B(n_154),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_1),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_215),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_2),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_161),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_164),
.Y(n_263)
);

AND2x6_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_167),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_165),
.B(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_169),
.Y(n_266)
);

CKINVDCx6p67_ASAP7_75t_R g267 ( 
.A(n_158),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_177),
.B(n_178),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_186),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_188),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_190),
.B(n_5),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_266),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_267),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_245),
.Y(n_288)
);

BUFx6f_ASAP7_75t_SL g289 ( 
.A(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_162),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_207),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_204),
.B1(n_198),
.B2(n_217),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_192),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_257),
.B(n_199),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_207),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_266),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_217),
.B1(n_237),
.B2(n_224),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_262),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_250),
.B(n_196),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_276),
.B(n_208),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_197),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_255),
.A2(n_224),
.B1(n_237),
.B2(n_210),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_255),
.A2(n_238),
.B1(n_202),
.B2(n_233),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_219),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_265),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_295),
.A2(n_258),
.B1(n_249),
.B2(n_250),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_247),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_291),
.B(n_247),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_249),
.B1(n_211),
.B2(n_203),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_304),
.A2(n_269),
.B1(n_264),
.B2(n_274),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_271),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_307),
.A2(n_272),
.B(n_274),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_285),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_272),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_284),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_286),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_269),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_303),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_269),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_269),
.Y(n_339)
);

OAI221xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_263),
.B1(n_273),
.B2(n_206),
.C(n_212),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_264),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_264),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_283),
.B(n_160),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_283),
.B(n_168),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_280),
.B(n_264),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_280),
.B(n_263),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_279),
.B(n_171),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_318),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_296),
.A2(n_214),
.B1(n_175),
.B2(n_176),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_316),
.Y(n_353)
);

INVx5_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_273),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_313),
.B1(n_312),
.B2(n_309),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_305),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_305),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_270),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_298),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_270),
.Y(n_363)
);

O2A1O1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_319),
.A2(n_312),
.B(n_313),
.C(n_315),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_356),
.A2(n_289),
.B1(n_213),
.B2(n_220),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_335),
.A2(n_309),
.B1(n_170),
.B2(n_223),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_321),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_341),
.B(n_342),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_327),
.B(n_282),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_329),
.A2(n_311),
.B(n_306),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_340),
.B1(n_352),
.B2(n_359),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_256),
.B(n_209),
.C(n_226),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_R g373 ( 
.A(n_328),
.B(n_331),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_333),
.A2(n_221),
.B(n_230),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_SL g377 ( 
.A(n_363),
.B(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_361),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_346),
.B(n_181),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_336),
.A2(n_232),
.B(n_182),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_317),
.B(n_296),
.C(n_309),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_339),
.A2(n_205),
.B(n_185),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_362),
.Y(n_384)
);

O2A1O1Ixp33_ASAP7_75t_L g385 ( 
.A1(n_355),
.A2(n_317),
.B(n_309),
.C(n_277),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_277),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_363),
.B1(n_330),
.B2(n_348),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_353),
.B(n_351),
.Y(n_389)
);

AOI22x1_ASAP7_75t_L g390 ( 
.A1(n_348),
.A2(n_236),
.B1(n_225),
.B2(n_222),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_343),
.B(n_183),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_193),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_349),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_324),
.A2(n_218),
.B(n_201),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_334),
.A2(n_200),
.B(n_80),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_338),
.B(n_9),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_SL g397 ( 
.A1(n_320),
.A2(n_79),
.B(n_152),
.C(n_150),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_5),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_332),
.B(n_7),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_323),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_337),
.B(n_75),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_320),
.A2(n_82),
.B1(n_148),
.B2(n_13),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_337),
.B(n_7),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_375),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_8),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_354),
.Y(n_407)
);

AO21x2_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_354),
.B(n_15),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_354),
.B(n_8),
.C(n_18),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_382),
.Y(n_410)
);

OAI21x1_ASAP7_75t_SL g411 ( 
.A1(n_396),
.A2(n_17),
.B(n_19),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

AO31x2_ASAP7_75t_L g413 ( 
.A1(n_372),
.A2(n_20),
.A3(n_22),
.B(n_23),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_374),
.A2(n_24),
.B(n_27),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_30),
.Y(n_415)
);

AOI221x1_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C(n_42),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_45),
.B(n_48),
.C(n_49),
.Y(n_417)
);

O2A1O1Ixp33_ASAP7_75t_SL g418 ( 
.A1(n_397),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_385),
.A2(n_56),
.B(n_57),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_379),
.A2(n_60),
.B(n_61),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_62),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

AO21x2_ASAP7_75t_L g424 ( 
.A1(n_373),
.A2(n_64),
.B(n_66),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g426 ( 
.A1(n_366),
.A2(n_83),
.B(n_84),
.Y(n_426)
);

AOI221xp5_ASAP7_75t_SL g427 ( 
.A1(n_388),
.A2(n_86),
.B1(n_87),
.B2(n_93),
.C(n_95),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_389),
.A2(n_97),
.B(n_100),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_370),
.A2(n_395),
.B(n_380),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_369),
.B(n_102),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_392),
.B(n_109),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_398),
.A2(n_117),
.B1(n_118),
.B2(n_122),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_123),
.Y(n_434)
);

AO22x2_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_124),
.B1(n_125),
.B2(n_128),
.Y(n_435)
);

AO21x2_ASAP7_75t_L g436 ( 
.A1(n_407),
.A2(n_408),
.B(n_419),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_412),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_403),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_431),
.A2(n_394),
.B1(n_367),
.B2(n_383),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_427),
.A2(n_390),
.B(n_377),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_367),
.B1(n_404),
.B2(n_400),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_131),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_415),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_133),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_406),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_134),
.Y(n_447)
);

AO31x2_ASAP7_75t_L g448 ( 
.A1(n_409),
.A2(n_137),
.A3(n_144),
.B(n_146),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_422),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_428),
.A2(n_429),
.B(n_411),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_423),
.B(n_430),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_437),
.Y(n_458)
);

AO21x2_ASAP7_75t_L g459 ( 
.A1(n_452),
.A2(n_408),
.B(n_417),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_454),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_451),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_442),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_435),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_452),
.A2(n_418),
.B(n_424),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_413),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_461),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_469),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_439),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_445),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_439),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_444),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_444),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_473),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_421),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_467),
.B(n_421),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_449),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_449),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_453),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_463),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_458),
.Y(n_492)
);

INVx2_ASAP7_75t_SL g493 ( 
.A(n_468),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_472),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_490),
.B(n_472),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_449),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_479),
.B(n_453),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_448),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_482),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_455),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_492),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_488),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_491),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_448),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_482),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_447),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_486),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_510),
.B(n_478),
.Y(n_512)
);

AOI32xp33_ASAP7_75t_L g513 ( 
.A1(n_499),
.A2(n_485),
.A3(n_432),
.B1(n_433),
.B2(n_483),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_481),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_500),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_487),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_503),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_493),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_501),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_518),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_515),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_495),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_512),
.C(n_513),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_514),
.Y(n_525)
);

OAI321xp33_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_524),
.A3(n_513),
.B1(n_525),
.B2(n_516),
.C(n_497),
.Y(n_526)
);

AOI221xp5_ASAP7_75t_L g527 ( 
.A1(n_523),
.A2(n_519),
.B1(n_507),
.B2(n_505),
.C(n_496),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_525),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_528),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_L g530 ( 
.A1(n_527),
.A2(n_495),
.B(n_440),
.Y(n_530)
);

OAI211xp5_ASAP7_75t_SL g531 ( 
.A1(n_526),
.A2(n_420),
.B(n_504),
.C(n_443),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_SL g532 ( 
.A(n_529),
.B(n_509),
.C(n_502),
.Y(n_532)
);

OAI311xp33_ASAP7_75t_L g533 ( 
.A1(n_530),
.A2(n_502),
.A3(n_457),
.B1(n_416),
.C1(n_496),
.Y(n_533)
);

NAND4xp75_ASAP7_75t_L g534 ( 
.A(n_531),
.B(n_493),
.C(n_441),
.D(n_414),
.Y(n_534)
);

NAND2x1p5_ASAP7_75t_L g535 ( 
.A(n_532),
.B(n_509),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_424),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_535),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_536),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_482),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_539),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_539),
.A2(n_537),
.B1(n_533),
.B2(n_457),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_540),
.A2(n_426),
.B(n_441),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_147),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_543),
.A2(n_441),
.B(n_436),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_542),
.A2(n_448),
.B1(n_413),
.B2(n_471),
.Y(n_545)
);

AOI21xp33_ASAP7_75t_L g546 ( 
.A1(n_544),
.A2(n_155),
.B(n_436),
.Y(n_546)
);

AO221x2_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_545),
.B1(n_448),
.B2(n_471),
.C(n_459),
.Y(n_547)
);

AOI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_547),
.A2(n_471),
.B(n_459),
.Y(n_548)
);


endmodule