module real_aes_8319_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_335;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g182 ( .A1(n_0), .A2(n_183), .B(n_184), .C(n_188), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_1), .B(n_178), .Y(n_189) );
INVx1_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_3), .B(n_143), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_4), .A2(n_124), .B(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_5), .A2(n_129), .B(n_134), .C(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_6), .A2(n_124), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_7), .B(n_178), .Y(n_478) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_8), .A2(n_157), .B(n_207), .Y(n_206) );
AND2x6_ASAP7_75t_L g129 ( .A(n_9), .B(n_130), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_10), .A2(n_129), .B(n_134), .C(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g533 ( .A(n_11), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_12), .B(n_41), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_12), .B(n_41), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_13), .B(n_187), .Y(n_510) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_15), .A2(n_100), .B1(n_108), .B2(n_740), .Y(n_99) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_16), .B(n_143), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_17), .A2(n_144), .B(n_518), .C(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_18), .B(n_178), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_19), .B(n_171), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_20), .A2(n_134), .B(n_165), .C(n_170), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_21), .A2(n_186), .B(n_201), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_22), .B(n_187), .Y(n_463) );
OAI222xp33_ASAP7_75t_L g443 ( .A1(n_23), .A2(n_444), .B1(n_726), .B2(n_727), .C1(n_733), .C2(n_737), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_23), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_24), .B(n_187), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_25), .Y(n_459) );
INVx1_ASAP7_75t_L g484 ( .A(n_26), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_27), .A2(n_134), .B(n_170), .C(n_210), .Y(n_209) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_29), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_30), .Y(n_737) );
INVx1_ASAP7_75t_L g560 ( .A(n_31), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_32), .A2(n_124), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g127 ( .A(n_33), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_34), .A2(n_132), .B(n_137), .C(n_147), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_35), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_36), .A2(n_186), .B(n_475), .C(n_477), .Y(n_474) );
INVxp67_ASAP7_75t_L g561 ( .A(n_37), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_38), .B(n_212), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_39), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_40), .A2(n_134), .B(n_170), .C(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_42), .A2(n_188), .B(n_531), .C(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_43), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_44), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_45), .B(n_143), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_46), .B(n_124), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_47), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_48), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_49), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_50), .A2(n_132), .B(n_147), .C(n_221), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_51), .A2(n_115), .B1(n_116), .B2(n_434), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_51), .Y(n_115) );
INVx1_ASAP7_75t_L g185 ( .A(n_52), .Y(n_185) );
INVx1_ASAP7_75t_L g222 ( .A(n_53), .Y(n_222) );
INVx1_ASAP7_75t_L g496 ( .A(n_54), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_55), .B(n_124), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_56), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_57), .Y(n_529) );
INVx1_ASAP7_75t_L g130 ( .A(n_58), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_59), .B(n_124), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_60), .B(n_178), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_61), .A2(n_169), .B(n_232), .C(n_234), .Y(n_231) );
INVx1_ASAP7_75t_L g152 ( .A(n_62), .Y(n_152) );
INVx1_ASAP7_75t_SL g476 ( .A(n_63), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_64), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_65), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_66), .B(n_178), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_67), .B(n_144), .Y(n_198) );
INVx1_ASAP7_75t_L g462 ( .A(n_68), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_69), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_70), .B(n_140), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_71), .A2(n_134), .B(n_147), .C(n_258), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_72), .Y(n_230) );
INVx1_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_74), .A2(n_124), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_75), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_76), .A2(n_124), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_77), .A2(n_163), .B(n_556), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_78), .Y(n_481) );
INVx1_ASAP7_75t_L g516 ( .A(n_79), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_80), .B(n_139), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_81), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_82), .A2(n_124), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g519 ( .A(n_83), .Y(n_519) );
INVx2_ASAP7_75t_L g150 ( .A(n_84), .Y(n_150) );
INVx1_ASAP7_75t_L g509 ( .A(n_85), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_86), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_87), .B(n_187), .Y(n_199) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_88), .B(n_104), .C(n_105), .Y(n_103) );
OR2x2_ASAP7_75t_L g436 ( .A(n_88), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g446 ( .A(n_88), .B(n_438), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_88), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_89), .A2(n_134), .B(n_147), .C(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_90), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVxp67_ASAP7_75t_L g235 ( .A(n_92), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_93), .B(n_157), .Y(n_534) );
INVx2_ASAP7_75t_L g499 ( .A(n_94), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_95), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g194 ( .A(n_96), .Y(n_194) );
INVx1_ASAP7_75t_L g259 ( .A(n_97), .Y(n_259) );
AND2x2_ASAP7_75t_L g224 ( .A(n_98), .B(n_149), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_100), .Y(n_740) );
CKINVDCx12_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
AND2x2_ASAP7_75t_L g438 ( .A(n_104), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI21x1_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_113), .B(n_442), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g739 ( .A(n_111), .Y(n_739) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_435), .B(n_440), .Y(n_113) );
INVx2_ASAP7_75t_L g434 ( .A(n_116), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_116), .A2(n_728), .B1(n_731), .B2(n_732), .Y(n_727) );
OR3x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_348), .C(n_391), .Y(n_116) );
NAND5xp2_ASAP7_75t_L g117 ( .A(n_118), .B(n_275), .C(n_305), .D(n_322), .E(n_337), .Y(n_117) );
AOI221xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_190), .B1(n_237), .B2(n_243), .C(n_247), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_159), .Y(n_119) );
OR2x2_ASAP7_75t_L g252 ( .A(n_120), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g292 ( .A(n_120), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_120), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_120), .B(n_245), .Y(n_327) );
OR2x2_ASAP7_75t_L g339 ( .A(n_120), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_120), .B(n_298), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_120), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_120), .B(n_276), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_120), .B(n_284), .Y(n_390) );
AND2x2_ASAP7_75t_L g422 ( .A(n_120), .B(n_176), .Y(n_422) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_120), .Y(n_430) );
INVx5_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_121), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g249 ( .A(n_121), .B(n_225), .Y(n_249) );
BUFx2_ASAP7_75t_L g272 ( .A(n_121), .Y(n_272) );
AND2x2_ASAP7_75t_L g301 ( .A(n_121), .B(n_160), .Y(n_301) );
AND2x2_ASAP7_75t_L g356 ( .A(n_121), .B(n_253), .Y(n_356) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_154), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_131), .B(n_149), .Y(n_122) );
BUFx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_125), .B(n_129), .Y(n_195) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
INVx1_ASAP7_75t_L g202 ( .A(n_127), .Y(n_202) );
INVx1_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_128), .Y(n_141) );
INVx3_ASAP7_75t_L g144 ( .A(n_128), .Y(n_144) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_128), .Y(n_187) );
INVx1_ASAP7_75t_L g212 ( .A(n_128), .Y(n_212) );
INVx4_ASAP7_75t_SL g148 ( .A(n_129), .Y(n_148) );
BUFx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_SL g180 ( .A1(n_133), .A2(n_148), .B(n_181), .C(n_182), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_133), .A2(n_148), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_133), .A2(n_148), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_133), .A2(n_148), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_133), .A2(n_148), .B(n_516), .C(n_517), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_133), .A2(n_148), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g556 ( .A1(n_133), .A2(n_148), .B(n_557), .C(n_558), .Y(n_556) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx3_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_135), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_142), .C(n_145), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_139), .A2(n_145), .B(n_222), .C(n_223), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_139), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
O2A1O1Ixp5_ASAP7_75t_L g508 ( .A1(n_139), .A2(n_464), .B(n_509), .C(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g233 ( .A(n_141), .Y(n_233) );
INVx2_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_143), .B(n_235), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_143), .A2(n_168), .B(n_484), .C(n_485), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_143), .A2(n_233), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_144), .B(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
INVx1_ASAP7_75t_L g520 ( .A(n_146), .Y(n_520) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx1_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_149), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_149), .A2(n_195), .B(n_481), .C(n_482), .Y(n_480) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_149), .A2(n_527), .B(n_534), .Y(n_526) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g158 ( .A(n_150), .B(n_151), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx3_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_156), .A2(n_193), .B(n_203), .Y(n_192) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_156), .A2(n_256), .B(n_264), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_156), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_156), .A2(n_458), .B(n_465), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_156), .B(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_156), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_157), .A2(n_208), .B(n_209), .Y(n_207) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_157), .Y(n_227) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_159), .B(n_310), .Y(n_319) );
OAI32xp33_ASAP7_75t_L g333 ( .A1(n_159), .A2(n_269), .A3(n_334), .B1(n_335), .B2(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_159), .B(n_335), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_159), .B(n_252), .Y(n_376) );
INVx1_ASAP7_75t_SL g405 ( .A(n_159), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_159), .B(n_192), .C(n_356), .D(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
INVx5_ASAP7_75t_L g246 ( .A(n_160), .Y(n_246) );
AND2x2_ASAP7_75t_L g276 ( .A(n_160), .B(n_177), .Y(n_276) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_160), .Y(n_355) );
AND2x2_ASAP7_75t_L g425 ( .A(n_160), .B(n_372), .Y(n_425) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_173), .Y(n_160) );
AOI21xp5_ASAP7_75t_SL g161 ( .A1(n_162), .A2(n_164), .B(n_171), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .Y(n_165) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_169), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_172), .B(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_175), .A2(n_505), .B(n_511), .Y(n_504) );
AND2x4_ASAP7_75t_L g298 ( .A(n_176), .B(n_246), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_176), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g332 ( .A(n_176), .B(n_253), .Y(n_332) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g245 ( .A(n_177), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g284 ( .A(n_177), .B(n_255), .Y(n_284) );
AND2x2_ASAP7_75t_L g293 ( .A(n_177), .B(n_254), .Y(n_293) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_189), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_186), .B(n_476), .Y(n_475) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g531 ( .A(n_187), .Y(n_531) );
INVx2_ASAP7_75t_L g464 ( .A(n_188), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_190), .A2(n_362), .B1(n_364), .B2(n_366), .C1(n_369), .C2(n_370), .Y(n_361) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_214), .Y(n_190) );
AND2x2_ASAP7_75t_L g294 ( .A(n_191), .B(n_295), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_191), .B(n_272), .C(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_206), .Y(n_191) );
INVx5_ASAP7_75t_SL g242 ( .A(n_192), .Y(n_242) );
OAI322xp33_ASAP7_75t_L g247 ( .A1(n_192), .A2(n_248), .A3(n_250), .B1(n_251), .B2(n_266), .C1(n_269), .C2(n_271), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_192), .B(n_240), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_192), .B(n_226), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_195), .A2(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_195), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_200), .A2(n_211), .B(n_213), .Y(n_210) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
INVx2_ASAP7_75t_L g554 ( .A(n_205), .Y(n_554) );
INVx2_ASAP7_75t_L g240 ( .A(n_206), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_206), .B(n_216), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_214), .B(n_279), .Y(n_334) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR2x2_ASAP7_75t_L g313 ( .A(n_215), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_225), .Y(n_215) );
OR2x2_ASAP7_75t_L g241 ( .A(n_216), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_216), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g281 ( .A(n_216), .B(n_226), .Y(n_281) );
AND2x2_ASAP7_75t_L g304 ( .A(n_216), .B(n_240), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_216), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_216), .B(n_279), .Y(n_320) );
AND2x2_ASAP7_75t_L g328 ( .A(n_216), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_216), .B(n_288), .Y(n_378) );
INVx5_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g268 ( .A(n_217), .B(n_242), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_217), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_217), .B(n_226), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_217), .B(n_342), .Y(n_383) );
OR2x2_ASAP7_75t_L g399 ( .A(n_217), .B(n_343), .Y(n_399) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_217), .B(n_360), .Y(n_406) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_217), .Y(n_413) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
AND2x2_ASAP7_75t_L g267 ( .A(n_225), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g317 ( .A(n_225), .B(n_240), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_225), .B(n_242), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_225), .B(n_279), .Y(n_401) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_226), .B(n_242), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_226), .B(n_240), .Y(n_289) );
OR2x2_ASAP7_75t_L g343 ( .A(n_226), .B(n_240), .Y(n_343) );
AND2x2_ASAP7_75t_L g360 ( .A(n_226), .B(n_239), .Y(n_360) );
INVxp67_ASAP7_75t_L g382 ( .A(n_226), .Y(n_382) );
AND2x2_ASAP7_75t_L g409 ( .A(n_226), .B(n_279), .Y(n_409) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_226), .Y(n_416) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_236), .Y(n_226) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_227), .A2(n_471), .B(n_478), .Y(n_470) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_227), .A2(n_494), .B(n_500), .Y(n_493) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_227), .A2(n_514), .B(n_521), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_259), .B(n_260), .C(n_261), .Y(n_258) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_233), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_233), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_239), .B(n_290), .Y(n_363) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g279 ( .A(n_240), .B(n_242), .Y(n_279) );
OR2x2_ASAP7_75t_L g346 ( .A(n_240), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g290 ( .A(n_241), .Y(n_290) );
OR2x2_ASAP7_75t_L g351 ( .A(n_241), .B(n_343), .Y(n_351) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g250 ( .A(n_245), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_245), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g251 ( .A(n_246), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_246), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_246), .B(n_253), .Y(n_286) );
INVx2_ASAP7_75t_L g331 ( .A(n_246), .Y(n_331) );
AND2x2_ASAP7_75t_L g344 ( .A(n_246), .B(n_284), .Y(n_344) );
AND2x2_ASAP7_75t_L g369 ( .A(n_246), .B(n_293), .Y(n_369) );
INVx1_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
INVx2_ASAP7_75t_SL g308 ( .A(n_252), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_253), .Y(n_311) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx2_ASAP7_75t_L g372 ( .A(n_255), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_263), .Y(n_256) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx3_ASAP7_75t_L g477 ( .A(n_262), .Y(n_477) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g341 ( .A(n_268), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_268), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_268), .A2(n_350), .B1(n_352), .B2(n_357), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_268), .B(n_360), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_269), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g303 ( .A(n_270), .Y(n_303) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OR2x2_ASAP7_75t_L g285 ( .A(n_272), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_272), .B(n_276), .Y(n_336) );
AND2x2_ASAP7_75t_L g359 ( .A(n_272), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g335 ( .A(n_274), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_277), .B(n_282), .C(n_296), .Y(n_275) );
INVx1_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_276), .A2(n_408), .B1(n_410), .B2(n_411), .C(n_414), .Y(n_407) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g426 ( .A(n_279), .Y(n_426) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g375 ( .A(n_281), .B(n_314), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B(n_287), .C(n_291), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OAI32xp33_ASAP7_75t_L g400 ( .A1(n_289), .A2(n_290), .A3(n_353), .B1(n_390), .B2(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
AND2x2_ASAP7_75t_L g432 ( .A(n_292), .B(n_331), .Y(n_432) );
AND2x2_ASAP7_75t_L g379 ( .A(n_293), .B(n_331), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_293), .B(n_301), .Y(n_397) );
AOI31xp33_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_299), .A3(n_300), .B(n_302), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_298), .B(n_310), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_298), .B(n_308), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_298), .A2(n_328), .B1(n_418), .B2(n_421), .C(n_423), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x2_ASAP7_75t_L g323 ( .A(n_303), .B(n_324), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_315), .B2(n_318), .C1(n_320), .C2(n_321), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g388 ( .A(n_307), .Y(n_388) );
INVx1_ASAP7_75t_L g410 ( .A(n_310), .Y(n_410) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_313), .A2(n_424), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx1_ASAP7_75t_L g329 ( .A(n_314), .Y(n_329) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_326), .B1(n_328), .B2(n_330), .C(n_333), .Y(n_322) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g367 ( .A(n_325), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g419 ( .A(n_325), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g394 ( .A(n_330), .Y(n_394) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
INVx1_ASAP7_75t_L g340 ( .A(n_332), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_335), .B(n_422), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B1(n_344), .B2(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g431 ( .A(n_344), .Y(n_431) );
INVxp33_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_346), .B(n_390), .Y(n_389) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_381), .A3(n_382), .B1(n_383), .B2(n_384), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g348 ( .A(n_349), .B(n_361), .C(n_373), .D(n_385), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp33_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_356), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_386), .B1(n_403), .B2(n_406), .C(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g421 ( .A(n_372), .B(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_377), .B2(n_379), .C(n_380), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_382), .B(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND4xp25_ASAP7_75t_L g391 ( .A(n_392), .B(n_402), .C(n_417), .D(n_428), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B(n_398), .C(n_400), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g433 ( .A(n_420), .Y(n_433) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_433), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_434), .A2(n_445), .B1(n_447), .B2(n_450), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_435), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_437), .B(n_449), .Y(n_736) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g448 ( .A(n_438), .B(n_449), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_440), .A2(n_443), .B(n_738), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g730 ( .A(n_446), .Y(n_730) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx6_ASAP7_75t_L g731 ( .A(n_448), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_450), .Y(n_732) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_451), .B(n_681), .Y(n_450) );
NOR4xp25_ASAP7_75t_L g451 ( .A(n_452), .B(n_618), .C(n_652), .D(n_668), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_453), .B(n_547), .C(n_582), .D(n_598), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_488), .B1(n_522), .B2(n_535), .C1(n_540), .C2(n_546), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI31xp33_ASAP7_75t_L g714 ( .A1(n_455), .A2(n_715), .A3(n_716), .B(n_718), .Y(n_714) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_467), .Y(n_455) );
AND2x2_ASAP7_75t_L g689 ( .A(n_456), .B(n_469), .Y(n_689) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_SL g539 ( .A(n_457), .Y(n_539) );
AND2x2_ASAP7_75t_L g546 ( .A(n_457), .B(n_479), .Y(n_546) );
AND2x2_ASAP7_75t_L g603 ( .A(n_457), .B(n_470), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_467), .B(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_468), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_468), .B(n_550), .Y(n_593) );
AND2x2_ASAP7_75t_L g686 ( .A(n_468), .B(n_626), .Y(n_686) );
OAI321xp33_ASAP7_75t_L g720 ( .A1(n_468), .A2(n_539), .A3(n_693), .B1(n_721), .B2(n_723), .C(n_724), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_468), .B(n_525), .C(n_633), .D(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AND2x2_ASAP7_75t_L g588 ( .A(n_469), .B(n_537), .Y(n_588) );
AND2x2_ASAP7_75t_L g607 ( .A(n_469), .B(n_539), .Y(n_607) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g538 ( .A(n_470), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g563 ( .A(n_470), .B(n_479), .Y(n_563) );
AND2x2_ASAP7_75t_L g649 ( .A(n_470), .B(n_537), .Y(n_649) );
INVx3_ASAP7_75t_SL g537 ( .A(n_479), .Y(n_537) );
AND2x2_ASAP7_75t_L g581 ( .A(n_479), .B(n_568), .Y(n_581) );
OR2x2_ASAP7_75t_L g614 ( .A(n_479), .B(n_539), .Y(n_614) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_479), .Y(n_621) );
AND2x2_ASAP7_75t_L g650 ( .A(n_479), .B(n_538), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_479), .B(n_623), .Y(n_665) );
AND2x2_ASAP7_75t_L g697 ( .A(n_479), .B(n_689), .Y(n_697) );
AND2x2_ASAP7_75t_L g706 ( .A(n_479), .B(n_551), .Y(n_706) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_501), .Y(n_489) );
INVx1_ASAP7_75t_SL g674 ( .A(n_490), .Y(n_674) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g542 ( .A(n_491), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g524 ( .A(n_492), .B(n_503), .Y(n_524) );
AND2x2_ASAP7_75t_L g610 ( .A(n_492), .B(n_526), .Y(n_610) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g580 ( .A(n_493), .B(n_513), .Y(n_580) );
OR2x2_ASAP7_75t_L g591 ( .A(n_493), .B(n_526), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_493), .B(n_526), .Y(n_617) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_493), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_501), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_501), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g590 ( .A(n_502), .B(n_591), .Y(n_590) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_502), .A2(n_580), .A3(n_586), .B1(n_617), .B2(n_667), .C1(n_677), .C2(n_679), .Y(n_676) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_503), .B(n_525), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_503), .B(n_526), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_503), .B(n_543), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_503), .B(n_617), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_503), .Y(n_655) );
AND2x2_ASAP7_75t_L g667 ( .A(n_503), .B(n_513), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_503), .B(n_542), .Y(n_699) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g564 ( .A(n_504), .B(n_513), .Y(n_564) );
BUFx3_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
AND3x2_ASAP7_75t_L g660 ( .A(n_504), .B(n_640), .C(n_661), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_513), .B(n_524), .C(n_525), .Y(n_523) );
INVx1_ASAP7_75t_SL g543 ( .A(n_513), .Y(n_543) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_513), .Y(n_645) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g639 ( .A(n_524), .B(n_640), .Y(n_639) );
INVxp67_ASAP7_75t_L g646 ( .A(n_524), .Y(n_646) );
AND2x2_ASAP7_75t_L g684 ( .A(n_525), .B(n_662), .Y(n_684) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g565 ( .A(n_526), .Y(n_565) );
AND2x2_ASAP7_75t_L g640 ( .A(n_526), .B(n_543), .Y(n_640) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OR2x2_ASAP7_75t_L g584 ( .A(n_537), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g703 ( .A(n_537), .B(n_603), .Y(n_703) );
AND2x2_ASAP7_75t_L g717 ( .A(n_537), .B(n_539), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_538), .B(n_551), .Y(n_658) );
AND2x2_ASAP7_75t_L g705 ( .A(n_538), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g568 ( .A(n_539), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g585 ( .A(n_539), .B(n_551), .Y(n_585) );
INVx1_ASAP7_75t_L g595 ( .A(n_539), .Y(n_595) );
AND2x2_ASAP7_75t_L g626 ( .A(n_539), .B(n_551), .Y(n_626) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_541), .A2(n_669), .B1(n_673), .B2(n_675), .C(n_676), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x2_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_545), .B(n_579), .Y(n_722) );
AOI322xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_564), .A3(n_565), .B1(n_566), .B2(n_572), .C1(n_574), .C2(n_581), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_563), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_550), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_550), .B(n_613), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_550), .A2(n_563), .B(n_637), .C(n_638), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_550), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_550), .B(n_607), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_550), .B(n_689), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_550), .B(n_717), .Y(n_716) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_551), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_551), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g678 ( .A(n_551), .B(n_565), .Y(n_678) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B(n_562), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_553), .A2(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g570 ( .A(n_555), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_562), .Y(n_571) );
INVx1_ASAP7_75t_L g653 ( .A(n_563), .Y(n_653) );
OAI31xp33_ASAP7_75t_L g663 ( .A1(n_563), .A2(n_588), .A3(n_664), .B(n_666), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_563), .B(n_569), .Y(n_715) );
INVx1_ASAP7_75t_SL g576 ( .A(n_564), .Y(n_576) );
AND2x2_ASAP7_75t_L g609 ( .A(n_564), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g690 ( .A(n_564), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g600 ( .A(n_565), .Y(n_600) );
AND2x2_ASAP7_75t_L g627 ( .A(n_565), .B(n_580), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_565), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g719 ( .A(n_565), .B(n_667), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_567), .B(n_637), .Y(n_710) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g624 ( .A(n_569), .Y(n_624) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_575), .B(n_577), .Y(n_574) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_576), .A2(n_619), .B(n_625), .C(n_641), .Y(n_618) );
OR2x2_ASAP7_75t_L g693 ( .A(n_576), .B(n_674), .Y(n_693) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g630 ( .A(n_578), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_578), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g599 ( .A(n_580), .B(n_600), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .B(n_589), .C(n_592), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_SL g633 ( .A(n_585), .Y(n_633) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_588), .B(n_626), .Y(n_631) );
INVx1_ASAP7_75t_L g637 ( .A(n_588), .Y(n_637) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g596 ( .A(n_591), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g629 ( .A(n_591), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g691 ( .A(n_591), .Y(n_691) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B(n_596), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_594), .A2(n_605), .B(n_608), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_601), .B(n_604), .C(n_611), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_599), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_602), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g615 ( .A(n_603), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_605), .A2(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_610), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g635 ( .A(n_610), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_615), .B(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g666 ( .A(n_617), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_623), .B(n_649), .Y(n_675) );
AND2x2_ASAP7_75t_L g688 ( .A(n_623), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g702 ( .A(n_623), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g712 ( .A(n_623), .B(n_650), .Y(n_712) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_628), .C(n_636), .Y(n_625) );
INVx1_ASAP7_75t_L g672 ( .A(n_626), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_632), .B2(n_634), .Y(n_628) );
OR2x2_ASAP7_75t_L g634 ( .A(n_630), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_630), .B(n_691), .Y(n_713) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g707 ( .A(n_640), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_647), .B1(n_650), .B2(n_651), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g725 ( .A(n_645), .Y(n_725) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g671 ( .A(n_649), .Y(n_671) );
OAI211xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B(n_656), .C(n_663), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_671), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NOR5xp2_ASAP7_75t_L g681 ( .A(n_682), .B(n_700), .C(n_708), .D(n_714), .E(n_720), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_685), .B(n_687), .C(n_694), .Y(n_682) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_692), .Y(n_687) );
OAI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_697), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B(n_707), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g723 ( .A(n_703), .Y(n_723) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_711), .B(n_713), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
endmodule