module fake_aes_5020_n_29 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
AND2x2_ASAP7_75t_L g12 ( .A(n_2), .B(n_3), .Y(n_12) );
INVx4_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
AND2x2_ASAP7_75t_SL g14 ( .A(n_5), .B(n_6), .Y(n_14) );
BUFx8_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_13), .B(n_0), .Y(n_17) );
NAND2x1p5_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .Y(n_18) );
OAI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_12), .B(n_13), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_16), .B1(n_12), .B2(n_14), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_1), .Y(n_21) );
OAI222xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_13), .B1(n_15), .B2(n_14), .C1(n_19), .C2(n_1), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_22), .Y(n_23) );
INVxp67_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND4xp25_ASAP7_75t_L g25 ( .A(n_24), .B(n_15), .C(n_4), .D(n_5), .Y(n_25) );
NOR3xp33_ASAP7_75t_L g26 ( .A(n_24), .B(n_19), .C(n_15), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_25), .B1(n_4), .B2(n_9), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_7), .B1(n_10), .B2(n_11), .Y(n_29) );
endmodule