module fake_jpeg_17296_n_20 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_20;

wire n_13;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_2),
.Y(n_10)
);

CKINVDCx12_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_4),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_2),
.A2(n_9),
.B1(n_7),
.B2(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_13),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_16),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.Y(n_16)
);

AOI322xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_13),
.A3(n_11),
.B1(n_8),
.B2(n_5),
.C1(n_4),
.C2(n_3),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_1),
.B1(n_3),
.B2(n_17),
.C(n_15),
.Y(n_20)
);


endmodule