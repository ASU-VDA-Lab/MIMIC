module real_jpeg_10918_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_269;
wire n_96;
wire n_273;
wire n_89;

BUFx24_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_53),
.B1(n_55),
.B2(n_72),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_1),
.A2(n_27),
.B1(n_31),
.B2(n_72),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_72),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_65),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_76),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_76),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_76),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_4),
.B(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_232),
.B(n_256),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_9),
.A2(n_54),
.B1(n_65),
.B2(n_71),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_27),
.B1(n_31),
.B2(n_54),
.Y(n_190)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_11),
.A2(n_65),
.B1(n_71),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_53),
.B1(n_55),
.B2(n_92),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_92),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_27),
.B1(n_31),
.B2(n_92),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_13),
.A2(n_39),
.B1(n_53),
.B2(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_27),
.B1(n_31),
.B2(n_39),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_14),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_15),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_15),
.A2(n_27),
.B1(n_31),
.B2(n_47),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_15),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_16),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_16),
.A2(n_53),
.B(n_67),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_16),
.A2(n_65),
.B1(n_71),
.B2(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_74),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_16),
.A2(n_37),
.B(n_41),
.C(n_200),
.D(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_16),
.B(n_37),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_16),
.B(n_60),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_16),
.A2(n_25),
.B(n_215),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_16),
.A2(n_55),
.B(n_56),
.C(n_149),
.D(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_16),
.B(n_55),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_20),
.B(n_100),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_83),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_21),
.A2(n_22),
.B1(n_77),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_51),
.C(n_62),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_35),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_25),
.A2(n_26),
.B(n_33),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_25),
.A2(n_26),
.B1(n_86),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_25),
.A2(n_26),
.B1(n_143),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_25),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_25),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_25),
.B(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_26),
.A2(n_222),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_26),
.B(n_140),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_27),
.A2(n_44),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_31),
.B(n_42),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_31),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_36),
.A2(n_40),
.B1(n_48),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_37),
.A2(n_248),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_38),
.B(n_58),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_46),
.B1(n_48),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_40),
.A2(n_48),
.B1(n_212),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_40),
.A2(n_246),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_45),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_41),
.B(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_48),
.A2(n_88),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_48),
.B(n_164),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_48),
.A2(n_162),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_48),
.B(n_140),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_57),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_59),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_70),
.B(n_73),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_65),
.A2(n_66),
.B(n_140),
.C(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_69),
.A2(n_91),
.B(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_73),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_77),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_79),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_93),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_85),
.B(n_87),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_99),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_96),
.A2(n_146),
.B1(n_147),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_96),
.A2(n_97),
.B(n_170),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_123),
.B2(n_124),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_112),
.B2(n_113),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_111),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_109),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_122),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_153),
.B(n_279),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_150),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_129),
.B(n_150),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_133),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_132),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_134),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_144),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_136),
.B1(n_144),
.B2(n_145),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_192),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_176),
.B(n_191),
.Y(n_155)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_156),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_173),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_173),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.CI(n_171),
.CON(n_157),
.SN(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.C(n_168),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_161),
.B1(n_168),
.B2(n_169),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_177),
.B(n_178),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_183),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_179),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_181),
.A2(n_183),
.B1(n_184),
.B2(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_181),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_188),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_185),
.A2(n_186),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_187),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_190),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_277),
.C(n_278),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_271),
.B(n_276),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_259),
.B(n_270),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_240),
.B(n_258),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_218),
.B(n_239),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_200),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_201),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_238),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_225),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_242),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_257),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_250),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_251),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_267),
.C(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);


endmodule