module fake_jpeg_4485_n_37 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_37);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_17),
.B(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_10),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_0),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_9),
.B1(n_1),
.B2(n_3),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_33),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_32),
.B(n_23),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_18),
.B(n_19),
.Y(n_37)
);


endmodule