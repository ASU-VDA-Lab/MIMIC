module fake_aes_6860_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx4_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
BUFx3_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OA21x2_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
OAI21xp5_ASAP7_75t_SL g9 ( .A1(n_7), .A2(n_3), .B(n_4), .Y(n_9) );
AOI211xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B(n_3), .C(n_2), .Y(n_10) );
AOI221xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_5), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_11), .B(n_5), .Y(n_13) );
endmodule