module real_jpeg_4673_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_1),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_1),
.A2(n_125),
.B1(n_153),
.B2(n_288),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_1),
.A2(n_153),
.B1(n_281),
.B2(n_320),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_1),
.A2(n_61),
.B1(n_153),
.B2(n_231),
.Y(n_375)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_2),
.A2(n_271),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_2),
.B(n_315),
.C(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_2),
.B(n_110),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_2),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_2),
.B(n_92),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_2),
.B(n_382),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_4),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_59),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_4),
.A2(n_59),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_6),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_6),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_6),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_9),
.A2(n_47),
.B1(n_87),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_87),
.B1(n_119),
.B2(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_10),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_11),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_11),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_11),
.A2(n_55),
.B1(n_124),
.B2(n_186),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_11),
.A2(n_124),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_11),
.A2(n_124),
.B1(n_389),
.B2(n_391),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_12),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_12),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_12),
.A2(n_157),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_12),
.A2(n_157),
.B1(n_231),
.B2(n_308),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_12),
.A2(n_157),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_13),
.A2(n_60),
.B1(n_202),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_13),
.A2(n_202),
.B1(n_325),
.B2(n_352),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_13),
.A2(n_202),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_14),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_15),
.A2(n_37),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_16),
.A2(n_45),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_249),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_248),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_215),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_20),
.B(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_164),
.C(n_181),
.Y(n_20)
);

FAx1_ASAP7_75t_L g290 ( 
.A(n_21),
.B(n_164),
.CI(n_181),
.CON(n_290),
.SN(n_290)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_22),
.B(n_94),
.C(n_134),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_23),
.B(n_53),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_42),
.B2(n_44),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_24),
.A2(n_44),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_24),
.A2(n_277),
.B1(n_283),
.B2(n_284),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_24),
.A2(n_319),
.B(n_322),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_24),
.A2(n_271),
.B(n_322),
.Y(n_348)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_25),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_25),
.B(n_324),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_25),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_25),
.A2(n_195),
.B1(n_278),
.B2(n_388),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_26),
.Y(n_356)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_27),
.Y(n_196)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_28),
.Y(n_327)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_30),
.Y(n_279)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_30),
.Y(n_392)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_31),
.Y(n_194)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_35),
.Y(n_345)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_35),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_36),
.Y(n_193)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_38),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_41),
.Y(n_321)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_42),
.Y(n_364)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_51),
.Y(n_282)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_52),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_65),
.B1(n_86),
.B2(n_92),
.Y(n_53)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_54),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_58),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_58),
.Y(n_231)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_58),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_64),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_64),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_64),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_65),
.A2(n_86),
.B1(n_92),
.B2(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_65),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_65),
.A2(n_92),
.B1(n_167),
.B2(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_65),
.B(n_307),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_75),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_74),
.Y(n_397)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_75),
.A2(n_331),
.B(n_335),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_89),
.Y(n_232)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g400 ( 
.A(n_90),
.B(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_91),
.Y(n_313)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_92),
.B(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_134),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_118),
.B1(n_127),
.B2(n_128),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_95),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_95),
.A2(n_127),
.B1(n_287),
.B2(n_412),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_110),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_99),
.B1(n_104),
.B2(n_107),
.Y(n_96)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_97),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_99),
.Y(n_210)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_102),
.Y(n_226)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_102),
.Y(n_263)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_102),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_103),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_106),
.Y(n_399)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

AOI22x1_ASAP7_75t_L g206 ( 
.A1(n_110),
.A2(n_207),
.B1(n_208),
.B2(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_110),
.A2(n_207),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_122),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

AOI32xp33_ASAP7_75t_L g394 ( 
.A1(n_125),
.A2(n_381),
.A3(n_395),
.B1(n_398),
.B2(n_400),
.Y(n_394)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_127),
.B(n_209),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_127),
.A2(n_412),
.B(n_415),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_151),
.B(n_155),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_151),
.B1(n_199),
.B2(n_205),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_136),
.B(n_156),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_136),
.A2(n_433),
.B(n_435),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx8_ASAP7_75t_L g434 ( 
.A(n_139),
.Y(n_434)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_155),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_162),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_176),
.B2(n_180),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_166),
.B(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_180),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_197),
.C(n_206),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_183),
.B(n_190),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_184),
.A2(n_300),
.B(n_306),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_184),
.A2(n_188),
.B1(n_331),
.B2(n_375),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_184),
.A2(n_306),
.B(n_375),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_185),
.A2(n_188),
.B(n_335),
.Y(n_438)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_193),
.Y(n_326)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_197),
.A2(n_198),
.B1(n_206),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_199),
.A2(n_205),
.B(n_247),
.Y(n_260)
);

OAI32xp33_ASAP7_75t_L g262 ( 
.A1(n_200),
.A2(n_263),
.A3(n_264),
.B1(n_266),
.B2(n_270),
.Y(n_262)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_205),
.B(n_271),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_206),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_207),
.A2(n_286),
.B(n_289),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_207),
.A2(n_289),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_207),
.B(n_208),
.Y(n_415)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_212),
.Y(n_414)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_234),
.B2(n_235),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B(n_233),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_228),
.Y(n_233)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_291),
.B(n_463),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_290),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_252),
.B(n_290),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_258),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_257),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_258),
.B(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.C(n_285),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_259),
.A2(n_260),
.B1(n_285),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_261),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_275),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_262),
.A2(n_275),
.B1(n_276),
.B2(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_262),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_SL g433 ( 
.A1(n_270),
.A2(n_271),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g378 ( 
.A1(n_271),
.A2(n_379),
.B(n_380),
.Y(n_378)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_285),
.Y(n_448)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_290),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_441),
.B(n_460),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_421),
.B(n_440),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_403),
.B(n_420),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_369),
.B(n_402),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_338),
.B(n_368),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_317),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_317),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_309),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_299),
.A2(n_309),
.B1(n_310),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_328),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_329),
.C(n_337),
.Y(n_370)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_336),
.B2(n_337),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx11_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_360),
.B(n_367),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_349),
.B(n_359),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_348),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_358),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_358),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_355),
.B(n_357),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_387),
.B(n_393),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_365),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_371),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_385),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_376),
.C(n_385),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx5_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_404),
.B(n_405),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_410),
.B2(n_419),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_409),
.C(n_419),
.Y(n_422)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_410),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_416),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_417),
.C(n_418),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_422),
.B(n_423),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_430),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_425),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_427),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_428),
.C(n_430),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_436),
.B2(n_439),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_437),
.C(n_438),
.Y(n_451)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_455),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_444),
.A2(n_461),
.B(n_462),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_452),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_452),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.C(n_451),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_449),
.A2(n_450),
.B1(n_451),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_451),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_457),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);


endmodule