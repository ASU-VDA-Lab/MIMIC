module fake_ariane_1655_n_2220 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2220);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2220;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_1682;
wire n_1836;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_1985;
wire n_995;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_661;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_1924;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_1432;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_2185;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_632;
wire n_650;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_1578;
wire n_1455;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2168;
wire n_670;
wire n_1826;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_2075;
wire n_1726;
wire n_1945;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_1005;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_1281;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_802;
wire n_1151;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2143;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_748;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_1344;
wire n_1390;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_1150;
wire n_977;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_1136;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_937;
wire n_1474;
wire n_2081;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_849;
wire n_2095;
wire n_1820;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_573;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g564 ( 
.A(n_125),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_56),
.Y(n_565)
);

BUFx5_ASAP7_75t_L g566 ( 
.A(n_310),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_25),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_251),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_460),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_137),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_334),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_130),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_422),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_340),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_104),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_5),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_114),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_342),
.Y(n_578)
);

BUFx5_ASAP7_75t_L g579 ( 
.A(n_3),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_121),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_166),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_191),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_430),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_134),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_537),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_214),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_428),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_145),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_62),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_96),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_227),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_427),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_99),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_170),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_221),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_295),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_8),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_122),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_382),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_58),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_432),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_506),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_159),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_494),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_429),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

INVxp33_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_434),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_561),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_140),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_521),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_335),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_67),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_532),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_33),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_131),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_251),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_388),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_398),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_488),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_107),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_420),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_493),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_418),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_104),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_333),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_162),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_306),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_16),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_196),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_260),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_187),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_146),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_313),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_86),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_70),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_60),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_61),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_261),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_545),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_451),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_236),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_282),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_503),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_76),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_470),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_97),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_108),
.Y(n_648)
);

BUFx8_ASAP7_75t_SL g649 ( 
.A(n_540),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_234),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_122),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_486),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_482),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_44),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_309),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_118),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_112),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_379),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_107),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_524),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_153),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_403),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_1),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_148),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_483),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_554),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_465),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_305),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_57),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_115),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_61),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_279),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_94),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_400),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_229),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_68),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_421),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_459),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_108),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_261),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_85),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_55),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_109),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_134),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_175),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_68),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_46),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_153),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_511),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_461),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_20),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_152),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_480),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_278),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_347),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_283),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_226),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_536),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_373),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_513),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_395),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_198),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_257),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_139),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_360),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_237),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_151),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_277),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_27),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_416),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_237),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_258),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_53),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_125),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_453),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_546),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_116),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_241),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_292),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_222),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_452),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_563),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_411),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_278),
.Y(n_724)
);

BUFx10_ASAP7_75t_L g725 ( 
.A(n_248),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_135),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_219),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_284),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_28),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_520),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_161),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_476),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_391),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_329),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_203),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_202),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_168),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_225),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_389),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_302),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_37),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_243),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_338),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_228),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_528),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_535),
.Y(n_746)
);

BUFx10_ASAP7_75t_L g747 ( 
.A(n_228),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_311),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_4),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_529),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_241),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_238),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_62),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_157),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_43),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_355),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_385),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_455),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_36),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_231),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_276),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_357),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_326),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_462),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_566),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_566),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_568),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_568),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_566),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_566),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_621),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_638),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_685),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_606),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_566),
.Y(n_775)
);

INVxp33_ASAP7_75t_SL g776 ( 
.A(n_703),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_564),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_621),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_630),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_680),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_680),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_726),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_726),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_566),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_569),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_602),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_712),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_685),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_566),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_579),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_619),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_579),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_579),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_718),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_672),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_763),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_579),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_624),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_763),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_579),
.Y(n_801)
);

INVxp33_ASAP7_75t_SL g802 ( 
.A(n_574),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_718),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_579),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_716),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_579),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_576),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_581),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_649),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_584),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_649),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_591),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_595),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_596),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_596),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_755),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_616),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_755),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_596),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_636),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_656),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_693),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_657),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_596),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_661),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_668),
.Y(n_827)
);

CKINVDCx16_ASAP7_75t_R g828 ( 
.A(n_673),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_688),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_704),
.Y(n_831)
);

INVxp33_ASAP7_75t_SL g832 ( 
.A(n_567),
.Y(n_832)
);

CKINVDCx16_ASAP7_75t_R g833 ( 
.A(n_673),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_706),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_623),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_693),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_707),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_709),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_728),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_583),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_565),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_735),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_749),
.Y(n_843)
);

INVxp67_ASAP7_75t_SL g844 ( 
.A(n_663),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_663),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_594),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_583),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_760),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_600),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_597),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_663),
.Y(n_851)
);

INVxp33_ASAP7_75t_SL g852 ( 
.A(n_570),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_583),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_769),
.A2(n_640),
.B(n_626),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_840),
.B(n_607),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_769),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_844),
.B(n_674),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_840),
.B(n_677),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_770),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_765),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_815),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_770),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_816),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_773),
.A2(n_740),
.B1(n_748),
.B2(n_632),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_847),
.B(n_678),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_775),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_847),
.B(n_698),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_801),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_802),
.B(n_607),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_848),
.B(n_673),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_765),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_853),
.B(n_701),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_775),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_816),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_853),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_705),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_767),
.B(n_725),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_794),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_794),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_766),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_787),
.B(n_721),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_798),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_804),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_792),
.B(n_732),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_825),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_825),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_766),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_792),
.B(n_733),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_845),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_776),
.A2(n_802),
.B1(n_796),
.B2(n_777),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_835),
.B(n_597),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_798),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_845),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_785),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_785),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_820),
.Y(n_897)
);

INVx3_ASAP7_75t_L g898 ( 
.A(n_820),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_835),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_776),
.A2(n_729),
.B1(n_727),
.B2(n_648),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_774),
.B(n_768),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_774),
.B(n_627),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_790),
.Y(n_903)
);

AO22x1_ASAP7_75t_L g904 ( 
.A1(n_772),
.A2(n_631),
.B1(n_655),
.B2(n_627),
.Y(n_904)
);

CKINVDCx14_ASAP7_75t_R g905 ( 
.A(n_809),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_851),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_806),
.A2(n_758),
.B(n_743),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_851),
.Y(n_908)
);

XNOR2x2_ASAP7_75t_L g909 ( 
.A(n_773),
.B(n_737),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_791),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_809),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_786),
.A2(n_741),
.B1(n_708),
.B2(n_659),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_791),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_869),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_869),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_905),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_912),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_912),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_876),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_876),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_869),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_884),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_855),
.B(n_786),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_865),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_884),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_865),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_891),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_861),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_856),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_870),
.B(n_811),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_R g933 ( 
.A(n_859),
.B(n_811),
.Y(n_933)
);

XOR2x2_ASAP7_75t_L g934 ( 
.A(n_909),
.B(n_789),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_871),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_866),
.Y(n_936)
);

INVxp33_ASAP7_75t_SL g937 ( 
.A(n_871),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_861),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_900),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_856),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_872),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_872),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_868),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_913),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_878),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_860),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_873),
.B(n_799),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_901),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_881),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_R g950 ( 
.A(n_881),
.B(n_799),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_909),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_860),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_888),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_888),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_878),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_901),
.Y(n_956)
);

CKINVDCx16_ASAP7_75t_R g957 ( 
.A(n_901),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_863),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_901),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_863),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_895),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_858),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_902),
.B(n_805),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_902),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_902),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_902),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_857),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_877),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_882),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_885),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_889),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_896),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_914),
.B(n_805),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_892),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_R g976 ( 
.A(n_896),
.B(n_823),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_867),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_892),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_914),
.B(n_793),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_892),
.Y(n_980)
);

CKINVDCx16_ASAP7_75t_R g981 ( 
.A(n_892),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_903),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_904),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_903),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_911),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_911),
.B(n_823),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_910),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_R g988 ( 
.A(n_899),
.B(n_836),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_858),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_867),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_904),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_899),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_898),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_910),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_899),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_914),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_874),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_935),
.B(n_788),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_976),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_936),
.B(n_832),
.Y(n_1002)
);

INVx4_ASAP7_75t_L g1003 ( 
.A(n_916),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_930),
.B(n_959),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_R g1005 ( 
.A(n_917),
.B(n_836),
.Y(n_1005)
);

AND2x6_ASAP7_75t_L g1006 ( 
.A(n_941),
.B(n_578),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_918),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_938),
.B(n_874),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_942),
.B(n_880),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_916),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_937),
.B(n_832),
.Y(n_1011)
);

AND2x6_ASAP7_75t_L g1012 ( 
.A(n_953),
.B(n_578),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_953),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_919),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_937),
.B(n_852),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_931),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_949),
.B(n_880),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_954),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_920),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_967),
.B(n_807),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_962),
.B(n_883),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_920),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_921),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_986),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_SL g1025 ( 
.A(n_921),
.B(n_585),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_973),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_940),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_982),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_978),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_984),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_957),
.B(n_828),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_943),
.B(n_852),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_939),
.A2(n_655),
.B1(n_681),
.B2(n_631),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_985),
.B(n_883),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_987),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_945),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_963),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_968),
.B(n_833),
.Y(n_1038)
);

INVx4_ASAP7_75t_L g1039 ( 
.A(n_980),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_955),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_915),
.B(n_604),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_997),
.B(n_893),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_950),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_960),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_946),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_946),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_995),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_974),
.B(n_899),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_952),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_955),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_952),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_975),
.B(n_981),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_998),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_948),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_963),
.Y(n_1055)
);

AND2x6_ASAP7_75t_L g1056 ( 
.A(n_922),
.B(n_604),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_969),
.B(n_899),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_970),
.B(n_841),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_971),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_956),
.Y(n_1060)
);

NAND3x1_ASAP7_75t_L g1061 ( 
.A(n_924),
.B(n_795),
.C(n_789),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_923),
.B(n_899),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_965),
.B(n_808),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_926),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_958),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_963),
.Y(n_1066)
);

INVx6_ASAP7_75t_L g1067 ( 
.A(n_963),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_961),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_929),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_999),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_961),
.Y(n_1071)
);

NAND3x1_ASAP7_75t_L g1072 ( 
.A(n_928),
.B(n_803),
.C(n_795),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_977),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_989),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_966),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_972),
.B(n_893),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_991),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_983),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_991),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_979),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_989),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_947),
.B(n_599),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_939),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_994),
.B(n_907),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_989),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_989),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_990),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_990),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_990),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_990),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_932),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_992),
.B(n_907),
.Y(n_1092)
);

INVx5_ASAP7_75t_L g1093 ( 
.A(n_988),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_996),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_964),
.B(n_992),
.Y(n_1095)
);

BUFx10_ASAP7_75t_L g1096 ( 
.A(n_927),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_944),
.B(n_841),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_996),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_993),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_849),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_951),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_951),
.Y(n_1103)
);

AND2x6_ASAP7_75t_L g1104 ( 
.A(n_933),
.B(n_611),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_925),
.B(n_849),
.Y(n_1105)
);

BUFx10_ASAP7_75t_L g1106 ( 
.A(n_925),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_934),
.B(n_575),
.C(n_572),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_934),
.B(n_644),
.Y(n_1108)
);

AO22x2_ASAP7_75t_L g1109 ( 
.A1(n_934),
.A2(n_817),
.B1(n_819),
.B2(n_803),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_941),
.Y(n_1110)
);

AND2x6_ASAP7_75t_L g1111 ( 
.A(n_941),
.B(n_611),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_941),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_935),
.B(n_846),
.Y(n_1113)
);

CKINVDCx14_ASAP7_75t_R g1114 ( 
.A(n_917),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_931),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_916),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_930),
.B(n_907),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_917),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_967),
.B(n_810),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_930),
.B(n_907),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_930),
.B(n_793),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_930),
.B(n_854),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_916),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_957),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_930),
.B(n_854),
.Y(n_1125)
);

OAI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_939),
.A2(n_691),
.B1(n_719),
.B2(n_681),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_916),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_1001),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1076),
.B(n_653),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1067),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_1059),
.B(n_662),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1080),
.B(n_879),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_1052),
.B(n_818),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1018),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_L g1135 ( 
.A(n_1011),
.B(n_819),
.C(n_817),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1024),
.B(n_577),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_L g1137 ( 
.A(n_1093),
.B(n_580),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1015),
.B(n_582),
.Y(n_1138)
);

INVx8_ASAP7_75t_L g1139 ( 
.A(n_1124),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1026),
.Y(n_1140)
);

AND2x6_ASAP7_75t_SL g1141 ( 
.A(n_1058),
.B(n_812),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1076),
.B(n_898),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1045),
.Y(n_1143)
);

INVxp33_ASAP7_75t_L g1144 ( 
.A(n_1098),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1023),
.B(n_586),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1028),
.Y(n_1146)
);

NAND2x1p5_ASAP7_75t_L g1147 ( 
.A(n_1124),
.B(n_898),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1124),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1038),
.B(n_691),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1045),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1044),
.A2(n_588),
.B1(n_590),
.B2(n_589),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1023),
.B(n_593),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1030),
.B(n_1020),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1020),
.B(n_719),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1119),
.B(n_753),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1119),
.B(n_753),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1004),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1093),
.B(n_598),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1004),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1107),
.A2(n_608),
.B1(n_731),
.B2(n_725),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1063),
.B(n_886),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_886),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1104),
.B(n_886),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1078),
.B(n_813),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1054),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1022),
.B(n_610),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1019),
.B(n_613),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1060),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1002),
.B(n_615),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1032),
.B(n_617),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1044),
.B(n_625),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1104),
.B(n_628),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_1107),
.B(n_663),
.Y(n_1173)
);

INVx8_ASAP7_75t_L g1174 ( 
.A(n_1093),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1043),
.B(n_629),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1053),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1104),
.B(n_633),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1050),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1036),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1013),
.B(n_634),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1008),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1008),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1084),
.A2(n_660),
.B(n_696),
.C(n_669),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_1031),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1110),
.B(n_635),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1007),
.B(n_637),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1014),
.B(n_639),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1025),
.A2(n_642),
.B1(n_645),
.B2(n_643),
.Y(n_1188)
);

INVx8_ASAP7_75t_L g1189 ( 
.A(n_1006),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1113),
.B(n_771),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1095),
.B(n_647),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1112),
.B(n_650),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1105),
.A2(n_651),
.B1(n_670),
.B2(n_664),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1050),
.B(n_654),
.Y(n_1194)
);

AND2x6_ASAP7_75t_SL g1195 ( 
.A(n_1101),
.B(n_814),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1092),
.B(n_879),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1000),
.B(n_778),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1082),
.B(n_671),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_1118),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1092),
.B(n_879),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1029),
.B(n_821),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1121),
.B(n_879),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1096),
.B(n_779),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1039),
.B(n_675),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1035),
.B(n_676),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1091),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1047),
.B(n_679),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1123),
.B(n_682),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1073),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1039),
.B(n_684),
.Y(n_1210)
);

OR2x6_ASAP7_75t_L g1211 ( 
.A(n_1100),
.B(n_843),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1042),
.A2(n_1125),
.B(n_1122),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1123),
.B(n_686),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1073),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1040),
.B(n_780),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1042),
.A2(n_879),
.B(n_573),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1075),
.B(n_1097),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1075),
.Y(n_1218)
);

NAND3xp33_ASAP7_75t_L g1219 ( 
.A(n_1005),
.B(n_1069),
.C(n_1064),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1122),
.A2(n_879),
.B(n_592),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1077),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1126),
.A2(n_608),
.B1(n_731),
.B2(n_725),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1003),
.B(n_692),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1016),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1006),
.B(n_694),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1006),
.B(n_697),
.Y(n_1226)
);

NOR3xp33_ASAP7_75t_L g1227 ( 
.A(n_1114),
.B(n_711),
.C(n_702),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1003),
.B(n_713),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1006),
.B(n_717),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1096),
.B(n_781),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1100),
.A2(n_734),
.B1(n_738),
.B2(n_720),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1012),
.B(n_724),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1012),
.B(n_742),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1100),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1009),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1037),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1037),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1102),
.A2(n_752),
.B1(n_754),
.B2(n_744),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_SL g1239 ( 
.A(n_1106),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1010),
.B(n_751),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1084),
.A2(n_660),
.B(n_761),
.C(n_759),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1012),
.B(n_782),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1103),
.A2(n_608),
.B1(n_736),
.B2(n_731),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1012),
.B(n_783),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1121),
.A2(n_714),
.B1(n_683),
.B2(n_822),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1111),
.B(n_784),
.Y(n_1246)
);

INVxp33_ASAP7_75t_L g1247 ( 
.A(n_1109),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1070),
.A2(n_641),
.B(n_826),
.C(n_824),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1010),
.B(n_714),
.C(n_683),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1111),
.A2(n_587),
.B1(n_646),
.B2(n_622),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1083),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1061),
.B(n_839),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1111),
.B(n_1127),
.Y(n_1253)
);

NOR3xp33_ASAP7_75t_L g1254 ( 
.A(n_1033),
.B(n_1116),
.C(n_1127),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1009),
.B(n_665),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1111),
.B(n_722),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1017),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1017),
.B(n_897),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1021),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1021),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1106),
.B(n_747),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1034),
.B(n_897),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1109),
.B(n_797),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1037),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1099),
.B(n_747),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1108),
.B(n_800),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1071),
.A2(n_714),
.B1(n_683),
.B2(n_827),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1041),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1125),
.A2(n_1120),
.B(n_1117),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1094),
.B(n_829),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1034),
.B(n_830),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1041),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1048),
.A2(n_601),
.B(n_571),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1094),
.B(n_831),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1079),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1027),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1088),
.B(n_834),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1057),
.B(n_714),
.C(n_837),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1067),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1046),
.B(n_838),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1055),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1049),
.B(n_897),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1087),
.B(n_605),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1051),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1065),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1068),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1041),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1041),
.B(n_842),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1056),
.B(n_850),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1056),
.B(n_897),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1056),
.B(n_897),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1056),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1089),
.B(n_609),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1115),
.B(n_906),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1055),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1117),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1089),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1090),
.B(n_906),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1081),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1085),
.B(n_906),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1055),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1066),
.B(n_612),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1066),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1089),
.B(n_614),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1074),
.B(n_618),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1074),
.B(n_908),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1074),
.B(n_908),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1212),
.A2(n_1086),
.B(n_1062),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_1072),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1153),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1144),
.B(n_1086),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1157),
.B(n_1159),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1138),
.B(n_1086),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1269),
.A2(n_1062),
.B(n_764),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1139),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1178),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1217),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1129),
.B(n_908),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1224),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1270),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1220),
.A2(n_862),
.B(n_858),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1269),
.A2(n_658),
.B(n_652),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_L g1323 ( 
.A(n_1199),
.B(n_1206),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1202),
.A2(n_667),
.B(n_666),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_L g1325 ( 
.A(n_1139),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1128),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1133),
.B(n_908),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1166),
.A2(n_3),
.B(n_0),
.C(n_2),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1202),
.A2(n_690),
.B(n_689),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1134),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1133),
.B(n_858),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1296),
.A2(n_700),
.B(n_699),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1181),
.B(n_4),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1239),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_R g1335 ( 
.A(n_1174),
.B(n_710),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1258),
.A2(n_695),
.B(n_862),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1182),
.B(n_5),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1173),
.A2(n_723),
.B1(n_730),
.B2(n_715),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1140),
.Y(n_1339)
);

INVx11_ASAP7_75t_L g1340 ( 
.A(n_1128),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1279),
.B(n_1211),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1235),
.B(n_6),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1284),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1211),
.B(n_862),
.Y(n_1344)
);

INVx11_ASAP7_75t_L g1345 ( 
.A(n_1139),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1174),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1257),
.B(n_6),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1191),
.A2(n_745),
.B1(n_750),
.B2(n_739),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1259),
.B(n_7),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1218),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1146),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1171),
.B(n_756),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1260),
.B(n_7),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1258),
.A2(n_762),
.B(n_757),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1197),
.B(n_862),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1190),
.B(n_8),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1255),
.B(n_9),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1255),
.B(n_1271),
.Y(n_1358)
);

CKINVDCx10_ASAP7_75t_R g1359 ( 
.A(n_1239),
.Y(n_1359)
);

INVxp67_ASAP7_75t_R g1360 ( 
.A(n_1148),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1297),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1262),
.A2(n_746),
.B(n_620),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1254),
.A2(n_864),
.B1(n_875),
.B2(n_862),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1285),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1216),
.A2(n_746),
.B(n_620),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_1149),
.B(n_1277),
.C(n_1170),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1196),
.A2(n_875),
.B(n_864),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1169),
.A2(n_875),
.B(n_887),
.C(n_864),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1280),
.B(n_9),
.Y(n_1369)
);

AO21x1_ASAP7_75t_L g1370 ( 
.A1(n_1245),
.A2(n_695),
.B(n_864),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1165),
.Y(n_1371)
);

NAND2x1p5_ASAP7_75t_L g1372 ( 
.A(n_1179),
.B(n_875),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1266),
.B(n_10),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1168),
.B(n_10),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1132),
.A2(n_746),
.B(n_620),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1132),
.A2(n_746),
.B(n_620),
.Y(n_1377)
);

OAI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1183),
.A2(n_695),
.B(n_887),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1142),
.A2(n_890),
.B(n_887),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1141),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1195),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1156),
.B(n_1164),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1176),
.Y(n_1383)
);

NOR2x1p5_ASAP7_75t_SL g1384 ( 
.A(n_1143),
.B(n_695),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1189),
.B(n_887),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1286),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1186),
.B(n_11),
.C(n_12),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1164),
.B(n_11),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1274),
.B(n_12),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1298),
.A2(n_894),
.B(n_890),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1201),
.B(n_13),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1187),
.B(n_13),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1196),
.A2(n_894),
.B(n_890),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1201),
.B(n_890),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1231),
.B(n_890),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1241),
.A2(n_695),
.B(n_894),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1200),
.A2(n_894),
.B(n_330),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1219),
.A2(n_894),
.B(n_695),
.C(n_16),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1275),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1150),
.A2(n_695),
.B(n_14),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1251),
.B(n_14),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1184),
.B(n_15),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1167),
.B(n_15),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1203),
.B(n_17),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1230),
.B(n_17),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1256),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1250),
.A2(n_21),
.B(n_18),
.C(n_19),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1194),
.B(n_1261),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1276),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1238),
.A2(n_1248),
.B(n_1213),
.C(n_1208),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1161),
.B(n_22),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1174),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1256),
.B(n_22),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1162),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1290),
.A2(n_332),
.B(n_331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1222),
.B(n_23),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1131),
.B(n_24),
.Y(n_1417)
);

INVx11_ASAP7_75t_L g1418 ( 
.A(n_1234),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1306),
.A2(n_337),
.B(n_336),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1205),
.B(n_24),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1215),
.B(n_25),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1237),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1237),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1207),
.B(n_26),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1302),
.B(n_26),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1297),
.B(n_1151),
.Y(n_1426)
);

NOR3xp33_ASAP7_75t_L g1427 ( 
.A(n_1193),
.B(n_27),
.C(n_28),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1306),
.A2(n_1307),
.B(n_1300),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1130),
.B(n_29),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1253),
.A2(n_341),
.B(n_339),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1130),
.B(n_30),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1209),
.B(n_30),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1214),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1263),
.B(n_31),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1282),
.A2(n_344),
.B(n_343),
.Y(n_1435)
);

CKINVDCx8_ASAP7_75t_R g1436 ( 
.A(n_1252),
.Y(n_1436)
);

NOR2x2_ASAP7_75t_L g1437 ( 
.A(n_1252),
.B(n_31),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1160),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_1252),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1221),
.B(n_34),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1294),
.A2(n_1189),
.B(n_1223),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1237),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1264),
.Y(n_1443)
);

NOR3xp33_ASAP7_75t_L g1444 ( 
.A(n_1265),
.B(n_35),
.C(n_36),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1180),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1299),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1288),
.B(n_38),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1189),
.A2(n_1240),
.B(n_1228),
.Y(n_1448)
);

NAND2xp33_ASAP7_75t_L g1449 ( 
.A(n_1264),
.B(n_39),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1185),
.B(n_1192),
.Y(n_1450)
);

AO21x1_ASAP7_75t_L g1451 ( 
.A1(n_1245),
.A2(n_346),
.B(n_345),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1147),
.B(n_1243),
.Y(n_1452)
);

INVx11_ASAP7_75t_L g1453 ( 
.A(n_1137),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1147),
.B(n_39),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1136),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1172),
.B(n_40),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1291),
.A2(n_349),
.B(n_348),
.Y(n_1457)
);

BUFx12f_ASAP7_75t_L g1458 ( 
.A(n_1264),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1177),
.B(n_40),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1281),
.B(n_41),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1268),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1242),
.B(n_42),
.Y(n_1462)
);

AO22x1_ASAP7_75t_L g1463 ( 
.A1(n_1227),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1281),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1281),
.B(n_45),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1295),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1244),
.B(n_48),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1236),
.A2(n_351),
.B(n_350),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1305),
.A2(n_353),
.B(n_352),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1295),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1301),
.A2(n_356),
.B(n_354),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1303),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1289),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1188),
.A2(n_48),
.B(n_49),
.Y(n_1474)
);

AOI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1163),
.A2(n_1278),
.B(n_1246),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1225),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1295),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1145),
.A2(n_359),
.B(n_358),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1247),
.B(n_50),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1226),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1158),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1272),
.A2(n_54),
.B1(n_51),
.B2(n_52),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1152),
.B(n_52),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1229),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1204),
.B(n_55),
.Y(n_1485)
);

NOR2x1p5_ASAP7_75t_SL g1486 ( 
.A(n_1249),
.B(n_361),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1232),
.B(n_56),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1233),
.B(n_57),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1210),
.B(n_1175),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1283),
.A2(n_1304),
.B(n_1293),
.Y(n_1490)
);

O2A1O1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1273),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1287),
.B(n_59),
.Y(n_1492)
);

INVx5_ASAP7_75t_L g1493 ( 
.A(n_1458),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1408),
.B(n_1292),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1341),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1464),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1325),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1308),
.A2(n_1267),
.B(n_363),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1367),
.A2(n_364),
.B(n_362),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1309),
.A2(n_1352),
.B1(n_1338),
.B2(n_1474),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1350),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1317),
.B(n_63),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1358),
.B(n_63),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1316),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_SL g1505 ( 
.A(n_1392),
.B(n_64),
.C(n_65),
.Y(n_1505)
);

O2A1O1Ixp5_ASAP7_75t_L g1506 ( 
.A1(n_1425),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1371),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1326),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1312),
.B(n_67),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1341),
.B(n_69),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1310),
.B(n_69),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1366),
.B(n_70),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1313),
.B(n_71),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1330),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1382),
.B(n_71),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1421),
.B(n_72),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1359),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_R g1518 ( 
.A(n_1325),
.B(n_365),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1385),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1379),
.A2(n_367),
.B(n_366),
.Y(n_1520)
);

NOR2xp67_ASAP7_75t_SL g1521 ( 
.A(n_1380),
.B(n_72),
.Y(n_1521)
);

AOI22x1_ASAP7_75t_L g1522 ( 
.A1(n_1324),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1319),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_369),
.B(n_368),
.Y(n_1524)
);

AO32x1_ASAP7_75t_L g1525 ( 
.A1(n_1445),
.A2(n_75),
.A3(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1315),
.B(n_370),
.Y(n_1526)
);

O2A1O1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1403),
.A2(n_1373),
.B(n_1387),
.C(n_1427),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1328),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.C(n_80),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1311),
.B(n_78),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1376),
.B(n_79),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1450),
.B(n_1414),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1339),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1351),
.B(n_1383),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1356),
.B(n_81),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1428),
.A2(n_372),
.B(n_371),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1410),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1397),
.A2(n_375),
.B(n_374),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1348),
.B(n_82),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1348),
.B(n_83),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1399),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1338),
.B(n_84),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1385),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1474),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1446),
.B(n_87),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1335),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1365),
.A2(n_377),
.B(n_376),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1357),
.B(n_88),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_R g1548 ( 
.A(n_1359),
.B(n_378),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1409),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1417),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1550)
);

BUFx3_ASAP7_75t_L g1551 ( 
.A(n_1315),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1453),
.B(n_89),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1455),
.B(n_90),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1327),
.B(n_91),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_R g1555 ( 
.A(n_1346),
.B(n_380),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1420),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1343),
.Y(n_1557)
);

CKINVDCx8_ASAP7_75t_R g1558 ( 
.A(n_1315),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1340),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1364),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1369),
.B(n_92),
.Y(n_1561)
);

BUFx2_ASAP7_75t_SL g1562 ( 
.A(n_1323),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1404),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1332),
.B(n_93),
.Y(n_1564)
);

AOI33xp33_ASAP7_75t_L g1565 ( 
.A1(n_1438),
.A2(n_97),
.A3(n_99),
.B1(n_95),
.B2(n_96),
.B3(n_98),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1434),
.B(n_1381),
.Y(n_1566)
);

NAND3xp33_ASAP7_75t_L g1567 ( 
.A(n_1406),
.B(n_1320),
.C(n_1407),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1346),
.B(n_381),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1418),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1385),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1386),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1314),
.A2(n_384),
.B(n_383),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1484),
.B(n_95),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1390),
.A2(n_387),
.B(n_386),
.Y(n_1574)
);

NOR3xp33_ASAP7_75t_L g1575 ( 
.A(n_1463),
.B(n_98),
.C(n_100),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1368),
.A2(n_392),
.B(n_390),
.Y(n_1576)
);

O2A1O1Ixp5_ASAP7_75t_L g1577 ( 
.A1(n_1426),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1389),
.A2(n_105),
.B1(n_102),
.B2(n_103),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1437),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1355),
.B(n_103),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1424),
.A2(n_109),
.B(n_105),
.C(n_106),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1413),
.A2(n_111),
.B1(n_106),
.B2(n_110),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1331),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1416),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1346),
.B(n_562),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1422),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1435),
.A2(n_394),
.B(n_393),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1336),
.A2(n_397),
.B(n_396),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1400),
.A2(n_1491),
.B(n_1398),
.C(n_1459),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1405),
.B(n_113),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1388),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1433),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1452),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1391),
.B(n_116),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1334),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1466),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_SL g1597 ( 
.A1(n_1333),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_L g1598 ( 
.A(n_1481),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1322),
.A2(n_401),
.B(n_399),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1337),
.B(n_117),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1489),
.B(n_119),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1394),
.A2(n_123),
.B1(n_120),
.B2(n_121),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1422),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1444),
.A2(n_124),
.B(n_120),
.C(n_123),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1363),
.A2(n_404),
.B(n_402),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1363),
.A2(n_406),
.B(n_405),
.Y(n_1606)
);

AOI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1321),
.A2(n_408),
.B(n_407),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1456),
.A2(n_127),
.B(n_124),
.C(n_126),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1345),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1439),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1406),
.B(n_128),
.C(n_129),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1342),
.B(n_129),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1347),
.B(n_130),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1472),
.Y(n_1614)
);

O2A1O1Ixp33_ASAP7_75t_L g1615 ( 
.A1(n_1402),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1349),
.B(n_132),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1485),
.B(n_1483),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1360),
.B(n_133),
.Y(n_1618)
);

AO21x1_ASAP7_75t_L g1619 ( 
.A1(n_1447),
.A2(n_135),
.B(n_136),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1479),
.B(n_136),
.Y(n_1620)
);

A2O1A1Ixp33_ASAP7_75t_L g1621 ( 
.A1(n_1476),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1344),
.B(n_138),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1449),
.A2(n_410),
.B(n_409),
.Y(n_1623)
);

A2O1A1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1476),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1441),
.A2(n_413),
.B(n_412),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1374),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1353),
.B(n_141),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1481),
.Y(n_1628)
);

OAI21xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1454),
.A2(n_1465),
.B(n_1460),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1423),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1423),
.Y(n_1631)
);

CKINVDCx8_ASAP7_75t_R g1632 ( 
.A(n_1481),
.Y(n_1632)
);

OR2x6_ASAP7_75t_L g1633 ( 
.A(n_1448),
.B(n_142),
.Y(n_1633)
);

O2A1O1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1401),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1318),
.A2(n_415),
.B(n_414),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1490),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1412),
.B(n_560),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1423),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1477),
.B(n_147),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1411),
.A2(n_1492),
.B1(n_1429),
.B2(n_1431),
.Y(n_1640)
);

INVx4_ASAP7_75t_L g1641 ( 
.A(n_1477),
.Y(n_1641)
);

O2A1O1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1461),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1432),
.A2(n_154),
.B1(n_150),
.B2(n_152),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1477),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1462),
.A2(n_154),
.B(n_155),
.Y(n_1645)
);

NOR2xp67_ASAP7_75t_L g1646 ( 
.A(n_1442),
.B(n_417),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1482),
.A2(n_159),
.B(n_156),
.C(n_158),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1467),
.A2(n_158),
.B(n_160),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1362),
.A2(n_423),
.B(n_419),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1440),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1344),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1361),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1436),
.B(n_163),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1442),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1443),
.B(n_424),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1443),
.B(n_559),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1470),
.B(n_163),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1372),
.Y(n_1658)
);

INVx8_ASAP7_75t_L g1659 ( 
.A(n_1470),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1473),
.B(n_164),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1480),
.A2(n_1488),
.B(n_1487),
.C(n_1478),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1480),
.B(n_164),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1395),
.B(n_165),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1329),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1354),
.B(n_167),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1375),
.A2(n_426),
.B(n_425),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1378),
.Y(n_1667)
);

INVx4_ASAP7_75t_L g1668 ( 
.A(n_1384),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1396),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1451),
.A2(n_172),
.B1(n_169),
.B2(n_171),
.Y(n_1670)
);

O2A1O1Ixp5_ASAP7_75t_L g1671 ( 
.A1(n_1539),
.A2(n_1370),
.B(n_1430),
.C(n_1469),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1531),
.B(n_171),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1579),
.B(n_172),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1495),
.B(n_1486),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1607),
.A2(n_1377),
.B(n_1415),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1549),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1667),
.A2(n_1475),
.B(n_1419),
.Y(n_1677)
);

AO31x2_ASAP7_75t_L g1678 ( 
.A1(n_1669),
.A2(n_1468),
.A3(n_1471),
.B(n_1457),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1589),
.A2(n_433),
.B(n_431),
.Y(n_1679)
);

INVx3_ASAP7_75t_SL g1680 ( 
.A(n_1559),
.Y(n_1680)
);

AOI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1605),
.A2(n_173),
.B(n_174),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_L g1682 ( 
.A1(n_1499),
.A2(n_436),
.B(n_435),
.Y(n_1682)
);

AO31x2_ASAP7_75t_L g1683 ( 
.A1(n_1640),
.A2(n_438),
.A3(n_439),
.B(n_437),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1588),
.A2(n_441),
.B(n_440),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1606),
.A2(n_1572),
.B(n_1599),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1576),
.A2(n_1625),
.B(n_1535),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1566),
.B(n_174),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1567),
.A2(n_175),
.B(n_176),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1512),
.A2(n_443),
.B(n_442),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1497),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1504),
.B(n_177),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1520),
.A2(n_445),
.B(n_444),
.Y(n_1692)
);

NAND3x1_ASAP7_75t_L g1693 ( 
.A(n_1601),
.B(n_178),
.C(n_179),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1516),
.A2(n_178),
.B(n_179),
.Y(n_1694)
);

AO31x2_ASAP7_75t_L g1695 ( 
.A1(n_1661),
.A2(n_447),
.A3(n_448),
.B(n_446),
.Y(n_1695)
);

NOR2xp67_ASAP7_75t_L g1696 ( 
.A(n_1493),
.B(n_449),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1574),
.A2(n_454),
.B(n_450),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1650),
.A2(n_457),
.B(n_456),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1524),
.A2(n_463),
.B(n_458),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_SL g1700 ( 
.A(n_1633),
.B(n_464),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1583),
.B(n_180),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1497),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1501),
.B(n_180),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1507),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1500),
.A2(n_181),
.B(n_182),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1510),
.B(n_181),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1493),
.B(n_466),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1537),
.A2(n_468),
.B(n_467),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1626),
.A2(n_471),
.B(n_469),
.Y(n_1709)
);

O2A1O1Ixp5_ASAP7_75t_L g1710 ( 
.A1(n_1564),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1614),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_L g1712 ( 
.A1(n_1587),
.A2(n_1635),
.B(n_1498),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1493),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1623),
.A2(n_183),
.B(n_184),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1503),
.B(n_185),
.Y(n_1715)
);

A2O1A1Ixp33_ASAP7_75t_L g1716 ( 
.A1(n_1527),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1649),
.A2(n_473),
.B(n_472),
.Y(n_1717)
);

NOR4xp25_ASAP7_75t_L g1718 ( 
.A(n_1505),
.B(n_189),
.C(n_186),
.D(n_188),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1497),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1543),
.A2(n_188),
.B(n_189),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1546),
.A2(n_475),
.B(n_474),
.Y(n_1721)
);

AO31x2_ASAP7_75t_L g1722 ( 
.A1(n_1668),
.A2(n_558),
.A3(n_557),
.B(n_556),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1563),
.B(n_190),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1666),
.A2(n_478),
.B(n_477),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1536),
.A2(n_190),
.B(n_191),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1514),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1552),
.B(n_192),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1638),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1621),
.A2(n_193),
.B(n_194),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1629),
.A2(n_195),
.B(n_196),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1569),
.Y(n_1731)
);

NOR2xp67_ASAP7_75t_L g1732 ( 
.A(n_1496),
.B(n_479),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1509),
.B(n_195),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1655),
.A2(n_484),
.B(n_481),
.Y(n_1734)
);

BUFx10_ASAP7_75t_L g1735 ( 
.A(n_1517),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_SL g1736 ( 
.A1(n_1645),
.A2(n_197),
.B(n_198),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1541),
.A2(n_197),
.B(n_199),
.Y(n_1737)
);

OA21x2_ASAP7_75t_L g1738 ( 
.A1(n_1670),
.A2(n_487),
.B(n_485),
.Y(n_1738)
);

AO31x2_ASAP7_75t_L g1739 ( 
.A1(n_1668),
.A2(n_555),
.A3(n_553),
.B(n_552),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1550),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1617),
.A2(n_200),
.B(n_201),
.C(n_202),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1633),
.A2(n_1648),
.B(n_1663),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1624),
.A2(n_203),
.B(n_204),
.Y(n_1743)
);

AO31x2_ASAP7_75t_L g1744 ( 
.A1(n_1619),
.A2(n_551),
.A3(n_550),
.B(n_549),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1525),
.A2(n_204),
.B(n_205),
.Y(n_1745)
);

BUFx2_ASAP7_75t_SL g1746 ( 
.A(n_1496),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1519),
.A2(n_490),
.B(n_489),
.Y(n_1747)
);

OAI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1519),
.A2(n_492),
.B(n_491),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1533),
.B(n_205),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1591),
.B(n_206),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1510),
.B(n_206),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1525),
.A2(n_207),
.B(n_208),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1547),
.A2(n_496),
.B(n_495),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1594),
.A2(n_207),
.B(n_208),
.C(n_209),
.Y(n_1754)
);

AOI221x1_ASAP7_75t_L g1755 ( 
.A1(n_1575),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.C(n_212),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1551),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1611),
.A2(n_211),
.B(n_212),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1542),
.A2(n_498),
.B(n_497),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1558),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1502),
.B(n_213),
.Y(n_1760)
);

OAI21x1_ASAP7_75t_L g1761 ( 
.A1(n_1542),
.A2(n_500),
.B(n_499),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1532),
.B(n_213),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1570),
.B(n_214),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1538),
.A2(n_215),
.B(n_216),
.Y(n_1764)
);

AO31x2_ASAP7_75t_L g1765 ( 
.A1(n_1540),
.A2(n_548),
.A3(n_544),
.B(n_543),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1525),
.A2(n_215),
.B(n_217),
.Y(n_1766)
);

AO31x2_ASAP7_75t_L g1767 ( 
.A1(n_1523),
.A2(n_542),
.A3(n_541),
.B(n_539),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1622),
.B(n_218),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1596),
.B(n_220),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1530),
.A2(n_220),
.B(n_221),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1662),
.B(n_222),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1515),
.B(n_223),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1570),
.A2(n_538),
.B(n_534),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1620),
.B(n_223),
.Y(n_1774)
);

BUFx10_ASAP7_75t_L g1775 ( 
.A(n_1595),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1511),
.B(n_224),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1654),
.B(n_224),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1660),
.B(n_225),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1600),
.A2(n_226),
.B(n_227),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1586),
.B(n_229),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1496),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1628),
.B(n_230),
.Y(n_1782)
);

INVx4_ASAP7_75t_SL g1783 ( 
.A(n_1508),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1565),
.B(n_230),
.Y(n_1784)
);

INVx5_ASAP7_75t_L g1785 ( 
.A(n_1609),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1529),
.B(n_231),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1557),
.Y(n_1787)
);

A2O1A1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1665),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1609),
.B(n_232),
.Y(n_1789)
);

NOR2xp67_ASAP7_75t_L g1790 ( 
.A(n_1631),
.B(n_501),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1612),
.A2(n_233),
.B(n_235),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1573),
.B(n_235),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1494),
.B(n_236),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1598),
.B(n_238),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1561),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1598),
.B(n_239),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1592),
.Y(n_1797)
);

A2O1A1Ixp33_ASAP7_75t_L g1798 ( 
.A1(n_1590),
.A2(n_1627),
.B(n_1613),
.C(n_1616),
.Y(n_1798)
);

AO31x2_ASAP7_75t_L g1799 ( 
.A1(n_1560),
.A2(n_533),
.A3(n_531),
.B(n_530),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1571),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1545),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1577),
.A2(n_243),
.B(n_244),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1652),
.B(n_244),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1506),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1522),
.A2(n_527),
.B(n_526),
.Y(n_1806)
);

OAI21x1_ASAP7_75t_L g1807 ( 
.A1(n_1586),
.A2(n_525),
.B(n_523),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1618),
.B(n_245),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1632),
.Y(n_1809)
);

OAI21x1_ASAP7_75t_L g1810 ( 
.A1(n_1603),
.A2(n_522),
.B(n_519),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1580),
.Y(n_1811)
);

OAI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1642),
.A2(n_245),
.B(n_246),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1534),
.B(n_246),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1653),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1659),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1659),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1544),
.B(n_247),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1513),
.A2(n_249),
.B(n_250),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1647),
.A2(n_250),
.B(n_252),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1603),
.B(n_252),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1581),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.C(n_256),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1676),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1704),
.Y(n_1823)
);

OAI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1675),
.A2(n_1664),
.B(n_1584),
.Y(n_1824)
);

O2A1O1Ixp33_ASAP7_75t_SL g1825 ( 
.A1(n_1716),
.A2(n_1636),
.B(n_1556),
.C(n_1608),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1704),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1760),
.A2(n_1651),
.B1(n_1593),
.B2(n_1582),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1726),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1742),
.A2(n_1610),
.B1(n_1602),
.B2(n_1578),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1686),
.A2(n_1630),
.B(n_1644),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1781),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1787),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1671),
.A2(n_1528),
.B(n_1639),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1712),
.A2(n_1644),
.B(n_1630),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1728),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1685),
.A2(n_1646),
.B(n_1657),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1682),
.A2(n_1643),
.B(n_1615),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1803),
.B(n_1652),
.Y(n_1838)
);

CKINVDCx16_ASAP7_75t_R g1839 ( 
.A(n_1735),
.Y(n_1839)
);

AOI22x1_ASAP7_75t_L g1840 ( 
.A1(n_1812),
.A2(n_1562),
.B1(n_1652),
.B2(n_1641),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1705),
.A2(n_1521),
.B1(n_1637),
.B2(n_1518),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1730),
.A2(n_1634),
.B(n_1597),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1718),
.A2(n_1604),
.B1(n_1548),
.B2(n_1637),
.C(n_1555),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1805),
.A2(n_1656),
.B(n_1585),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_SL g1846 ( 
.A1(n_1688),
.A2(n_253),
.B(n_254),
.C(n_255),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1759),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1674),
.B(n_1526),
.Y(n_1848)
);

AND2x4_ASAP7_75t_L g1849 ( 
.A(n_1783),
.B(n_1526),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1725),
.A2(n_1819),
.B1(n_1694),
.B2(n_1727),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1811),
.B(n_1568),
.Y(n_1851)
);

OAI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1798),
.A2(n_1568),
.B(n_1658),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1681),
.A2(n_256),
.B(n_257),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1714),
.A2(n_258),
.B(n_259),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1757),
.A2(n_259),
.B(n_260),
.Y(n_1855)
);

O2A1O1Ixp33_ASAP7_75t_SL g1856 ( 
.A1(n_1788),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1797),
.Y(n_1857)
);

NAND2x1p5_ASAP7_75t_L g1858 ( 
.A(n_1809),
.B(n_502),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1806),
.A2(n_518),
.B(n_517),
.Y(n_1859)
);

OR2x6_ASAP7_75t_L g1860 ( 
.A(n_1674),
.B(n_504),
.Y(n_1860)
);

INVxp67_ASAP7_75t_SL g1861 ( 
.A(n_1677),
.Y(n_1861)
);

OR2x6_ASAP7_75t_L g1862 ( 
.A(n_1809),
.B(n_505),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1800),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1711),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1759),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1680),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_SL g1867 ( 
.A1(n_1789),
.A2(n_262),
.B(n_263),
.C(n_264),
.Y(n_1867)
);

INVx6_ASAP7_75t_L g1868 ( 
.A(n_1759),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1684),
.A2(n_516),
.B(n_515),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1700),
.A2(n_265),
.B(n_266),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1811),
.B(n_265),
.Y(n_1871)
);

OAI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1692),
.A2(n_514),
.B(n_510),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1677),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1805),
.A2(n_509),
.B(n_508),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1767),
.Y(n_1875)
);

AO21x2_ASAP7_75t_L g1876 ( 
.A1(n_1802),
.A2(n_507),
.B(n_267),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1762),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1767),
.Y(n_1878)
);

AO22x1_ASAP7_75t_L g1879 ( 
.A1(n_1764),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1695),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1749),
.Y(n_1881)
);

BUFx12f_ASAP7_75t_L g1882 ( 
.A(n_1735),
.Y(n_1882)
);

INVx2_ASAP7_75t_SL g1883 ( 
.A(n_1783),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1720),
.A2(n_268),
.B(n_269),
.Y(n_1884)
);

HB1xp67_ASAP7_75t_L g1885 ( 
.A(n_1695),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1771),
.B(n_1672),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1734),
.A2(n_269),
.B(n_270),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1754),
.B(n_270),
.C(n_271),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1750),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_L g1890 ( 
.A1(n_1708),
.A2(n_271),
.B(n_272),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1756),
.B(n_272),
.Y(n_1891)
);

OAI21x1_ASAP7_75t_L g1892 ( 
.A1(n_1699),
.A2(n_273),
.B(n_274),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1697),
.A2(n_273),
.B(n_274),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1741),
.A2(n_275),
.B(n_276),
.C(n_277),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1729),
.A2(n_275),
.B(n_279),
.Y(n_1895)
);

OAI21x1_ASAP7_75t_L g1896 ( 
.A1(n_1717),
.A2(n_1724),
.B(n_1721),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1781),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1747),
.A2(n_280),
.B(n_281),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1691),
.B(n_280),
.Y(n_1899)
);

OA21x2_ASAP7_75t_L g1900 ( 
.A1(n_1745),
.A2(n_281),
.B(n_282),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1770),
.A2(n_283),
.B(n_284),
.C(n_285),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1695),
.Y(n_1902)
);

OAI21x1_ASAP7_75t_L g1903 ( 
.A1(n_1748),
.A2(n_285),
.B(n_286),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1799),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1808),
.B(n_286),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1701),
.B(n_287),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1701),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1678),
.Y(n_1908)
);

CKINVDCx11_ASAP7_75t_R g1909 ( 
.A(n_1775),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1781),
.B(n_287),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1731),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_SL g1912 ( 
.A1(n_1700),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1758),
.A2(n_288),
.B(n_289),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1799),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1793),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1752),
.A2(n_290),
.B(n_291),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1822),
.B(n_1703),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1911),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1911),
.B(n_1713),
.Y(n_1919)
);

OA21x2_ASAP7_75t_L g1920 ( 
.A1(n_1861),
.A2(n_1766),
.B(n_1755),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1866),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1822),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1824),
.A2(n_1896),
.B(n_1836),
.Y(n_1923)
);

BUFx2_ASAP7_75t_SL g1924 ( 
.A(n_1866),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1823),
.B(n_1683),
.Y(n_1925)
);

OA21x2_ASAP7_75t_L g1926 ( 
.A1(n_1861),
.A2(n_1761),
.B(n_1773),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1880),
.A2(n_1689),
.B(n_1738),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1830),
.A2(n_1810),
.B(n_1807),
.Y(n_1928)
);

AOI21x1_ASAP7_75t_L g1929 ( 
.A1(n_1879),
.A2(n_1874),
.B(n_1900),
.Y(n_1929)
);

CKINVDCx8_ASAP7_75t_R g1930 ( 
.A(n_1839),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1880),
.A2(n_1689),
.B(n_1738),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1823),
.B(n_1683),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1826),
.Y(n_1933)
);

BUFx3_ASAP7_75t_L g1934 ( 
.A(n_1882),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1828),
.B(n_1683),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1850),
.A2(n_1693),
.B1(n_1740),
.B2(n_1814),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1832),
.B(n_1723),
.Y(n_1937)
);

AOI221xp5_ASAP7_75t_L g1938 ( 
.A1(n_1850),
.A2(n_1784),
.B1(n_1795),
.B2(n_1821),
.C(n_1673),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1838),
.B(n_1801),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1857),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1909),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1863),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1909),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1835),
.B(n_1813),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1848),
.B(n_1763),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1827),
.A2(n_1736),
.B1(n_1687),
.B2(n_1737),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1864),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1873),
.A2(n_1710),
.B(n_1779),
.Y(n_1948)
);

OA21x2_ASAP7_75t_L g1949 ( 
.A1(n_1873),
.A2(n_1791),
.B(n_1733),
.Y(n_1949)
);

NAND2x1_ASAP7_75t_L g1950 ( 
.A(n_1860),
.B(n_1780),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1881),
.B(n_1769),
.Y(n_1951)
);

AO21x2_ASAP7_75t_L g1952 ( 
.A1(n_1908),
.A2(n_1698),
.B(n_1709),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1885),
.A2(n_1679),
.B(n_1743),
.Y(n_1953)
);

OAI21x1_ASAP7_75t_L g1954 ( 
.A1(n_1834),
.A2(n_1818),
.B(n_1804),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1894),
.A2(n_1763),
.B(n_1753),
.Y(n_1955)
);

AO31x2_ASAP7_75t_L g1956 ( 
.A1(n_1875),
.A2(n_1715),
.A3(n_1772),
.B(n_1776),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1840),
.A2(n_1820),
.B(n_1786),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1882),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1908),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1885),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1902),
.A2(n_1778),
.B(n_1780),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1878),
.A2(n_1792),
.B(n_1777),
.Y(n_1962)
);

NAND2x1p5_ASAP7_75t_L g1963 ( 
.A(n_1849),
.B(n_1785),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1868),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1874),
.A2(n_1794),
.B(n_1796),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1940),
.B(n_1902),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1922),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1918),
.B(n_1886),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1922),
.B(n_1915),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1959),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1956),
.B(n_1877),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1923),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1933),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1926),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1959),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1925),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1919),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1917),
.B(n_1889),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1942),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1956),
.B(n_1886),
.Y(n_1980)
);

OR2x6_ASAP7_75t_L g1981 ( 
.A(n_1927),
.B(n_1848),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1960),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1960),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1925),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1947),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1919),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1918),
.B(n_1904),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1926),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1956),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1980),
.A2(n_1938),
.B1(n_1829),
.B2(n_1936),
.Y(n_1990)
);

AOI22xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1981),
.A2(n_1949),
.B1(n_1961),
.B2(n_1874),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1968),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1967),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1980),
.A2(n_1938),
.B1(n_1856),
.B2(n_1846),
.C(n_1901),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1981),
.A2(n_1955),
.B(n_1953),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1982),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1968),
.A2(n_1946),
.B1(n_1912),
.B2(n_1950),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1981),
.A2(n_1876),
.B1(n_1842),
.B2(n_1895),
.Y(n_1998)
);

INVx4_ASAP7_75t_L g1999 ( 
.A(n_1972),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1977),
.B(n_1944),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1974),
.Y(n_2001)
);

AOI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1981),
.A2(n_1876),
.B1(n_1842),
.B2(n_1962),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1981),
.A2(n_1962),
.B1(n_1884),
.B2(n_1888),
.Y(n_2003)
);

OAI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1981),
.A2(n_1961),
.B1(n_1848),
.B2(n_1860),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1967),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1977),
.Y(n_2006)
);

OAI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1981),
.A2(n_1860),
.B1(n_1953),
.B2(n_1929),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1966),
.Y(n_2008)
);

CKINVDCx6p67_ASAP7_75t_R g2009 ( 
.A(n_1969),
.Y(n_2009)
);

OAI211xp5_ASAP7_75t_L g2010 ( 
.A1(n_1982),
.A2(n_1912),
.B(n_1855),
.C(n_1844),
.Y(n_2010)
);

NOR4xp25_ASAP7_75t_L g2011 ( 
.A(n_1978),
.B(n_1951),
.C(n_1899),
.D(n_1846),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_2000),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_2000),
.Y(n_2013)
);

NAND3xp33_ASAP7_75t_L g2014 ( 
.A(n_1990),
.B(n_1901),
.C(n_1894),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_2008),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_2006),
.B(n_1977),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_2009),
.B(n_1986),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_2006),
.B(n_1986),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1992),
.B(n_1969),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_1996),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_SL g2021 ( 
.A1(n_2014),
.A2(n_1995),
.B1(n_1997),
.B2(n_2010),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_2017),
.B(n_2012),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_2019),
.B(n_2008),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_2020),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_2013),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2015),
.B(n_1993),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_2021),
.B(n_2011),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_2024),
.B(n_1941),
.Y(n_2028)
);

OAI31xp33_ASAP7_75t_L g2029 ( 
.A1(n_2025),
.A2(n_2014),
.A3(n_2007),
.B(n_1998),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_2026),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2022),
.B(n_2011),
.Y(n_2031)
);

AND2x2_ASAP7_75t_SL g2032 ( 
.A(n_2023),
.B(n_1994),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_SL g2033 ( 
.A1(n_2026),
.A2(n_1988),
.B1(n_1974),
.B2(n_1949),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_2024),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_2023),
.B(n_1969),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2030),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2028),
.B(n_2009),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2034),
.B(n_2016),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_2032),
.B(n_1905),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_2027),
.A2(n_1991),
.B1(n_2003),
.B2(n_2002),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2035),
.Y(n_2041)
);

AOI221x1_ASAP7_75t_L g2042 ( 
.A1(n_2031),
.A2(n_1971),
.B1(n_1870),
.B2(n_1999),
.C(n_1871),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2029),
.B(n_1993),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2033),
.B(n_2016),
.Y(n_2044)
);

NAND4xp25_ASAP7_75t_SL g2045 ( 
.A(n_2029),
.B(n_1706),
.C(n_1751),
.D(n_1930),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_L g2046 ( 
.A1(n_2027),
.A2(n_1774),
.B(n_1965),
.C(n_1906),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_2038),
.B(n_2037),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2038),
.B(n_1924),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_2036),
.B(n_1934),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_2039),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2041),
.B(n_2005),
.Y(n_2051)
);

INVxp67_ASAP7_75t_SL g2052 ( 
.A(n_2043),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_2046),
.B(n_2045),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2042),
.B(n_2005),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2051),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_2048),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2053),
.A2(n_2040),
.B1(n_2046),
.B2(n_2044),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2052),
.A2(n_2040),
.B1(n_2004),
.B2(n_1971),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2057),
.A2(n_2050),
.B1(n_2054),
.B2(n_2047),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2055),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2056),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2058),
.A2(n_2049),
.B1(n_1883),
.B2(n_1974),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2062),
.A2(n_2049),
.B1(n_1921),
.B2(n_1943),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2059),
.A2(n_1958),
.B(n_1867),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_2061),
.Y(n_2065)
);

O2A1O1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_2060),
.A2(n_1867),
.B(n_1856),
.C(n_1768),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2059),
.B(n_2001),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2065),
.Y(n_2068)
);

O2A1O1Ixp33_ASAP7_75t_L g2069 ( 
.A1(n_2064),
.A2(n_1817),
.B(n_1854),
.C(n_1862),
.Y(n_2069)
);

AOI21xp33_ASAP7_75t_SL g2070 ( 
.A1(n_2067),
.A2(n_1891),
.B(n_1775),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_2063),
.Y(n_2071)
);

O2A1O1Ixp33_ASAP7_75t_L g2072 ( 
.A1(n_2066),
.A2(n_1862),
.B(n_1853),
.C(n_1891),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_SL g2073 ( 
.A1(n_2067),
.A2(n_1816),
.B(n_2001),
.C(n_1983),
.Y(n_2073)
);

A2O1A1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_2064),
.A2(n_1988),
.B(n_1974),
.C(n_1843),
.Y(n_2074)
);

O2A1O1Ixp33_ASAP7_75t_SL g2075 ( 
.A1(n_2067),
.A2(n_1983),
.B(n_1785),
.C(n_1986),
.Y(n_2075)
);

NOR3xp33_ASAP7_75t_L g2076 ( 
.A(n_2065),
.B(n_1782),
.C(n_1707),
.Y(n_2076)
);

NOR3xp33_ASAP7_75t_L g2077 ( 
.A(n_2065),
.B(n_1732),
.C(n_1696),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_2077),
.A2(n_1988),
.B1(n_1974),
.B2(n_2018),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2068),
.B(n_1999),
.Y(n_2079)
);

O2A1O1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_2071),
.A2(n_1862),
.B(n_1825),
.C(n_1858),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2074),
.A2(n_1999),
.B1(n_2018),
.B2(n_1988),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2069),
.A2(n_1746),
.B1(n_1988),
.B2(n_1852),
.C(n_1937),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2076),
.A2(n_1849),
.B1(n_1910),
.B2(n_1838),
.Y(n_2083)
);

NAND3xp33_ASAP7_75t_SL g2084 ( 
.A(n_2072),
.B(n_1858),
.C(n_1963),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_2070),
.A2(n_1972),
.B1(n_1884),
.B2(n_1920),
.Y(n_2085)
);

OAI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_2073),
.A2(n_1785),
.B(n_1815),
.C(n_1970),
.Y(n_2086)
);

OAI32xp33_ASAP7_75t_L g2087 ( 
.A1(n_2075),
.A2(n_1841),
.A3(n_1978),
.B1(n_1963),
.B2(n_1972),
.Y(n_2087)
);

OAI211xp5_ASAP7_75t_L g2088 ( 
.A1(n_2068),
.A2(n_1970),
.B(n_1975),
.C(n_1972),
.Y(n_2088)
);

A2O1A1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_2069),
.A2(n_1957),
.B(n_1931),
.C(n_1972),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2068),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2090),
.B(n_1970),
.Y(n_2091)
);

INVx2_ASAP7_75t_SL g2092 ( 
.A(n_2079),
.Y(n_2092)
);

AOI221x1_ASAP7_75t_L g2093 ( 
.A1(n_2084),
.A2(n_1910),
.B1(n_1939),
.B2(n_1985),
.C(n_294),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2083),
.B(n_1978),
.Y(n_2094)
);

AOI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_2082),
.A2(n_1825),
.B1(n_1931),
.B2(n_1985),
.C(n_1979),
.Y(n_2095)
);

A2O1A1Ixp33_ASAP7_75t_SL g2096 ( 
.A1(n_2088),
.A2(n_291),
.B(n_292),
.C(n_293),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_2086),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2081),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2089),
.B(n_2080),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2078),
.B(n_1975),
.Y(n_2100)
);

AOI322xp5_ASAP7_75t_L g2101 ( 
.A1(n_2085),
.A2(n_1907),
.A3(n_1935),
.B1(n_1989),
.B2(n_1975),
.C1(n_1932),
.C2(n_1987),
.Y(n_2101)
);

AOI21xp33_ASAP7_75t_L g2102 ( 
.A1(n_2087),
.A2(n_1989),
.B(n_1884),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_2090),
.B(n_1719),
.Y(n_2103)
);

AOI311xp33_ASAP7_75t_L g2104 ( 
.A1(n_2096),
.A2(n_2099),
.A3(n_2098),
.B(n_2095),
.C(n_2092),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2091),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2097),
.A2(n_1900),
.B1(n_1916),
.B2(n_1868),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2093),
.Y(n_2107)
);

OAI21xp33_ASAP7_75t_L g2108 ( 
.A1(n_2103),
.A2(n_1841),
.B(n_1847),
.Y(n_2108)
);

OAI21xp33_ASAP7_75t_SL g2109 ( 
.A1(n_2100),
.A2(n_2101),
.B(n_2094),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_2102),
.A2(n_1916),
.B1(n_1900),
.B2(n_1868),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_L g2111 ( 
.A1(n_2099),
.A2(n_1979),
.B1(n_1973),
.B2(n_1935),
.C(n_1932),
.Y(n_2111)
);

OAI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_2096),
.A2(n_1916),
.B1(n_1865),
.B2(n_1719),
.C(n_1948),
.Y(n_2112)
);

XOR2x2_ASAP7_75t_L g2113 ( 
.A(n_2097),
.B(n_1790),
.Y(n_2113)
);

OAI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2098),
.A2(n_293),
.B(n_294),
.C(n_295),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_2091),
.Y(n_2115)
);

NOR2x1_ASAP7_75t_L g2116 ( 
.A(n_2105),
.B(n_296),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2107),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2114),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2115),
.Y(n_2119)
);

NOR2x1_ASAP7_75t_L g2120 ( 
.A(n_2104),
.B(n_2112),
.Y(n_2120)
);

NOR2x1_ASAP7_75t_L g2121 ( 
.A(n_2108),
.B(n_296),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2109),
.B(n_2113),
.Y(n_2122)
);

NOR2x1_ASAP7_75t_L g2123 ( 
.A(n_2110),
.B(n_297),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2111),
.B(n_1973),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2106),
.Y(n_2125)
);

OAI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2107),
.A2(n_1719),
.B1(n_1702),
.B2(n_1690),
.Y(n_2126)
);

NOR2x1_ASAP7_75t_L g2127 ( 
.A(n_2105),
.B(n_297),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2107),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2107),
.A2(n_1948),
.B1(n_1920),
.B2(n_1702),
.Y(n_2129)
);

NOR3xp33_ASAP7_75t_SL g2130 ( 
.A(n_2122),
.B(n_298),
.C(n_299),
.Y(n_2130)
);

INVxp33_ASAP7_75t_SL g2131 ( 
.A(n_2119),
.Y(n_2131)
);

NAND4xp75_ASAP7_75t_L g2132 ( 
.A(n_2120),
.B(n_298),
.C(n_299),
.D(n_300),
.Y(n_2132)
);

XNOR2xp5_ASAP7_75t_L g2133 ( 
.A(n_2116),
.B(n_300),
.Y(n_2133)
);

XNOR2xp5_ASAP7_75t_L g2134 ( 
.A(n_2127),
.B(n_301),
.Y(n_2134)
);

XOR2xp5_ASAP7_75t_L g2135 ( 
.A(n_2118),
.B(n_301),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2121),
.B(n_302),
.Y(n_2136)
);

NAND4xp75_ASAP7_75t_L g2137 ( 
.A(n_2117),
.B(n_303),
.C(n_304),
.D(n_305),
.Y(n_2137)
);

NAND2x1p5_ASAP7_75t_L g2138 ( 
.A(n_2128),
.B(n_2123),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2125),
.Y(n_2139)
);

XNOR2xp5_ASAP7_75t_L g2140 ( 
.A(n_2126),
.B(n_303),
.Y(n_2140)
);

NAND4xp75_ASAP7_75t_L g2141 ( 
.A(n_2124),
.B(n_304),
.C(n_306),
.D(n_307),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2129),
.Y(n_2142)
);

NOR2x1_ASAP7_75t_L g2143 ( 
.A(n_2119),
.B(n_307),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2116),
.Y(n_2144)
);

NAND2x1p5_ASAP7_75t_SL g2145 ( 
.A(n_2119),
.B(n_308),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2116),
.Y(n_2146)
);

AOI221xp5_ASAP7_75t_SL g2147 ( 
.A1(n_2119),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.C(n_311),
.Y(n_2147)
);

OAI31xp33_ASAP7_75t_L g2148 ( 
.A1(n_2138),
.A2(n_1690),
.A3(n_1831),
.B(n_1897),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2144),
.A2(n_1952),
.B1(n_1976),
.B2(n_1984),
.Y(n_2149)
);

OAI211xp5_ASAP7_75t_L g2150 ( 
.A1(n_2147),
.A2(n_312),
.B(n_313),
.C(n_314),
.Y(n_2150)
);

NOR2x1_ASAP7_75t_L g2151 ( 
.A(n_2132),
.B(n_312),
.Y(n_2151)
);

NAND3xp33_ASAP7_75t_SL g2152 ( 
.A(n_2146),
.B(n_314),
.C(n_315),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2143),
.A2(n_1872),
.B(n_1887),
.Y(n_2153)
);

AOI221x1_ASAP7_75t_L g2154 ( 
.A1(n_2145),
.A2(n_2139),
.B1(n_2136),
.B2(n_2142),
.C(n_2131),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2133),
.B(n_1744),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2135),
.A2(n_1833),
.B1(n_1831),
.B2(n_1897),
.Y(n_2156)
);

OAI221xp5_ASAP7_75t_L g2157 ( 
.A1(n_2134),
.A2(n_1833),
.B1(n_316),
.B2(n_317),
.C(n_318),
.Y(n_2157)
);

NAND4xp25_ASAP7_75t_L g2158 ( 
.A(n_2130),
.B(n_315),
.C(n_316),
.D(n_317),
.Y(n_2158)
);

CKINVDCx6p67_ASAP7_75t_R g2159 ( 
.A(n_2154),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_2151),
.B(n_2140),
.Y(n_2160)
);

XNOR2xp5_ASAP7_75t_L g2161 ( 
.A(n_2158),
.B(n_2137),
.Y(n_2161)
);

NAND3xp33_ASAP7_75t_L g2162 ( 
.A(n_2150),
.B(n_2141),
.C(n_319),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2155),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2153),
.B(n_318),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2152),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2157),
.A2(n_319),
.B(n_320),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2156),
.A2(n_1833),
.B1(n_1892),
.B2(n_1890),
.Y(n_2167)
);

XNOR2x1_ASAP7_75t_L g2168 ( 
.A(n_2148),
.B(n_320),
.Y(n_2168)
);

XNOR2xp5_ASAP7_75t_L g2169 ( 
.A(n_2149),
.B(n_321),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2151),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_2159),
.B(n_321),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2170),
.Y(n_2172)
);

OAI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_2165),
.A2(n_2162),
.B1(n_2168),
.B2(n_2161),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_2164),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2160),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2169),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2163),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2166),
.Y(n_2178)
);

XNOR2x1_ASAP7_75t_L g2179 ( 
.A(n_2167),
.B(n_322),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2159),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_2180),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2171),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2172),
.Y(n_2183)
);

AND2x2_ASAP7_75t_SL g2184 ( 
.A(n_2175),
.B(n_322),
.Y(n_2184)
);

AOI22x1_ASAP7_75t_L g2185 ( 
.A1(n_2177),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2174),
.Y(n_2186)
);

CKINVDCx20_ASAP7_75t_R g2187 ( 
.A(n_2173),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2178),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2179),
.Y(n_2189)
);

OR3x2_ASAP7_75t_L g2190 ( 
.A(n_2176),
.B(n_323),
.C(n_324),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_2183),
.A2(n_1893),
.B(n_1913),
.Y(n_2191)
);

AND2x2_ASAP7_75t_SL g2192 ( 
.A(n_2184),
.B(n_2188),
.Y(n_2192)
);

AO22x2_ASAP7_75t_L g2193 ( 
.A1(n_2182),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2181),
.B(n_327),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2187),
.A2(n_1964),
.B1(n_1851),
.B2(n_328),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2190),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2185),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2186),
.B(n_328),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2189),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2184),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2192),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_2200),
.B(n_2199),
.Y(n_2202)
);

INVxp33_ASAP7_75t_L g2203 ( 
.A(n_2196),
.Y(n_2203)
);

XNOR2xp5_ASAP7_75t_L g2204 ( 
.A(n_2194),
.B(n_329),
.Y(n_2204)
);

AOI21xp33_ASAP7_75t_L g2205 ( 
.A1(n_2197),
.A2(n_1903),
.B(n_1898),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2198),
.Y(n_2206)
);

AO22x2_ASAP7_75t_L g2207 ( 
.A1(n_2195),
.A2(n_1945),
.B1(n_1987),
.B2(n_1966),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2193),
.Y(n_2208)
);

AOI22x1_ASAP7_75t_L g2209 ( 
.A1(n_2202),
.A2(n_2191),
.B1(n_1945),
.B2(n_1739),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2201),
.A2(n_1869),
.B1(n_1837),
.B2(n_1954),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_2203),
.A2(n_1966),
.B1(n_1859),
.B2(n_1987),
.Y(n_2211)
);

NAND3xp33_ASAP7_75t_L g2212 ( 
.A(n_2208),
.B(n_1722),
.C(n_1739),
.Y(n_2212)
);

AOI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2206),
.A2(n_1845),
.B1(n_1984),
.B2(n_1976),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2212),
.A2(n_2204),
.B1(n_2207),
.B2(n_2205),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_2214),
.A2(n_2209),
.B1(n_2213),
.B2(n_2211),
.Y(n_2215)
);

AOI22xp5_ASAP7_75t_SL g2216 ( 
.A1(n_2215),
.A2(n_2210),
.B1(n_1722),
.B2(n_1739),
.Y(n_2216)
);

AOI22xp5_ASAP7_75t_SL g2217 ( 
.A1(n_2215),
.A2(n_1722),
.B1(n_1765),
.B2(n_1744),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2216),
.B(n_1765),
.Y(n_2218)
);

AOI221xp5_ASAP7_75t_L g2219 ( 
.A1(n_2218),
.A2(n_2217),
.B1(n_1765),
.B2(n_1845),
.C(n_1984),
.Y(n_2219)
);

AOI211xp5_ASAP7_75t_L g2220 ( 
.A1(n_2219),
.A2(n_1744),
.B(n_1928),
.C(n_1914),
.Y(n_2220)
);


endmodule