module fake_ibex_1672_n_3532 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3532);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3532;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3411;
wire n_3025;
wire n_2955;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_667;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2436;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_3030;
wire n_3097;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3510;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_660;
wire n_2590;
wire n_3119;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_3034;
wire n_2612;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2979;
wire n_2376;
wire n_3398;
wire n_2476;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2654;
wire n_2463;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_991;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2437;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_648;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_1455;
wire n_804;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2816;
wire n_2803;
wire n_2433;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_3236;
wire n_2658;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_946;
wire n_1362;
wire n_707;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_3173;
wire n_3102;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_750;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_3223;
wire n_3318;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_1532;
wire n_791;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_3067;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_2928;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3286;
wire n_3124;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2148;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2302;
wire n_2453;
wire n_2082;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_2168;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_1383;
wire n_990;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2970;
wire n_1393;
wire n_2497;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

INVx1_ASAP7_75t_L g646 ( 
.A(n_91),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_270),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_205),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_415),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_24),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_570),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_366),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_305),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_404),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_199),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_35),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_637),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_272),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_216),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_536),
.Y(n_660)
);

INVxp33_ASAP7_75t_SL g661 ( 
.A(n_15),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_542),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_413),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_622),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_463),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_412),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_174),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_46),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_102),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_499),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_23),
.Y(n_671)
);

BUFx2_ASAP7_75t_L g672 ( 
.A(n_638),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_538),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_294),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_619),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_229),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_94),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_284),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_56),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_95),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_541),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_614),
.Y(n_682)
);

CKINVDCx14_ASAP7_75t_R g683 ( 
.A(n_539),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_237),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_264),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_464),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_157),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_32),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_242),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_254),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_271),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_423),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_302),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_73),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_253),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_321),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_117),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_386),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_559),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_366),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_80),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_17),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_53),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_380),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_531),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_340),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_453),
.Y(n_707)
);

CKINVDCx16_ASAP7_75t_R g708 ( 
.A(n_510),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_644),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_150),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_424),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_552),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_293),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_409),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_357),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_399),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_448),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_377),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_16),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_588),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_523),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_387),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_485),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_550),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_428),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_108),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_219),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_440),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_458),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_159),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_595),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_428),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_551),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_470),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_447),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_92),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_563),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_199),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_106),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_346),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_181),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_45),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_504),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_341),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_345),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_407),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_601),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_599),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_367),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_123),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_358),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_609),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_573),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_560),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_537),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_554),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_130),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_124),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_628),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_239),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_109),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_488),
.B(n_313),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_602),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_179),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_70),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_312),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_200),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_60),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_639),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_4),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_632),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_45),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_99),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_534),
.Y(n_774)
);

BUFx2_ASAP7_75t_L g775 ( 
.A(n_39),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_295),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_338),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_482),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_310),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_275),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_196),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_634),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_413),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_163),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_430),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_327),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_252),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_371),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_37),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_498),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_56),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_438),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_154),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_321),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_152),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_326),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_51),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_507),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_403),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_623),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_320),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_226),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_640),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_481),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_433),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_348),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_515),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_101),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_270),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_641),
.Y(n_810)
);

CKINVDCx20_ASAP7_75t_R g811 ( 
.A(n_285),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_613),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_245),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_52),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_331),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_597),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_589),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_66),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_630),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_64),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_286),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_216),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_211),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_467),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_439),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_492),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_576),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_491),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_156),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_506),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_299),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_273),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_535),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_482),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_310),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_346),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_624),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_5),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_243),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_402),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_512),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_95),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_128),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_567),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_188),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_34),
.Y(n_847)
);

CKINVDCx14_ASAP7_75t_R g848 ( 
.A(n_92),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_618),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_400),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_373),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_610),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_549),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_60),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_49),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_370),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_416),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_203),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_168),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_458),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_493),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_304),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_74),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_103),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_131),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_471),
.Y(n_866)
);

INVxp33_ASAP7_75t_SL g867 ( 
.A(n_49),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_139),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_594),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_530),
.Y(n_870)
);

BUFx2_ASAP7_75t_SL g871 ( 
.A(n_396),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_385),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_509),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_511),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_489),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_26),
.Y(n_876)
);

CKINVDCx14_ASAP7_75t_R g877 ( 
.A(n_5),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_212),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_438),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_625),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_344),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_411),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_26),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_607),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_506),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_631),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_591),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_388),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_345),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_88),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_34),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_156),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_626),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_352),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_67),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_575),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_141),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_546),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_642),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_437),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_574),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_309),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_324),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_249),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_23),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_127),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_40),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_93),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_158),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_612),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_267),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_357),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_633),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_616),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_518),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_508),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_103),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_627),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_209),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_308),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_572),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_365),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_582),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_281),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_261),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_435),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_37),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_350),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_69),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_600),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_360),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_128),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_11),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_358),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_30),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_556),
.Y(n_936)
);

CKINVDCx16_ASAP7_75t_R g937 ( 
.A(n_440),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_488),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_492),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_220),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_264),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_226),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_433),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_120),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_302),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_35),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_90),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_503),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_317),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_192),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_273),
.Y(n_951)
);

BUFx2_ASAP7_75t_SL g952 ( 
.A(n_568),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_261),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_571),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_596),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_334),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_584),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_215),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_185),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_395),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_101),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_405),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_225),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_10),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_343),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_306),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_432),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_27),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_444),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_636),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_517),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_324),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_145),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_195),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_402),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_374),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_643),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_645),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_540),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_254),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_255),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_2),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_134),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_33),
.B(n_381),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_376),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_418),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_335),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_224),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_519),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_404),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_331),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_248),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_330),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_369),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_514),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_548),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_278),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_73),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_292),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_617),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_494),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_301),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_598),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_308),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_102),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_339),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_123),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_407),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_64),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_629),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_501),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_502),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_253),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_46),
.B(n_285),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_390),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_191),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_483),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_280),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_496),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_392),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_370),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_309),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_452),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_347),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_185),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_389),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_327),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_495),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_593),
.Y(n_1029)
);

NOR2xp67_ASAP7_75t_L g1030 ( 
.A(n_62),
.B(n_141),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_365),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_377),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_909),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_739),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_697),
.B(n_765),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_686),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_739),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_739),
.Y(n_1038)
);

INVxp33_ASAP7_75t_L g1039 ( 
.A(n_711),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_763),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_763),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_775),
.B(n_799),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_816),
.B(n_1),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_909),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_763),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_763),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_739),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_848),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_649),
.A2(n_4),
.B1(n_0),
.B2(n_3),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_842),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_739),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_739),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_731),
.A2(n_516),
.B(n_513),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_739),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_870),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_842),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_870),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_870),
.Y(n_1058)
);

BUFx12f_ASAP7_75t_L g1059 ( 
.A(n_714),
.Y(n_1059)
);

BUFx12f_ASAP7_75t_L g1060 ( 
.A(n_714),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_870),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_995),
.B(n_3),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_719),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_655),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_720),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_877),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_720),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_714),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_662),
.B(n_520),
.Y(n_1069)
);

BUFx8_ASAP7_75t_SL g1070 ( 
.A(n_649),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_738),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_691),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_738),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_655),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_720),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_655),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_655),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_674),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_674),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_689),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_689),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_665),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_703),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_691),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_659),
.A2(n_13),
.B1(n_9),
.B2(n_12),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_796),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_722),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_749),
.Y(n_1088)
);

INVx3_ASAP7_75t_L g1089 ( 
.A(n_722),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_703),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_749),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_SL g1092 ( 
.A(n_681),
.B(n_521),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_705),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_732),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_749),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_825),
.B(n_14),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_732),
.Y(n_1097)
);

AND2x2_ASAP7_75t_SL g1098 ( 
.A(n_810),
.B(n_13),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_865),
.B(n_15),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_783),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_884),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_741),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_R g1103 ( 
.A1(n_659),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_1103)
);

AND2x4_ASAP7_75t_L g1104 ( 
.A(n_796),
.B(n_18),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_783),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_749),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_884),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_908),
.B(n_19),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_731),
.A2(n_524),
.B(n_522),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_884),
.Y(n_1110)
);

BUFx8_ASAP7_75t_SL g1111 ( 
.A(n_718),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_784),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_784),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_938),
.B(n_19),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_995),
.B(n_18),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_772),
.Y(n_1116)
);

BUFx8_ASAP7_75t_SL g1117 ( 
.A(n_718),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_772),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_772),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_846),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_850),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_740),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_850),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_955),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_772),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_959),
.B(n_20),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_833),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_955),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_833),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1009),
.B(n_22),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_781),
.B(n_24),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_708),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_821),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_846),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_735),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1104),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1036),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1104),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1126),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1070),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1126),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1111),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1086),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1121),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1110),
.B(n_672),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1117),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1123),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1089),
.Y(n_1148)
);

CKINVDCx16_ASAP7_75t_R g1149 ( 
.A(n_1082),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_1059),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1060),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1093),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1132),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1110),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1065),
.B(n_914),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1063),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1120),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1065),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1039),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1040),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1102),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1133),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1067),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1101),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1050),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1033),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1103),
.Y(n_1167)
);

INVxp33_ASAP7_75t_SL g1168 ( 
.A(n_1035),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1033),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1120),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1128),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_R g1172 ( 
.A(n_1068),
.B(n_683),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1072),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1042),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1044),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1075),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_L g1177 ( 
.A(n_1075),
.B(n_1107),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1075),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_1124),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1084),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1056),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1107),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_L g1183 ( 
.A(n_1107),
.B(n_862),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1087),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1034),
.A2(n_813),
.B(n_733),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_1085),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_R g1187 ( 
.A(n_1068),
.B(n_747),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1100),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1098),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1056),
.Y(n_1190)
);

XOR2xp5_ASAP7_75t_L g1191 ( 
.A(n_1049),
.B(n_747),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1122),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1105),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1112),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1048),
.Y(n_1195)
);

BUFx10_ASAP7_75t_L g1196 ( 
.A(n_1062),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1113),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1134),
.Y(n_1198)
);

NOR2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1131),
.B(n_677),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1037),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1066),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1043),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1071),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1096),
.Y(n_1204)
);

HB1xp67_ASAP7_75t_L g1205 ( 
.A(n_1099),
.Y(n_1205)
);

NOR2xp67_ASAP7_75t_L g1206 ( 
.A(n_1078),
.B(n_924),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1040),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1108),
.Y(n_1208)
);

CKINVDCx16_ASAP7_75t_R g1209 ( 
.A(n_1092),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1114),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1130),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1078),
.B(n_874),
.Y(n_1212)
);

AND3x2_ASAP7_75t_L g1213 ( 
.A(n_1115),
.B(n_767),
.C(n_761),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1073),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1079),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1038),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1079),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1080),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1069),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1080),
.B(n_959),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_L g1221 ( 
.A(n_1081),
.B(n_1018),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1081),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1047),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1051),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_R g1225 ( 
.A(n_1083),
.B(n_748),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1083),
.Y(n_1226)
);

AND3x2_ASAP7_75t_L g1227 ( 
.A(n_1090),
.B(n_676),
.C(n_670),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1090),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1094),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1052),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1097),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1054),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1097),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_1135),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1135),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1057),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1057),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1057),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1064),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1053),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1064),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1053),
.A2(n_867),
.B1(n_661),
.B2(n_937),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1109),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1064),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1074),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1109),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1074),
.Y(n_1247)
);

NOR2x1p5_ASAP7_75t_L g1248 ( 
.A(n_1076),
.B(n_677),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1076),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1077),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1077),
.B(n_970),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1077),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1088),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1088),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_SL g1255 ( 
.A1(n_1088),
.A2(n_740),
.B1(n_790),
.B2(n_786),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1091),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1091),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1091),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1095),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_R g1260 ( 
.A(n_1095),
.B(n_748),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1095),
.Y(n_1261)
);

BUFx10_ASAP7_75t_L g1262 ( 
.A(n_1106),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1106),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1106),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1129),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1040),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1116),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_1116),
.B(n_1018),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1116),
.B(n_733),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1118),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1118),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1118),
.B(n_939),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1119),
.B(n_813),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1119),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1119),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1125),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1125),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1127),
.B(n_955),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1129),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1129),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1041),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1041),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1041),
.Y(n_1283)
);

CKINVDCx16_ASAP7_75t_R g1284 ( 
.A(n_1045),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1045),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1045),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1046),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1046),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1046),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1055),
.Y(n_1290)
);

NAND2xp33_ASAP7_75t_R g1291 ( 
.A(n_1055),
.B(n_661),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_R g1292 ( 
.A(n_1055),
.B(n_828),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_R g1293 ( 
.A(n_1058),
.B(n_913),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_1058),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1058),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1061),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1061),
.B(n_913),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1082),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1070),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1070),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1070),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1070),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1070),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_R g1304 ( 
.A(n_1093),
.B(n_918),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1070),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1070),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_R g1307 ( 
.A(n_1093),
.B(n_918),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1070),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1089),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_R g1310 ( 
.A(n_1093),
.B(n_994),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1104),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1070),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1070),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1070),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1070),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1082),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1104),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1082),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1104),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1070),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_R g1321 ( 
.A(n_1093),
.B(n_771),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1211),
.B(n_771),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_SL g1323 ( 
.A(n_1179),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1159),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1288),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1231),
.B(n_1000),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1137),
.B(n_692),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1143),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_1137),
.Y(n_1329)
);

BUFx8_ASAP7_75t_L g1330 ( 
.A(n_1150),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1144),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1151),
.B(n_871),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1147),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1170),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1168),
.B(n_1003),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1199),
.B(n_1021),
.Y(n_1336)
);

NAND2xp33_ASAP7_75t_L g1337 ( 
.A(n_1172),
.B(n_1243),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1205),
.B(n_1145),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1196),
.B(n_1010),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1156),
.B(n_692),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1220),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1202),
.B(n_660),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1145),
.B(n_867),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1240),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1138),
.B(n_529),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1156),
.B(n_685),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1246),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1215),
.B(n_664),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1173),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1180),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1220),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1204),
.B(n_675),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1162),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1138),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1218),
.B(n_699),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_1208),
.B(n_709),
.Y(n_1356)
);

NOR3xp33_ASAP7_75t_L g1357 ( 
.A(n_1255),
.B(n_1032),
.C(n_905),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1210),
.B(n_712),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1185),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1226),
.B(n_721),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1161),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1228),
.B(n_1229),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1184),
.Y(n_1363)
);

AO221x1_ASAP7_75t_L g1364 ( 
.A1(n_1189),
.A2(n_794),
.B1(n_811),
.B2(n_790),
.C(n_786),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1304),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1161),
.B(n_1183),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1148),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1136),
.B(n_1139),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1174),
.B(n_684),
.C(n_678),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1141),
.A2(n_892),
.B(n_958),
.C(n_851),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1234),
.A2(n_811),
.B1(n_814),
.B2(n_794),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1233),
.B(n_724),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1235),
.B(n_737),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1179),
.B(n_651),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1188),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1194),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1309),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1262),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1321),
.B(n_999),
.Y(n_1379)
);

OR2x6_ASAP7_75t_L g1380 ( 
.A(n_1206),
.B(n_1248),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1190),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1166),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1155),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1311),
.B(n_752),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1317),
.B(n_755),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1217),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1149),
.B(n_1192),
.C(n_1209),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1319),
.B(n_756),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1291),
.B(n_684),
.C(n_678),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1221),
.Y(n_1390)
);

INVxp33_ASAP7_75t_L g1391 ( 
.A(n_1225),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1175),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1163),
.B(n_759),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1193),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1157),
.B(n_769),
.Y(n_1395)
);

NOR3xp33_ASAP7_75t_L g1396 ( 
.A(n_1195),
.B(n_701),
.C(n_696),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1272),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1219),
.B(n_774),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1197),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1198),
.Y(n_1400)
);

BUFx5_ASAP7_75t_L g1401 ( 
.A(n_1224),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1155),
.B(n_1212),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1165),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1181),
.B(n_800),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_SL g1405 ( 
.A(n_1158),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1164),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1291),
.B(n_687),
.C(n_685),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1283),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1181),
.B(n_803),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1284),
.B(n_812),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1176),
.B(n_817),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1178),
.B(n_834),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1182),
.B(n_978),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1269),
.B(n_532),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1177),
.B(n_845),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1213),
.B(n_849),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1269),
.B(n_1273),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1213),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1222),
.B(n_695),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1243),
.B(n_1232),
.C(n_1223),
.Y(n_1421)
);

NAND2xp33_ASAP7_75t_L g1422 ( 
.A(n_1292),
.B(n_880),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1278),
.B(n_886),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1227),
.B(n_898),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1251),
.B(n_1200),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1247),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1247),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1294),
.B(n_899),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1227),
.B(n_901),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1152),
.B(n_910),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1257),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1276),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1276),
.Y(n_1433)
);

NOR3xp33_ASAP7_75t_L g1434 ( 
.A(n_1201),
.B(n_727),
.C(n_713),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1171),
.B(n_1298),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1216),
.B(n_1230),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1237),
.B(n_915),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1268),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1187),
.B(n_923),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1292),
.B(n_930),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1214),
.B(n_936),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1262),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1239),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1293),
.B(n_1260),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1203),
.B(n_1153),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1273),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1236),
.B(n_957),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1304),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1287),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1238),
.B(n_971),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1277),
.B(n_1014),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1297),
.B(n_977),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1310),
.B(n_979),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1280),
.Y(n_1455)
);

AO221x1_ASAP7_75t_L g1456 ( 
.A1(n_1307),
.A2(n_872),
.B1(n_883),
.B2(n_826),
.C(n_814),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1241),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1310),
.B(n_989),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1244),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1290),
.Y(n_1460)
);

BUFx5_ASAP7_75t_L g1461 ( 
.A(n_1281),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1245),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1252),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1295),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1191),
.B(n_695),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1256),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_L g1467 ( 
.A(n_1263),
.B(n_1029),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1267),
.B(n_657),
.Y(n_1468)
);

INVxp33_ASAP7_75t_L g1469 ( 
.A(n_1140),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1270),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1271),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1142),
.B(n_687),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1146),
.B(n_688),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1274),
.B(n_688),
.Y(n_1474)
);

NAND2xp33_ASAP7_75t_L g1475 ( 
.A(n_1275),
.B(n_852),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1259),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1254),
.B(n_693),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1254),
.B(n_693),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1253),
.B(n_997),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1258),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1261),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1299),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1264),
.A2(n_892),
.B(n_958),
.C(n_851),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1160),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1186),
.B(n_952),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1282),
.B(n_999),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1285),
.B(n_1001),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1167),
.B(n_673),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1249),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1300),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1301),
.B(n_682),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1250),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1289),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1279),
.B(n_1001),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1286),
.B(n_1004),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1160),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1296),
.B(n_1004),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1302),
.B(n_753),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1207),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1207),
.B(n_754),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1266),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1266),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1303),
.B(n_1008),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1305),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1306),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1320),
.Y(n_1506)
);

BUFx5_ASAP7_75t_L g1507 ( 
.A(n_1308),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1312),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1313),
.B(n_1008),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1314),
.B(n_1011),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1315),
.B(n_1011),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1169),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1159),
.B(n_648),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1211),
.B(n_650),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1211),
.B(n_652),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1159),
.B(n_653),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1168),
.B(n_782),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1169),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1169),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1169),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1168),
.B(n_807),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1211),
.B(n_658),
.Y(n_1522)
);

INVxp33_ASAP7_75t_L g1523 ( 
.A(n_1137),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1211),
.B(n_663),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1211),
.B(n_666),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_SL g1526 ( 
.A(n_1159),
.B(n_818),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1159),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1159),
.B(n_773),
.Y(n_1528)
);

NOR3xp33_ASAP7_75t_L g1529 ( 
.A(n_1255),
.B(n_1015),
.C(n_894),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1159),
.B(n_820),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1240),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1173),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_L g1533 ( 
.A(n_1242),
.B(n_668),
.C(n_667),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1136),
.A2(n_647),
.B1(n_654),
.B2(n_646),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1159),
.B(n_838),
.Y(n_1535)
);

INVxp33_ASAP7_75t_L g1536 ( 
.A(n_1137),
.Y(n_1536)
);

INVx4_ASAP7_75t_L g1537 ( 
.A(n_1284),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1159),
.Y(n_1538)
);

NOR2xp67_ASAP7_75t_L g1539 ( 
.A(n_1242),
.B(n_533),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1169),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1159),
.B(n_853),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1150),
.B(n_762),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1169),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1173),
.Y(n_1544)
);

INVx8_ASAP7_75t_L g1545 ( 
.A(n_1154),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1159),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1284),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1211),
.B(n_669),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1159),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1211),
.B(n_671),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1240),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1136),
.A2(n_679),
.B1(n_680),
.B2(n_656),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1173),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1211),
.B(n_698),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1168),
.B(n_869),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1211),
.B(n_702),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_SL g1557 ( 
.A(n_1179),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1159),
.B(n_706),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1173),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1168),
.B(n_887),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1211),
.B(n_710),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1173),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1159),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1211),
.B(n_716),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1159),
.B(n_1022),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1159),
.B(n_893),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1159),
.B(n_717),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1211),
.B(n_723),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1173),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1527),
.B(n_872),
.C(n_826),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1338),
.B(n_725),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1030),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1354),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1361),
.A2(n_904),
.B1(n_907),
.B2(n_883),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1563),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1341),
.Y(n_1577)
);

NOR3xp33_ASAP7_75t_SL g1578 ( 
.A(n_1371),
.B(n_728),
.C(n_726),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1351),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1328),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1329),
.A2(n_907),
.B1(n_928),
.B2(n_904),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1403),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1344),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1331),
.Y(n_1584)
);

A2O1A1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1333),
.A2(n_694),
.B(n_700),
.C(n_690),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1370),
.A2(n_1402),
.B(n_1357),
.C(n_1529),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1538),
.B(n_928),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1335),
.B(n_1322),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1330),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1523),
.B(n_929),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1536),
.A2(n_736),
.B1(n_743),
.B2(n_730),
.Y(n_1591)
);

NOR2x2_ASAP7_75t_L g1592 ( 
.A(n_1542),
.B(n_929),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1378),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1392),
.Y(n_1594)
);

AND2x6_ASAP7_75t_L g1595 ( 
.A(n_1344),
.B(n_996),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1343),
.A2(n_751),
.B1(n_757),
.B2(n_750),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1517),
.B(n_758),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1546),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1334),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1545),
.B(n_735),
.Y(n_1600)
);

NOR2xp67_ASAP7_75t_L g1601 ( 
.A(n_1324),
.B(n_1549),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1521),
.A2(n_766),
.B1(n_770),
.B2(n_760),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1399),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1400),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_SL g1605 ( 
.A(n_1365),
.B(n_1017),
.C(n_940),
.Y(n_1605)
);

BUFx4f_ASAP7_75t_L g1606 ( 
.A(n_1545),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1382),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1378),
.Y(n_1608)
);

BUFx4f_ASAP7_75t_L g1609 ( 
.A(n_1545),
.Y(n_1609)
);

INVx3_ASAP7_75t_SL g1610 ( 
.A(n_1547),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1394),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1401),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1555),
.B(n_776),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1367),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_R g1615 ( 
.A(n_1449),
.B(n_933),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1560),
.B(n_777),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1377),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1327),
.B(n_933),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1330),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1533),
.A2(n_944),
.B1(n_964),
.B2(n_940),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1353),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1386),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1537),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1537),
.B(n_704),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1514),
.B(n_778),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1362),
.B(n_944),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1368),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1378),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1381),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1515),
.B(n_1554),
.Y(n_1630)
);

NAND2xp33_ASAP7_75t_L g1631 ( 
.A(n_1344),
.B(n_779),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1325),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1438),
.B(n_787),
.C(n_785),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1522),
.B(n_788),
.Y(n_1634)
);

INVx6_ASAP7_75t_L g1635 ( 
.A(n_1332),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1426),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1524),
.B(n_789),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1349),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1340),
.B(n_964),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1346),
.B(n_1379),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1525),
.B(n_1568),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1350),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1548),
.B(n_797),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1363),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1375),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1397),
.B(n_976),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1376),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1396),
.A2(n_715),
.B(n_729),
.C(n_707),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1550),
.B(n_798),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1418),
.A2(n_805),
.B1(n_809),
.B2(n_801),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1427),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1556),
.B(n_1561),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1421),
.A2(n_921),
.B(n_896),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1332),
.B(n_1542),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1532),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1336),
.B(n_734),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1544),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1553),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_R g1659 ( 
.A(n_1323),
.B(n_976),
.Y(n_1659)
);

NOR2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1431),
.B(n_991),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1559),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1528),
.A2(n_998),
.B1(n_991),
.B2(n_1017),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1558),
.B(n_998),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1432),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1562),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1336),
.B(n_742),
.Y(n_1666)
);

INVx6_ASAP7_75t_L g1667 ( 
.A(n_1507),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1482),
.B(n_1027),
.C(n_824),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1565),
.B(n_822),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1465),
.A2(n_831),
.B(n_835),
.C(n_827),
.Y(n_1670)
);

BUFx8_ASAP7_75t_L g1671 ( 
.A(n_1323),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1569),
.Y(n_1672)
);

AND2x6_ASAP7_75t_L g1673 ( 
.A(n_1347),
.B(n_996),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1564),
.B(n_1326),
.Y(n_1674)
);

INVx3_ASAP7_75t_SL g1675 ( 
.A(n_1504),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1490),
.Y(n_1676)
);

AND2x4_ASAP7_75t_SL g1677 ( 
.A(n_1513),
.B(n_744),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1408),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1420),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1383),
.B(n_1369),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_SL g1681 ( 
.A(n_1435),
.B(n_840),
.C(n_839),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1433),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1534),
.B(n_843),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_L g1684 ( 
.A(n_1434),
.B(n_858),
.C(n_847),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1516),
.B(n_860),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1442),
.A2(n_866),
.B1(n_873),
.B2(n_864),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1552),
.A2(n_745),
.B1(n_764),
.B2(n_746),
.Y(n_1687)
);

BUFx4f_ASAP7_75t_L g1688 ( 
.A(n_1505),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1567),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1347),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1457),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1390),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1539),
.B(n_876),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1348),
.B(n_881),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1494),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1436),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1495),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1512),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1497),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1355),
.B(n_882),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1419),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1447),
.A2(n_768),
.B1(n_793),
.B2(n_780),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1531),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1360),
.B(n_888),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1531),
.B(n_889),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_SL g1706 ( 
.A(n_1488),
.B(n_897),
.C(n_895),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1557),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1518),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1519),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1457),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1389),
.A2(n_911),
.B1(n_912),
.B2(n_906),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1551),
.B(n_916),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1457),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1406),
.B(n_922),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1462),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1477),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_SL g1717 ( 
.A1(n_1453),
.A2(n_984),
.B(n_954),
.C(n_791),
.Y(n_1717)
);

BUFx3_ASAP7_75t_L g1718 ( 
.A(n_1462),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1407),
.B(n_1503),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1478),
.Y(n_1720)
);

INVx5_ASAP7_75t_L g1721 ( 
.A(n_1466),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1455),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1466),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1443),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1557),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1520),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1446),
.A2(n_934),
.B1(n_935),
.B2(n_927),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1380),
.B(n_795),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1466),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1372),
.B(n_942),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1540),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1373),
.B(n_945),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1428),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1366),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1543),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_1508),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1444),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1339),
.B(n_947),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1380),
.B(n_802),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1444),
.Y(n_1740)
);

INVx5_ASAP7_75t_L g1741 ( 
.A(n_1366),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1384),
.B(n_1374),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1472),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1425),
.B(n_953),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1473),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1359),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1364),
.A2(n_806),
.B1(n_808),
.B2(n_804),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1479),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1509),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_SL g1750 ( 
.A(n_1506),
.B(n_960),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1526),
.A2(n_967),
.B1(n_968),
.B2(n_965),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1391),
.B(n_972),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1507),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1342),
.B(n_973),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1359),
.Y(n_1755)
);

BUFx4f_ASAP7_75t_L g1756 ( 
.A(n_1452),
.Y(n_1756)
);

INVx4_ASAP7_75t_L g1757 ( 
.A(n_1405),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1352),
.B(n_815),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1450),
.Y(n_1759)
);

AOI22x1_ASAP7_75t_L g1760 ( 
.A1(n_1501),
.A2(n_791),
.B1(n_792),
.B2(n_744),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1486),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1337),
.A2(n_829),
.B1(n_830),
.B2(n_823),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1487),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1530),
.A2(n_982),
.B1(n_985),
.B2(n_980),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1483),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1535),
.B(n_986),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1510),
.B(n_1511),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1481),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1441),
.B(n_987),
.Y(n_1769)
);

AND3x1_ASAP7_75t_L g1770 ( 
.A(n_1387),
.B(n_841),
.C(n_832),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1541),
.B(n_988),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1507),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1439),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1430),
.B(n_1012),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1485),
.B(n_1013),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1385),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1507),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1356),
.B(n_1023),
.Y(n_1778)
);

INVx5_ASAP7_75t_L g1779 ( 
.A(n_1452),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1566),
.A2(n_1026),
.B1(n_1016),
.B2(n_854),
.Y(n_1780)
);

AND2x6_ASAP7_75t_L g1781 ( 
.A(n_1459),
.B(n_792),
.Y(n_1781)
);

CKINVDCx8_ASAP7_75t_R g1782 ( 
.A(n_1416),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1460),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1456),
.A2(n_855),
.B1(n_856),
.B2(n_844),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1388),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1493),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1358),
.B(n_857),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1464),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1398),
.B(n_1007),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1474),
.B(n_859),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1393),
.B(n_861),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1424),
.A2(n_875),
.B1(n_878),
.B2(n_863),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1454),
.B(n_879),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1469),
.B(n_1458),
.Y(n_1794)
);

AND2x6_ASAP7_75t_SL g1795 ( 
.A(n_1491),
.B(n_885),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1470),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1471),
.Y(n_1797)
);

BUFx3_ASAP7_75t_L g1798 ( 
.A(n_1463),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1484),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1500),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1404),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1410),
.B(n_890),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1409),
.Y(n_1803)
);

INVx5_ASAP7_75t_L g1804 ( 
.A(n_1484),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1345),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1440),
.B(n_891),
.Y(n_1806)
);

BUFx8_ASAP7_75t_L g1807 ( 
.A(n_1405),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1413),
.B(n_1395),
.Y(n_1808)
);

AND2x2_ASAP7_75t_SL g1809 ( 
.A(n_1422),
.B(n_819),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_SL g1810 ( 
.A(n_1498),
.B(n_902),
.C(n_900),
.Y(n_1810)
);

INVx2_ASAP7_75t_SL g1811 ( 
.A(n_1437),
.Y(n_1811)
);

NAND2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1445),
.B(n_1468),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1415),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1423),
.B(n_917),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1429),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1411),
.B(n_919),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1475),
.A2(n_926),
.B1(n_931),
.B2(n_925),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1476),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1417),
.Y(n_1819)
);

BUFx4f_ASAP7_75t_L g1820 ( 
.A(n_1484),
.Y(n_1820)
);

BUFx4f_ASAP7_75t_L g1821 ( 
.A(n_1496),
.Y(n_1821)
);

INVx4_ASAP7_75t_L g1822 ( 
.A(n_1496),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1467),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1412),
.B(n_932),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1461),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1448),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1451),
.B(n_941),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1414),
.A2(n_946),
.B(n_943),
.Y(n_1828)
);

AND2x6_ASAP7_75t_L g1829 ( 
.A(n_1496),
.B(n_836),
.Y(n_1829)
);

NOR2xp67_ASAP7_75t_L g1830 ( 
.A(n_1414),
.B(n_21),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1480),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1489),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1492),
.B(n_951),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1499),
.A2(n_962),
.B(n_956),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1502),
.B(n_963),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1538),
.B(n_969),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1329),
.B(n_1006),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1403),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1354),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1354),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1354),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1421),
.A2(n_975),
.B(n_974),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1338),
.B(n_983),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1361),
.A2(n_992),
.B1(n_993),
.B2(n_990),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1338),
.B(n_1002),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1563),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1354),
.Y(n_1847)
);

INVx6_ASAP7_75t_L g1848 ( 
.A(n_1330),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1361),
.B(n_1005),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1329),
.B(n_1020),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1538),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1361),
.B(n_1024),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1456),
.A2(n_1028),
.B1(n_1025),
.B2(n_837),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1563),
.Y(n_1854)
);

OR2x6_ASAP7_75t_L g1855 ( 
.A(n_1654),
.B(n_836),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1626),
.B(n_837),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1610),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1696),
.A2(n_903),
.B1(n_920),
.B2(n_868),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1630),
.A2(n_1652),
.B(n_1641),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1580),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1674),
.A2(n_903),
.B(n_868),
.Y(n_1861)
);

NAND3xp33_ASAP7_75t_L g1862 ( 
.A(n_1810),
.B(n_948),
.C(n_920),
.Y(n_1862)
);

INVx4_ASAP7_75t_L g1863 ( 
.A(n_1606),
.Y(n_1863)
);

AND2x2_ASAP7_75t_SL g1864 ( 
.A(n_1606),
.B(n_948),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1588),
.A2(n_950),
.B(n_949),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_R g1866 ( 
.A(n_1619),
.B(n_25),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1584),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1696),
.B(n_961),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1586),
.A2(n_1819),
.B(n_1765),
.C(n_1748),
.Y(n_1869)
);

O2A1O1Ixp33_ASAP7_75t_L g1870 ( 
.A1(n_1717),
.A2(n_966),
.B(n_981),
.C(n_961),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1682),
.Y(n_1871)
);

AOI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1830),
.A2(n_1031),
.B(n_1019),
.Y(n_1872)
);

OR2x6_ASAP7_75t_L g1873 ( 
.A(n_1654),
.B(n_1019),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1671),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1640),
.B(n_1594),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1601),
.B(n_1031),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1755),
.A2(n_526),
.B(n_525),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1603),
.B(n_25),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1742),
.A2(n_1805),
.B(n_1828),
.Y(n_1879)
);

NOR2xp67_ASAP7_75t_SL g1880 ( 
.A(n_1848),
.B(n_27),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1604),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1803),
.B(n_28),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1599),
.B(n_28),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1607),
.B(n_1680),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1598),
.B(n_29),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1851),
.B(n_29),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1575),
.B(n_1581),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1671),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1826),
.B(n_31),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1761),
.B(n_1763),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1808),
.A2(n_528),
.B(n_527),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1636),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1678),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1675),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_L g1895 ( 
.A(n_1605),
.B(n_33),
.C(n_36),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1609),
.B(n_36),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1801),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1716),
.B(n_41),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1679),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1720),
.A2(n_544),
.B(n_543),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1676),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1648),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1611),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1695),
.A2(n_547),
.B(n_545),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1577),
.B(n_43),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1697),
.A2(n_555),
.B(n_553),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1589),
.B(n_44),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1579),
.B(n_47),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1609),
.B(n_47),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1750),
.B(n_48),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1614),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1699),
.A2(n_558),
.B(n_557),
.Y(n_1912)
);

BUFx12f_ASAP7_75t_L g1913 ( 
.A(n_1848),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1663),
.B(n_48),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1617),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1576),
.B(n_50),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1701),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1721),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1846),
.B(n_1854),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1582),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1838),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1590),
.A2(n_57),
.B1(n_54),
.B2(n_55),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1622),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1618),
.B(n_57),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1585),
.A2(n_61),
.B(n_58),
.C(n_59),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1789),
.A2(n_62),
.B(n_59),
.C(n_61),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1639),
.B(n_63),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1659),
.Y(n_1928)
);

CKINVDCx11_ASAP7_75t_R g1929 ( 
.A(n_1600),
.Y(n_1929)
);

AO21x2_ASAP7_75t_L g1930 ( 
.A1(n_1653),
.A2(n_562),
.B(n_561),
.Y(n_1930)
);

BUFx2_ASAP7_75t_L g1931 ( 
.A(n_1621),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1587),
.B(n_1749),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1843),
.B(n_65),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1733),
.B(n_65),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1845),
.B(n_66),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1745),
.B(n_67),
.Y(n_1936)
);

BUFx3_ASAP7_75t_L g1937 ( 
.A(n_1807),
.Y(n_1937)
);

NOR3xp33_ASAP7_75t_SL g1938 ( 
.A(n_1570),
.B(n_68),
.C(n_69),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1572),
.B(n_68),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1743),
.B(n_71),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1689),
.B(n_72),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1636),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1651),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1813),
.A2(n_565),
.B(n_564),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1713),
.B(n_74),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1646),
.B(n_75),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1794),
.B(n_75),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1790),
.B(n_76),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1625),
.A2(n_569),
.B(n_566),
.Y(n_1949)
);

OR2x6_ASAP7_75t_L g1950 ( 
.A(n_1600),
.B(n_76),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1722),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1844),
.B(n_77),
.Y(n_1952)
);

O2A1O1Ixp33_ASAP7_75t_L g1953 ( 
.A1(n_1793),
.A2(n_81),
.B(n_78),
.C(n_80),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1664),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1702),
.B(n_81),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1811),
.B(n_82),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1833),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1713),
.B(n_82),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1747),
.A2(n_1853),
.B(n_1784),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_R g1960 ( 
.A(n_1707),
.B(n_83),
.Y(n_1960)
);

AO32x2_ASAP7_75t_L g1961 ( 
.A1(n_1687),
.A2(n_85),
.A3(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_1961)
);

AO32x2_ASAP7_75t_L g1962 ( 
.A1(n_1723),
.A2(n_86),
.A3(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1736),
.B(n_87),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1814),
.B(n_88),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1583),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1638),
.Y(n_1966)
);

NOR2xp67_ASAP7_75t_SL g1967 ( 
.A(n_1635),
.B(n_89),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1662),
.B(n_89),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1656),
.A2(n_93),
.B1(n_90),
.B2(n_91),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1634),
.A2(n_578),
.B(n_577),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1620),
.A2(n_97),
.B1(n_94),
.B2(n_96),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1583),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1642),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1807),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_SL g1975 ( 
.A(n_1668),
.B(n_98),
.C(n_99),
.Y(n_1975)
);

AOI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1685),
.A2(n_104),
.B1(n_98),
.B2(n_100),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_L g1977 ( 
.A(n_1583),
.B(n_579),
.Y(n_1977)
);

OA22x2_ASAP7_75t_L g1978 ( 
.A1(n_1592),
.A2(n_105),
.B1(n_100),
.B2(n_104),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1721),
.B(n_106),
.Y(n_1979)
);

OAI22x1_ASAP7_75t_L g1980 ( 
.A1(n_1660),
.A2(n_110),
.B1(n_107),
.B2(n_109),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1849),
.B(n_107),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1677),
.B(n_1837),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1768),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1852),
.B(n_110),
.Y(n_1984)
);

NOR3xp33_ASAP7_75t_SL g1985 ( 
.A(n_1684),
.B(n_111),
.C(n_112),
.Y(n_1985)
);

NOR3xp33_ASAP7_75t_SL g1986 ( 
.A(n_1727),
.B(n_113),
.C(n_114),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1644),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1788),
.B(n_115),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1809),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1615),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1645),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1796),
.B(n_1797),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1637),
.A2(n_581),
.B(n_580),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1850),
.B(n_121),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1762),
.A2(n_125),
.B1(n_122),
.B2(n_124),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1836),
.B(n_126),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1643),
.A2(n_585),
.B(n_583),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1758),
.B(n_127),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1786),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1669),
.B(n_129),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1655),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1649),
.A2(n_587),
.B(n_586),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1714),
.B(n_129),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1758),
.B(n_1787),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1629),
.Y(n_2005)
);

AO21x2_ASAP7_75t_L g2006 ( 
.A1(n_1842),
.A2(n_592),
.B(n_590),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_L g2007 ( 
.A(n_1734),
.B(n_132),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1787),
.B(n_132),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1571),
.Y(n_2009)
);

A2O1A1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1834),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1779),
.B(n_133),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1824),
.B(n_135),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1715),
.Y(n_2013)
);

A2O1A1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1806),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1635),
.Y(n_2015)
);

BUFx12f_ASAP7_75t_L g2016 ( 
.A(n_1757),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1823),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1647),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1571),
.B(n_139),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1777),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1775),
.A2(n_143),
.B1(n_140),
.B2(n_142),
.Y(n_2021)
);

INVx8_ASAP7_75t_L g2022 ( 
.A(n_1829),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1827),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2023)
);

INVx4_ASAP7_75t_L g2024 ( 
.A(n_1691),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1657),
.Y(n_2025)
);

INVx6_ASAP7_75t_L g2026 ( 
.A(n_1757),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1779),
.B(n_144),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1781),
.B(n_146),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1658),
.Y(n_2029)
);

OAI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1741),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1781),
.B(n_147),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1737),
.B(n_148),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1779),
.B(n_149),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1632),
.Y(n_2034)
);

AOI21xp33_ASAP7_75t_L g2035 ( 
.A1(n_1738),
.A2(n_1778),
.B(n_1754),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1665),
.Y(n_2036)
);

CKINVDCx12_ASAP7_75t_R g2037 ( 
.A(n_1767),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_1578),
.B(n_150),
.Y(n_2038)
);

O2A1O1Ixp33_ASAP7_75t_L g2039 ( 
.A1(n_1597),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1661),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_1767),
.B(n_151),
.Y(n_2041)
);

CKINVDCx8_ASAP7_75t_R g2042 ( 
.A(n_1741),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1672),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1574),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1820),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1839),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1840),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1741),
.B(n_155),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1591),
.A2(n_158),
.B1(n_155),
.B2(n_157),
.Y(n_2049)
);

INVx4_ASAP7_75t_L g2050 ( 
.A(n_1710),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1841),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1694),
.A2(n_604),
.B(n_603),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1688),
.B(n_159),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1781),
.B(n_160),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1756),
.B(n_160),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1781),
.B(n_161),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1700),
.A2(n_606),
.B(n_605),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1704),
.A2(n_611),
.B(n_608),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1624),
.B(n_161),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1688),
.B(n_162),
.Y(n_2060)
);

A2O1A1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_1817),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_1718),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1791),
.B(n_164),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1847),
.Y(n_2064)
);

CKINVDCx20_ASAP7_75t_R g2065 ( 
.A(n_1725),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_L g2066 ( 
.A(n_1756),
.B(n_165),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1627),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1820),
.B(n_166),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1821),
.B(n_167),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1729),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_1613),
.B(n_1616),
.Y(n_2071)
);

NOR2xp33_ASAP7_75t_L g2072 ( 
.A(n_1798),
.B(n_167),
.Y(n_2072)
);

O2A1O1Ixp33_ASAP7_75t_L g2073 ( 
.A1(n_1816),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1774),
.B(n_169),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1791),
.B(n_170),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1730),
.A2(n_620),
.B(n_615),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_L g2077 ( 
.A1(n_1656),
.A2(n_173),
.B1(n_171),
.B2(n_172),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_R g2078 ( 
.A(n_1623),
.B(n_172),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1831),
.A2(n_1832),
.B(n_1744),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1802),
.B(n_175),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1821),
.B(n_176),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1802),
.B(n_176),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1683),
.B(n_177),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1731),
.Y(n_2084)
);

AO22x1_ASAP7_75t_L g2085 ( 
.A1(n_1595),
.A2(n_181),
.B1(n_178),
.B2(n_180),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1737),
.B(n_180),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1698),
.Y(n_2087)
);

NOR2xp67_ASAP7_75t_L g2088 ( 
.A(n_1650),
.B(n_182),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1708),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1624),
.B(n_183),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1596),
.B(n_184),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1740),
.B(n_1666),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1681),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1670),
.B(n_186),
.Y(n_2094)
);

AO32x1_ASAP7_75t_L g2095 ( 
.A1(n_1822),
.A2(n_188),
.A3(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1709),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1726),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1740),
.B(n_187),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1735),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1690),
.Y(n_2100)
);

CKINVDCx8_ASAP7_75t_R g2101 ( 
.A(n_1795),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1766),
.B(n_1771),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1760),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1782),
.B(n_190),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1666),
.B(n_191),
.Y(n_2105)
);

BUFx8_ASAP7_75t_SL g2106 ( 
.A(n_1728),
.Y(n_2106)
);

INVx4_ASAP7_75t_L g2107 ( 
.A(n_1804),
.Y(n_2107)
);

BUFx12f_ASAP7_75t_L g2108 ( 
.A(n_1573),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_1593),
.Y(n_2109)
);

INVx3_ASAP7_75t_SL g2110 ( 
.A(n_1728),
.Y(n_2110)
);

INVx1_ASAP7_75t_SL g2111 ( 
.A(n_1595),
.Y(n_2111)
);

BUFx3_ASAP7_75t_L g2112 ( 
.A(n_1593),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1783),
.B(n_193),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1692),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1760),
.Y(n_2115)
);

O2A1O1Ixp33_ASAP7_75t_L g2116 ( 
.A1(n_1693),
.A2(n_195),
.B(n_193),
.C(n_194),
.Y(n_2116)
);

O2A1O1Ixp33_ASAP7_75t_L g2117 ( 
.A1(n_1769),
.A2(n_198),
.B(n_194),
.C(n_197),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_SL g2118 ( 
.A(n_1703),
.B(n_635),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1792),
.B(n_197),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1612),
.A2(n_198),
.B(n_200),
.Y(n_2120)
);

OAI21xp33_ASAP7_75t_L g2121 ( 
.A1(n_1706),
.A2(n_201),
.B(n_202),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1667),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1667),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_1739),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2124)
);

NAND2x1p5_ASAP7_75t_L g2125 ( 
.A(n_1804),
.B(n_1608),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1732),
.A2(n_208),
.B(n_210),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1776),
.B(n_210),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1785),
.B(n_211),
.Y(n_2128)
);

OR2x6_ASAP7_75t_L g2129 ( 
.A(n_1759),
.B(n_510),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1773),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1719),
.B(n_212),
.Y(n_2131)
);

BUFx8_ASAP7_75t_L g2132 ( 
.A(n_1739),
.Y(n_2132)
);

INVx4_ASAP7_75t_L g2133 ( 
.A(n_1804),
.Y(n_2133)
);

CKINVDCx8_ASAP7_75t_R g2134 ( 
.A(n_1829),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1815),
.B(n_213),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_1724),
.B(n_214),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_1753),
.B(n_217),
.Y(n_2137)
);

AND3x2_ASAP7_75t_L g2138 ( 
.A(n_1770),
.B(n_217),
.C(n_218),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1602),
.B(n_1686),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1818),
.Y(n_2140)
);

AND2x4_ASAP7_75t_L g2141 ( 
.A(n_1772),
.B(n_220),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1780),
.B(n_221),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1751),
.B(n_221),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1829),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1764),
.B(n_222),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1812),
.B(n_223),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1628),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2147)
);

INVxp67_ASAP7_75t_L g2148 ( 
.A(n_1705),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1818),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1633),
.B(n_227),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1711),
.B(n_228),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1628),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_2152)
);

O2A1O1Ixp33_ASAP7_75t_L g2153 ( 
.A1(n_1752),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_1595),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1829),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_1825),
.B(n_233),
.Y(n_2156)
);

O2A1O1Ixp33_ASAP7_75t_SL g2157 ( 
.A1(n_1712),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2157)
);

INVxp67_ASAP7_75t_SL g2158 ( 
.A(n_1631),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1595),
.B(n_235),
.Y(n_2159)
);

O2A1O1Ixp33_ASAP7_75t_L g2160 ( 
.A1(n_1835),
.A2(n_239),
.B(n_236),
.C(n_238),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_1673),
.Y(n_2161)
);

AOI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_1800),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_2162)
);

BUFx2_ASAP7_75t_L g2163 ( 
.A(n_1673),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1673),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1682),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1630),
.A2(n_244),
.B(n_245),
.Y(n_2166)
);

OAI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1696),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1696),
.B(n_246),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1682),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1580),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1799),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_1598),
.Y(n_2172)
);

AO32x1_ASAP7_75t_L g2173 ( 
.A1(n_1805),
.A2(n_247),
.A3(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_1799),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_1848),
.Y(n_2175)
);

INVx2_ASAP7_75t_SL g2176 ( 
.A(n_1848),
.Y(n_2176)
);

INVx1_ASAP7_75t_SL g2177 ( 
.A(n_1610),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1682),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1618),
.B(n_250),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_1598),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_R g2181 ( 
.A(n_1619),
.B(n_251),
.Y(n_2181)
);

NOR3xp33_ASAP7_75t_SL g2182 ( 
.A(n_1605),
.B(n_252),
.C(n_255),
.Y(n_2182)
);

INVx3_ASAP7_75t_L g2183 ( 
.A(n_1713),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1826),
.B(n_256),
.Y(n_2184)
);

OAI22x1_ASAP7_75t_L g2185 ( 
.A1(n_1660),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_2185)
);

O2A1O1Ixp33_ASAP7_75t_L g2186 ( 
.A1(n_1717),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1799),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1626),
.B(n_262),
.Y(n_2188)
);

INVx4_ASAP7_75t_L g2189 ( 
.A(n_1610),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1601),
.B(n_263),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_SL g2191 ( 
.A(n_1606),
.B(n_265),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1630),
.A2(n_265),
.B(n_266),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1601),
.B(n_266),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_1590),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1630),
.A2(n_268),
.B(n_269),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_R g2196 ( 
.A(n_1619),
.B(n_271),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1696),
.B(n_272),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1696),
.B(n_274),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_SL g2199 ( 
.A1(n_1654),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2199)
);

NOR2xp33_ASAP7_75t_L g2200 ( 
.A(n_1626),
.B(n_276),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1696),
.B(n_277),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1696),
.B(n_277),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1580),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1580),
.Y(n_2204)
);

CKINVDCx6p67_ASAP7_75t_R g2205 ( 
.A(n_1675),
.Y(n_2205)
);

CKINVDCx11_ASAP7_75t_R g2206 ( 
.A(n_1619),
.Y(n_2206)
);

NAND3xp33_ASAP7_75t_L g2207 ( 
.A(n_1810),
.B(n_279),
.C(n_280),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_L g2208 ( 
.A(n_1626),
.B(n_282),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1618),
.B(n_283),
.Y(n_2209)
);

OR2x6_ASAP7_75t_L g2210 ( 
.A(n_1654),
.B(n_509),
.Y(n_2210)
);

BUFx3_ASAP7_75t_L g2211 ( 
.A(n_1610),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_1696),
.A2(n_286),
.B1(n_283),
.B2(n_284),
.Y(n_2212)
);

OAI21x1_ASAP7_75t_L g2213 ( 
.A1(n_1746),
.A2(n_287),
.B(n_288),
.Y(n_2213)
);

NOR2xp33_ASAP7_75t_R g2214 ( 
.A(n_1619),
.B(n_287),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1598),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_1626),
.B(n_289),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1696),
.B(n_290),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_1799),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1618),
.B(n_291),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_1701),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1580),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_1601),
.B(n_296),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1626),
.B(n_297),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_1619),
.Y(n_2224)
);

OAI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1696),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1580),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1618),
.B(n_300),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_1610),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1696),
.B(n_303),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1626),
.B(n_304),
.Y(n_2230)
);

NAND2x1p5_ASAP7_75t_L g2231 ( 
.A(n_1721),
.B(n_306),
.Y(n_2231)
);

AOI21xp5_ASAP7_75t_L g2232 ( 
.A1(n_1630),
.A2(n_307),
.B(n_311),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1682),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1696),
.B(n_307),
.Y(n_2234)
);

AOI21xp5_ASAP7_75t_L g2235 ( 
.A1(n_1630),
.A2(n_311),
.B(n_312),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_L g2236 ( 
.A(n_1810),
.B(n_314),
.C(n_315),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1580),
.Y(n_2237)
);

INVx2_ASAP7_75t_SL g2238 ( 
.A(n_1848),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_1713),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_1701),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_L g2241 ( 
.A1(n_1630),
.A2(n_318),
.B(n_319),
.Y(n_2241)
);

BUFx2_ASAP7_75t_L g2242 ( 
.A(n_1598),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_1626),
.B(n_319),
.Y(n_2243)
);

OR2x6_ASAP7_75t_L g2244 ( 
.A(n_1950),
.B(n_2022),
.Y(n_2244)
);

BUFx2_ASAP7_75t_SL g2245 ( 
.A(n_1937),
.Y(n_2245)
);

BUFx2_ASAP7_75t_SL g2246 ( 
.A(n_1874),
.Y(n_2246)
);

INVx1_ASAP7_75t_SL g2247 ( 
.A(n_2177),
.Y(n_2247)
);

AO21x2_ASAP7_75t_L g2248 ( 
.A1(n_2103),
.A2(n_320),
.B(n_322),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1932),
.B(n_322),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1890),
.Y(n_2250)
);

AOI21x1_ASAP7_75t_L g2251 ( 
.A1(n_2115),
.A2(n_323),
.B(n_325),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1893),
.Y(n_2252)
);

INVx5_ASAP7_75t_SL g2253 ( 
.A(n_2205),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1983),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1999),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1899),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_2107),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1860),
.Y(n_2258)
);

INVx6_ASAP7_75t_L g2259 ( 
.A(n_2189),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1867),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_2206),
.Y(n_2261)
);

OAI21x1_ASAP7_75t_L g2262 ( 
.A1(n_1872),
.A2(n_328),
.B(n_329),
.Y(n_2262)
);

INVxp67_ASAP7_75t_SL g2263 ( 
.A(n_2137),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1923),
.B(n_328),
.Y(n_2264)
);

INVx8_ASAP7_75t_L g2265 ( 
.A(n_1913),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_SL g2266 ( 
.A(n_1894),
.B(n_329),
.Y(n_2266)
);

CKINVDCx16_ASAP7_75t_R g2267 ( 
.A(n_1866),
.Y(n_2267)
);

BUFx12f_ASAP7_75t_L g2268 ( 
.A(n_1888),
.Y(n_2268)
);

CKINVDCx5p33_ASAP7_75t_R g2269 ( 
.A(n_2224),
.Y(n_2269)
);

INVx3_ASAP7_75t_L g2270 ( 
.A(n_2107),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1857),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_2133),
.Y(n_2272)
);

BUFx12f_ASAP7_75t_L g2273 ( 
.A(n_1929),
.Y(n_2273)
);

OAI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_1859),
.A2(n_332),
.B(n_333),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1887),
.B(n_333),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1881),
.Y(n_2276)
);

AO21x2_ASAP7_75t_L g2277 ( 
.A1(n_2131),
.A2(n_334),
.B(n_335),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1869),
.B(n_336),
.Y(n_2278)
);

BUFx3_ASAP7_75t_L g2279 ( 
.A(n_2211),
.Y(n_2279)
);

INVx3_ASAP7_75t_SL g2280 ( 
.A(n_2189),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_1901),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2171),
.Y(n_2282)
);

AO21x2_ASAP7_75t_L g2283 ( 
.A1(n_1879),
.A2(n_336),
.B(n_337),
.Y(n_2283)
);

BUFx2_ASAP7_75t_SL g2284 ( 
.A(n_1863),
.Y(n_2284)
);

INVxp67_ASAP7_75t_SL g2285 ( 
.A(n_2137),
.Y(n_2285)
);

BUFx2_ASAP7_75t_L g2286 ( 
.A(n_2228),
.Y(n_2286)
);

OA21x2_ASAP7_75t_L g2287 ( 
.A1(n_2213),
.A2(n_337),
.B(n_338),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2171),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2170),
.B(n_339),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2079),
.A2(n_340),
.B(n_341),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2133),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1918),
.Y(n_2292)
);

AOI22x1_ASAP7_75t_L g2293 ( 
.A1(n_1949),
.A2(n_342),
.B1(n_344),
.B2(n_347),
.Y(n_2293)
);

OR2x6_ASAP7_75t_L g2294 ( 
.A(n_1950),
.B(n_348),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_1884),
.A2(n_349),
.B(n_350),
.Y(n_2295)
);

BUFx2_ASAP7_75t_L g2296 ( 
.A(n_2180),
.Y(n_2296)
);

NAND2x1p5_ASAP7_75t_L g2297 ( 
.A(n_1863),
.B(n_349),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1923),
.B(n_351),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2171),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1918),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2203),
.B(n_351),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_2129),
.Y(n_2302)
);

OR2x6_ASAP7_75t_L g2303 ( 
.A(n_1950),
.B(n_2022),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2204),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_2045),
.B(n_353),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2221),
.B(n_354),
.Y(n_2306)
);

BUFx2_ASAP7_75t_SL g2307 ( 
.A(n_2042),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2226),
.B(n_354),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2237),
.B(n_355),
.Y(n_2309)
);

AOI22x1_ASAP7_75t_L g2310 ( 
.A1(n_1970),
.A2(n_356),
.B1(n_359),
.B2(n_360),
.Y(n_2310)
);

BUFx4f_ASAP7_75t_L g2311 ( 
.A(n_2210),
.Y(n_2311)
);

AOI22xp33_ASAP7_75t_L g2312 ( 
.A1(n_2038),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_2312)
);

BUFx12f_ASAP7_75t_L g2313 ( 
.A(n_2210),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2174),
.Y(n_2314)
);

OR2x6_ASAP7_75t_L g2315 ( 
.A(n_2022),
.B(n_2210),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1911),
.Y(n_2316)
);

OR2x6_ASAP7_75t_L g2317 ( 
.A(n_2129),
.B(n_363),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_1877),
.A2(n_364),
.B(n_367),
.Y(n_2318)
);

INVx4_ASAP7_75t_L g2319 ( 
.A(n_2016),
.Y(n_2319)
);

AO21x2_ASAP7_75t_L g2320 ( 
.A1(n_1930),
.A2(n_364),
.B(n_368),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_1915),
.B(n_368),
.Y(n_2321)
);

BUFx2_ASAP7_75t_SL g2322 ( 
.A(n_2065),
.Y(n_2322)
);

AO21x2_ASAP7_75t_L g2323 ( 
.A1(n_1930),
.A2(n_371),
.B(n_372),
.Y(n_2323)
);

INVx5_ASAP7_75t_L g2324 ( 
.A(n_2164),
.Y(n_2324)
);

BUFx2_ASAP7_75t_SL g2325 ( 
.A(n_2177),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2215),
.B(n_372),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2174),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1903),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1992),
.Y(n_2329)
);

BUFx8_ASAP7_75t_L g2330 ( 
.A(n_1990),
.Y(n_2330)
);

INVx6_ASAP7_75t_L g2331 ( 
.A(n_2034),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2009),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2125),
.Y(n_2333)
);

INVx1_ASAP7_75t_SL g2334 ( 
.A(n_2242),
.Y(n_2334)
);

INVx3_ASAP7_75t_L g2335 ( 
.A(n_2134),
.Y(n_2335)
);

AOI21xp5_ASAP7_75t_L g2336 ( 
.A1(n_1939),
.A2(n_375),
.B(n_376),
.Y(n_2336)
);

AOI22x1_ASAP7_75t_L g2337 ( 
.A1(n_1993),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_2337)
);

OAI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2168),
.A2(n_379),
.B(n_381),
.Y(n_2338)
);

BUFx3_ASAP7_75t_L g2339 ( 
.A(n_2125),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_2108),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2187),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1966),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2197),
.A2(n_382),
.B(n_383),
.Y(n_2343)
);

NAND2x1p5_ASAP7_75t_L g2344 ( 
.A(n_2045),
.B(n_382),
.Y(n_2344)
);

AO21x1_ASAP7_75t_L g2345 ( 
.A1(n_2156),
.A2(n_1989),
.B(n_2186),
.Y(n_2345)
);

OR2x2_ASAP7_75t_L g2346 ( 
.A(n_2004),
.B(n_1931),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1973),
.Y(n_2347)
);

INVx2_ASAP7_75t_SL g2348 ( 
.A(n_2132),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_1965),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2218),
.Y(n_2350)
);

OAI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2198),
.A2(n_384),
.B(n_385),
.Y(n_2351)
);

AO21x2_ASAP7_75t_L g2352 ( 
.A1(n_2006),
.A2(n_386),
.B(n_387),
.Y(n_2352)
);

BUFx2_ASAP7_75t_SL g2353 ( 
.A(n_2175),
.Y(n_2353)
);

OA21x2_ASAP7_75t_L g2354 ( 
.A1(n_1891),
.A2(n_390),
.B(n_391),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1987),
.Y(n_2355)
);

AO21x1_ASAP7_75t_L g2356 ( 
.A1(n_2156),
.A2(n_391),
.B(n_392),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_1964),
.A2(n_393),
.B(n_394),
.Y(n_2357)
);

AOI22x1_ASAP7_75t_L g2358 ( 
.A1(n_1997),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_2358)
);

BUFx12f_ASAP7_75t_L g2359 ( 
.A(n_2132),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1875),
.B(n_397),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2184),
.B(n_397),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_1972),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2005),
.Y(n_2363)
);

OAI21xp5_ASAP7_75t_L g2364 ( 
.A1(n_2201),
.A2(n_398),
.B(n_399),
.Y(n_2364)
);

AO21x2_ASAP7_75t_L g2365 ( 
.A1(n_2006),
.A2(n_398),
.B(n_400),
.Y(n_2365)
);

AOI22x1_ASAP7_75t_L g2366 ( 
.A1(n_2002),
.A2(n_401),
.B1(n_403),
.B2(n_405),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1991),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2001),
.Y(n_2368)
);

OAI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2183),
.A2(n_401),
.B(n_406),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_1864),
.B(n_406),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2025),
.Y(n_2371)
);

INVx3_ASAP7_75t_SL g2372 ( 
.A(n_2110),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2029),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2018),
.Y(n_2374)
);

CKINVDCx20_ASAP7_75t_R g2375 ( 
.A(n_2106),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_1933),
.A2(n_408),
.B(n_410),
.Y(n_2376)
);

INVx6_ASAP7_75t_L g2377 ( 
.A(n_2024),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2172),
.B(n_408),
.Y(n_2378)
);

INVx1_ASAP7_75t_SL g2379 ( 
.A(n_2013),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_1928),
.Y(n_2380)
);

BUFx2_ASAP7_75t_SL g2381 ( 
.A(n_2176),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2040),
.Y(n_2382)
);

NAND2x1p5_ASAP7_75t_L g2383 ( 
.A(n_2141),
.B(n_414),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2129),
.Y(n_2384)
);

INVx1_ASAP7_75t_SL g2385 ( 
.A(n_2013),
.Y(n_2385)
);

NAND2x1p5_ASAP7_75t_L g2386 ( 
.A(n_2141),
.B(n_417),
.Y(n_2386)
);

BUFx2_ASAP7_75t_R g2387 ( 
.A(n_2101),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2239),
.A2(n_418),
.B(n_419),
.Y(n_2388)
);

AO21x2_ASAP7_75t_L g2389 ( 
.A1(n_2202),
.A2(n_419),
.B(n_420),
.Y(n_2389)
);

OA21x2_ASAP7_75t_L g2390 ( 
.A1(n_1904),
.A2(n_420),
.B(n_421),
.Y(n_2390)
);

INVx6_ASAP7_75t_SL g2391 ( 
.A(n_1855),
.Y(n_2391)
);

OR2x6_ASAP7_75t_L g2392 ( 
.A(n_1855),
.B(n_421),
.Y(n_2392)
);

OA21x2_ASAP7_75t_L g2393 ( 
.A1(n_1906),
.A2(n_422),
.B(n_424),
.Y(n_2393)
);

OAI21x1_ASAP7_75t_L g2394 ( 
.A1(n_2239),
.A2(n_422),
.B(n_425),
.Y(n_2394)
);

INVx6_ASAP7_75t_L g2395 ( 
.A(n_2024),
.Y(n_2395)
);

OA21x2_ASAP7_75t_L g2396 ( 
.A1(n_1912),
.A2(n_425),
.B(n_426),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2184),
.B(n_426),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_1855),
.Y(n_2398)
);

INVx3_ASAP7_75t_SL g2399 ( 
.A(n_1873),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_1873),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2043),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2036),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2136),
.Y(n_2403)
);

OA21x2_ASAP7_75t_L g2404 ( 
.A1(n_1900),
.A2(n_427),
.B(n_429),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2071),
.B(n_2044),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_1920),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_2136),
.Y(n_2407)
);

OAI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2217),
.A2(n_427),
.B(n_429),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2229),
.A2(n_430),
.B(n_431),
.Y(n_2409)
);

INVx4_ASAP7_75t_L g2410 ( 
.A(n_1873),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_1996),
.B(n_431),
.Y(n_2411)
);

AO21x2_ASAP7_75t_L g2412 ( 
.A1(n_2234),
.A2(n_434),
.B(n_435),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_2181),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2046),
.B(n_434),
.Y(n_2414)
);

NAND2x1p5_ASAP7_75t_L g2415 ( 
.A(n_2050),
.B(n_436),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2047),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2051),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2064),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_1921),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_2032),
.Y(n_2420)
);

NAND2x1p5_ASAP7_75t_L g2421 ( 
.A(n_2050),
.B(n_439),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2026),
.Y(n_2422)
);

CKINVDCx8_ASAP7_75t_R g2423 ( 
.A(n_2093),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2084),
.B(n_441),
.Y(n_2424)
);

OA21x2_ASAP7_75t_L g2425 ( 
.A1(n_1944),
.A2(n_442),
.B(n_443),
.Y(n_2425)
);

HB1xp67_ASAP7_75t_L g2426 ( 
.A(n_2032),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_2026),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2096),
.Y(n_2428)
);

NAND2x1p5_ASAP7_75t_L g2429 ( 
.A(n_2144),
.B(n_2163),
.Y(n_2429)
);

INVx1_ASAP7_75t_SL g2430 ( 
.A(n_2078),
.Y(n_2430)
);

OAI21x1_ASAP7_75t_L g2431 ( 
.A1(n_2052),
.A2(n_2058),
.B(n_2057),
.Y(n_2431)
);

BUFx2_ASAP7_75t_SL g2432 ( 
.A(n_2238),
.Y(n_2432)
);

AOI22x1_ASAP7_75t_L g2433 ( 
.A1(n_2076),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_2196),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2231),
.Y(n_2435)
);

BUFx4_ASAP7_75t_SL g2436 ( 
.A(n_2155),
.Y(n_2436)
);

INVx5_ASAP7_75t_L g2437 ( 
.A(n_2100),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_1862),
.A2(n_449),
.B(n_450),
.Y(n_2438)
);

AOI22x1_ASAP7_75t_L g2439 ( 
.A1(n_1865),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_2439)
);

INVx4_ASAP7_75t_L g2440 ( 
.A(n_2231),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2097),
.Y(n_2441)
);

INVx4_ASAP7_75t_L g2442 ( 
.A(n_2100),
.Y(n_2442)
);

AO21x2_ASAP7_75t_L g2443 ( 
.A1(n_2086),
.A2(n_454),
.B(n_455),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_2070),
.Y(n_2444)
);

BUFx2_ASAP7_75t_R g2445 ( 
.A(n_1896),
.Y(n_2445)
);

HB1xp67_ASAP7_75t_L g2446 ( 
.A(n_2099),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2139),
.B(n_454),
.Y(n_2447)
);

OAI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_1862),
.A2(n_456),
.B(n_457),
.Y(n_2448)
);

INVx1_ASAP7_75t_SL g2449 ( 
.A(n_2059),
.Y(n_2449)
);

INVxp67_ASAP7_75t_SL g2450 ( 
.A(n_2100),
.Y(n_2450)
);

INVx3_ASAP7_75t_SL g2451 ( 
.A(n_2062),
.Y(n_2451)
);

CKINVDCx20_ASAP7_75t_R g2452 ( 
.A(n_2214),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2114),
.Y(n_2453)
);

OA21x2_ASAP7_75t_L g2454 ( 
.A1(n_2120),
.A2(n_456),
.B(n_459),
.Y(n_2454)
);

OR2x6_ASAP7_75t_L g2455 ( 
.A(n_1974),
.B(n_459),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2130),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2225),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_L g2458 ( 
.A1(n_1968),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_2458)
);

NOR2x1_ASAP7_75t_SL g2459 ( 
.A(n_1989),
.B(n_460),
.Y(n_2459)
);

AO21x2_ASAP7_75t_L g2460 ( 
.A1(n_2098),
.A2(n_461),
.B(n_462),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2225),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2087),
.Y(n_2462)
);

OAI21x1_ASAP7_75t_L g2463 ( 
.A1(n_1945),
.A2(n_463),
.B(n_464),
.Y(n_2463)
);

BUFx2_ASAP7_75t_R g2464 ( 
.A(n_1909),
.Y(n_2464)
);

HB1xp67_ASAP7_75t_L g2465 ( 
.A(n_1871),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1957),
.B(n_465),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_2089),
.B(n_465),
.Y(n_2467)
);

NAND2x1p5_ASAP7_75t_L g2468 ( 
.A(n_2111),
.B(n_466),
.Y(n_2468)
);

INVx2_ASAP7_75t_SL g2469 ( 
.A(n_2015),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2165),
.Y(n_2470)
);

OAI21xp5_ASAP7_75t_L g2471 ( 
.A1(n_1861),
.A2(n_466),
.B(n_467),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_SL g2472 ( 
.A(n_2112),
.Y(n_2472)
);

INVx1_ASAP7_75t_SL g2473 ( 
.A(n_2090),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_1963),
.Y(n_2474)
);

OAI21x1_ASAP7_75t_SL g2475 ( 
.A1(n_2122),
.A2(n_468),
.B(n_469),
.Y(n_2475)
);

OAI21x1_ASAP7_75t_L g2476 ( 
.A1(n_1958),
.A2(n_468),
.B(n_470),
.Y(n_2476)
);

INVx6_ASAP7_75t_SL g2477 ( 
.A(n_2037),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2169),
.Y(n_2478)
);

BUFx2_ASAP7_75t_SL g2479 ( 
.A(n_2088),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_2178),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2233),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1878),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2067),
.Y(n_2483)
);

INVxp67_ASAP7_75t_SL g2484 ( 
.A(n_2161),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_1883),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2102),
.B(n_472),
.Y(n_2486)
);

NAND2x1p5_ASAP7_75t_L g2487 ( 
.A(n_2111),
.B(n_473),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_1924),
.B(n_473),
.Y(n_2488)
);

OR2x6_ASAP7_75t_L g2489 ( 
.A(n_2085),
.B(n_474),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2154),
.B(n_474),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_1892),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_1960),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_1868),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2179),
.B(n_475),
.Y(n_2494)
);

AO21x2_ASAP7_75t_L g2495 ( 
.A1(n_2113),
.A2(n_476),
.B(n_477),
.Y(n_2495)
);

BUFx12f_ASAP7_75t_L g2496 ( 
.A(n_1940),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_SL g2497 ( 
.A(n_2140),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1905),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_1908),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_1942),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1882),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1898),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_1889),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2209),
.B(n_478),
.Y(n_2504)
);

OAI21xp5_ASAP7_75t_L g2505 ( 
.A1(n_2166),
.A2(n_479),
.B(n_480),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_1954),
.Y(n_2506)
);

AO21x2_ASAP7_75t_L g2507 ( 
.A1(n_1870),
.A2(n_480),
.B(n_481),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2199),
.Y(n_2508)
);

BUFx2_ASAP7_75t_L g2509 ( 
.A(n_1982),
.Y(n_2509)
);

CKINVDCx12_ASAP7_75t_R g2510 ( 
.A(n_2199),
.Y(n_2510)
);

BUFx3_ASAP7_75t_L g2511 ( 
.A(n_2109),
.Y(n_2511)
);

OAI21x1_ASAP7_75t_L g2512 ( 
.A1(n_2159),
.A2(n_483),
.B(n_484),
.Y(n_2512)
);

OR2x2_ASAP7_75t_L g2513 ( 
.A(n_2219),
.B(n_484),
.Y(n_2513)
);

BUFx12f_ASAP7_75t_L g2514 ( 
.A(n_2094),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2092),
.Y(n_2515)
);

INVx4_ASAP7_75t_L g2516 ( 
.A(n_2138),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2227),
.B(n_485),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_1943),
.B(n_486),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_1935),
.B(n_487),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_1988),
.Y(n_2520)
);

BUFx2_ASAP7_75t_R g2521 ( 
.A(n_2150),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_1995),
.Y(n_2522)
);

NAND2x1p5_ASAP7_75t_L g2523 ( 
.A(n_1880),
.B(n_490),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2149),
.Y(n_2524)
);

BUFx2_ASAP7_75t_L g2525 ( 
.A(n_2158),
.Y(n_2525)
);

BUFx2_ASAP7_75t_L g2526 ( 
.A(n_2003),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_1948),
.B(n_490),
.Y(n_2527)
);

OAI21x1_ASAP7_75t_L g2528 ( 
.A1(n_1979),
.A2(n_491),
.B(n_493),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_2072),
.Y(n_2529)
);

NAND2x1p5_ASAP7_75t_L g2530 ( 
.A(n_1967),
.B(n_494),
.Y(n_2530)
);

AO21x2_ASAP7_75t_L g2531 ( 
.A1(n_2012),
.A2(n_495),
.B(n_496),
.Y(n_2531)
);

BUFx3_ASAP7_75t_L g2532 ( 
.A(n_2028),
.Y(n_2532)
);

INVx4_ASAP7_75t_L g2533 ( 
.A(n_1978),
.Y(n_2533)
);

INVx4_ASAP7_75t_L g2534 ( 
.A(n_2191),
.Y(n_2534)
);

OAI21x1_ASAP7_75t_SL g2535 ( 
.A1(n_2122),
.A2(n_497),
.B(n_498),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_1961),
.Y(n_2536)
);

OAI21x1_ASAP7_75t_L g2537 ( 
.A1(n_2192),
.A2(n_497),
.B(n_499),
.Y(n_2537)
);

NOR2x1_ASAP7_75t_R g2538 ( 
.A(n_2191),
.B(n_500),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_2151),
.Y(n_2539)
);

AO21x1_ASAP7_75t_L g2540 ( 
.A1(n_2123),
.A2(n_500),
.B(n_501),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_1947),
.B(n_502),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_1995),
.Y(n_2542)
);

AOI22x1_ASAP7_75t_L g2543 ( 
.A1(n_2195),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_1856),
.B(n_505),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_1961),
.Y(n_2545)
);

INVxp67_ASAP7_75t_SL g2546 ( 
.A(n_2123),
.Y(n_2546)
);

INVx3_ASAP7_75t_SL g2547 ( 
.A(n_1919),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2000),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_1994),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2031),
.Y(n_2550)
);

OR2x6_ASAP7_75t_L g2551 ( 
.A(n_1959),
.B(n_507),
.Y(n_2551)
);

NOR2x1_ASAP7_75t_R g2552 ( 
.A(n_1910),
.B(n_508),
.Y(n_2552)
);

INVx2_ASAP7_75t_SL g2553 ( 
.A(n_1907),
.Y(n_2553)
);

BUFx2_ASAP7_75t_L g2554 ( 
.A(n_2054),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2056),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2483),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_L g2557 ( 
.A1(n_2551),
.A2(n_1914),
.B1(n_1927),
.B2(n_2243),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2483),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2536),
.Y(n_2559)
);

NAND2x1p5_ASAP7_75t_L g2560 ( 
.A(n_2340),
.B(n_2048),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2296),
.Y(n_2561)
);

BUFx3_ASAP7_75t_L g2562 ( 
.A(n_2265),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2325),
.Y(n_2563)
);

BUFx10_ASAP7_75t_L g2564 ( 
.A(n_2261),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2440),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2536),
.Y(n_2566)
);

INVx2_ASAP7_75t_SL g2567 ( 
.A(n_2265),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_2265),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2440),
.Y(n_2569)
);

AOI21x1_ASAP7_75t_L g2570 ( 
.A1(n_2345),
.A2(n_2193),
.B(n_2190),
.Y(n_2570)
);

CKINVDCx11_ASAP7_75t_R g2571 ( 
.A(n_2359),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2533),
.B(n_2035),
.Y(n_2572)
);

HB1xp67_ASAP7_75t_L g2573 ( 
.A(n_2334),
.Y(n_2573)
);

CKINVDCx20_ASAP7_75t_R g2574 ( 
.A(n_2375),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2545),
.Y(n_2575)
);

INVx6_ASAP7_75t_L g2576 ( 
.A(n_2340),
.Y(n_2576)
);

INVx5_ASAP7_75t_L g2577 ( 
.A(n_2359),
.Y(n_2577)
);

CKINVDCx14_ASAP7_75t_R g2578 ( 
.A(n_2375),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2545),
.Y(n_2579)
);

CKINVDCx20_ASAP7_75t_R g2580 ( 
.A(n_2261),
.Y(n_2580)
);

OAI22xp5_ASAP7_75t_L g2581 ( 
.A1(n_2263),
.A2(n_2207),
.B1(n_2236),
.B2(n_1959),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2250),
.B(n_2188),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2254),
.Y(n_2583)
);

INVx5_ASAP7_75t_L g2584 ( 
.A(n_2253),
.Y(n_2584)
);

OAI21xp5_ASAP7_75t_SL g2585 ( 
.A1(n_2430),
.A2(n_2236),
.B(n_2207),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2405),
.B(n_2200),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2332),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2405),
.B(n_2329),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2255),
.Y(n_2589)
);

OR2x6_ASAP7_75t_L g2590 ( 
.A(n_2294),
.B(n_2244),
.Y(n_2590)
);

CKINVDCx11_ASAP7_75t_R g2591 ( 
.A(n_2268),
.Y(n_2591)
);

NAND2x1p5_ASAP7_75t_L g2592 ( 
.A(n_2311),
.B(n_2319),
.Y(n_2592)
);

AOI22xp33_ASAP7_75t_L g2593 ( 
.A1(n_2551),
.A2(n_2216),
.B1(n_2208),
.B2(n_2230),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2258),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2333),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2268),
.Y(n_2596)
);

OAI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2263),
.A2(n_2021),
.B1(n_1976),
.B2(n_2223),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_SL g2598 ( 
.A1(n_2508),
.A2(n_2041),
.B1(n_2055),
.B2(n_2066),
.Y(n_2598)
);

AO21x1_ASAP7_75t_SL g2599 ( 
.A1(n_2435),
.A2(n_2063),
.B(n_1998),
.Y(n_2599)
);

OAI21x1_ASAP7_75t_L g2600 ( 
.A1(n_2431),
.A2(n_2241),
.B(n_2235),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2333),
.Y(n_2601)
);

OR2x2_ASAP7_75t_L g2602 ( 
.A(n_2346),
.B(n_1885),
.Y(n_2602)
);

AOI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2551),
.A2(n_1895),
.B1(n_1946),
.B2(n_2091),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2285),
.A2(n_1922),
.B1(n_2194),
.B2(n_1971),
.Y(n_2604)
);

AOI22xp5_ASAP7_75t_L g2605 ( 
.A1(n_2447),
.A2(n_1934),
.B1(n_1981),
.B2(n_1984),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2260),
.Y(n_2606)
);

AO21x1_ASAP7_75t_SL g2607 ( 
.A1(n_2435),
.A2(n_2008),
.B(n_2075),
.Y(n_2607)
);

BUFx3_ASAP7_75t_L g2608 ( 
.A(n_2280),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2437),
.Y(n_2609)
);

BUFx2_ASAP7_75t_L g2610 ( 
.A(n_2391),
.Y(n_2610)
);

BUFx3_ASAP7_75t_L g2611 ( 
.A(n_2280),
.Y(n_2611)
);

AOI21x1_ASAP7_75t_L g2612 ( 
.A1(n_2302),
.A2(n_2222),
.B(n_2069),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2276),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2304),
.Y(n_2614)
);

AOI21x1_ASAP7_75t_L g2615 ( 
.A1(n_2302),
.A2(n_2068),
.B(n_2081),
.Y(n_2615)
);

BUFx3_ASAP7_75t_L g2616 ( 
.A(n_2372),
.Y(n_2616)
);

AOI21x1_ASAP7_75t_L g2617 ( 
.A1(n_2384),
.A2(n_2019),
.B(n_2060),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2339),
.Y(n_2618)
);

NAND2x1p5_ASAP7_75t_L g2619 ( 
.A(n_2311),
.B(n_2053),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2339),
.Y(n_2620)
);

AOI22xp33_ASAP7_75t_L g2621 ( 
.A1(n_2533),
.A2(n_2074),
.B1(n_2121),
.B2(n_1980),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2508),
.B(n_2514),
.Y(n_2622)
);

AOI21x1_ASAP7_75t_L g2623 ( 
.A1(n_2384),
.A2(n_2146),
.B(n_1876),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2406),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2406),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2316),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2419),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2416),
.Y(n_2628)
);

AOI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_2313),
.A2(n_2185),
.B1(n_2083),
.B2(n_2145),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2332),
.Y(n_2630)
);

OAI22xp5_ASAP7_75t_L g2631 ( 
.A1(n_2285),
.A2(n_2049),
.B1(n_1951),
.B2(n_2220),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2417),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_SL g2633 ( 
.A(n_2294),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2418),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2447),
.A2(n_1936),
.B1(n_2007),
.B2(n_2135),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2317),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2534),
.B(n_2030),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2294),
.A2(n_2104),
.B1(n_1952),
.B2(n_1955),
.Y(n_2638)
);

AO21x1_ASAP7_75t_L g2639 ( 
.A1(n_2534),
.A2(n_2017),
.B(n_2020),
.Y(n_2639)
);

INVx6_ASAP7_75t_L g2640 ( 
.A(n_2259),
.Y(n_2640)
);

CKINVDCx20_ASAP7_75t_R g2641 ( 
.A(n_2253),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2453),
.Y(n_2642)
);

HB1xp67_ASAP7_75t_L g2643 ( 
.A(n_2317),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2363),
.Y(n_2644)
);

AO21x1_ASAP7_75t_SL g2645 ( 
.A1(n_2420),
.A2(n_2082),
.B(n_2080),
.Y(n_2645)
);

INVx4_ASAP7_75t_L g2646 ( 
.A(n_2372),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2456),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2317),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2252),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2256),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2328),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2342),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2259),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_SL g2654 ( 
.A1(n_2459),
.A2(n_1897),
.B1(n_2167),
.B2(n_2212),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2347),
.Y(n_2655)
);

BUFx8_ASAP7_75t_L g2656 ( 
.A(n_2273),
.Y(n_2656)
);

OAI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2244),
.A2(n_2240),
.B1(n_1917),
.B2(n_2124),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_SL g2658 ( 
.A1(n_2313),
.A2(n_2011),
.B1(n_2027),
.B2(n_2033),
.Y(n_2658)
);

NAND2x1p5_ASAP7_75t_L g2659 ( 
.A(n_2319),
.B(n_1916),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2355),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2367),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2510),
.A2(n_2119),
.B1(n_1986),
.B2(n_1938),
.Y(n_2662)
);

BUFx2_ASAP7_75t_L g2663 ( 
.A(n_2391),
.Y(n_2663)
);

AOI22xp33_ASAP7_75t_SL g2664 ( 
.A1(n_2479),
.A2(n_2383),
.B1(n_2386),
.B2(n_2361),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2539),
.A2(n_2142),
.B1(n_2143),
.B2(n_2105),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2446),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2437),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2374),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2249),
.B(n_2446),
.Y(n_2669)
);

HB1xp67_ASAP7_75t_L g2670 ( 
.A(n_2465),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2368),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2371),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2373),
.Y(n_2673)
);

CKINVDCx20_ASAP7_75t_R g2674 ( 
.A(n_2253),
.Y(n_2674)
);

INVx6_ASAP7_75t_L g2675 ( 
.A(n_2259),
.Y(n_2675)
);

INVxp67_ASAP7_75t_L g2676 ( 
.A(n_2286),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2275),
.A2(n_2023),
.B1(n_2126),
.B2(n_2232),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2257),
.Y(n_2678)
);

BUFx2_ASAP7_75t_L g2679 ( 
.A(n_2391),
.Y(n_2679)
);

BUFx8_ASAP7_75t_SL g2680 ( 
.A(n_2273),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2275),
.B(n_1858),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_SL g2682 ( 
.A(n_2455),
.Y(n_2682)
);

INVx3_ASAP7_75t_L g2683 ( 
.A(n_2257),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2382),
.Y(n_2684)
);

BUFx2_ASAP7_75t_SL g2685 ( 
.A(n_2348),
.Y(n_2685)
);

BUFx6f_ASAP7_75t_L g2686 ( 
.A(n_2437),
.Y(n_2686)
);

OAI21x1_ASAP7_75t_SL g2687 ( 
.A1(n_2475),
.A2(n_2073),
.B(n_1953),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2486),
.B(n_1886),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2402),
.Y(n_2689)
);

INVx1_ASAP7_75t_SL g2690 ( 
.A(n_2271),
.Y(n_2690)
);

INVx5_ASAP7_75t_L g2691 ( 
.A(n_2244),
.Y(n_2691)
);

BUFx12f_ASAP7_75t_L g2692 ( 
.A(n_2269),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2402),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2478),
.Y(n_2694)
);

NAND2x1p5_ASAP7_75t_L g2695 ( 
.A(n_2271),
.B(n_2279),
.Y(n_2695)
);

BUFx2_ASAP7_75t_R g2696 ( 
.A(n_2269),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2478),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2457),
.Y(n_2698)
);

OAI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2486),
.A2(n_1902),
.B(n_2117),
.Y(n_2699)
);

NAND2x1p5_ASAP7_75t_L g2700 ( 
.A(n_2279),
.B(n_1956),
.Y(n_2700)
);

OAI21x1_ASAP7_75t_SL g2701 ( 
.A1(n_2535),
.A2(n_1925),
.B(n_2039),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2461),
.Y(n_2702)
);

AO21x1_ASAP7_75t_L g2703 ( 
.A1(n_2468),
.A2(n_2152),
.B(n_2147),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2428),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2441),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2401),
.Y(n_2706)
);

OR2x6_ASAP7_75t_L g2707 ( 
.A(n_2303),
.B(n_2148),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2524),
.Y(n_2708)
);

BUFx8_ASAP7_75t_L g2709 ( 
.A(n_2492),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2524),
.Y(n_2710)
);

INVx6_ASAP7_75t_L g2711 ( 
.A(n_2330),
.Y(n_2711)
);

CKINVDCx11_ASAP7_75t_R g2712 ( 
.A(n_2423),
.Y(n_2712)
);

INVx3_ASAP7_75t_L g2713 ( 
.A(n_2270),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2400),
.B(n_1985),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2370),
.B(n_2182),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2510),
.A2(n_1975),
.B1(n_1941),
.B2(n_1969),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2462),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2392),
.A2(n_2077),
.B1(n_2127),
.B2(n_2128),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2283),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2283),
.Y(n_2720)
);

BUFx12f_ASAP7_75t_L g2721 ( 
.A(n_2330),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2470),
.Y(n_2722)
);

NAND2x1p5_ASAP7_75t_L g2723 ( 
.A(n_2400),
.B(n_2118),
.Y(n_2723)
);

NAND2x1p5_ASAP7_75t_L g2724 ( 
.A(n_2410),
.B(n_2118),
.Y(n_2724)
);

BUFx6f_ASAP7_75t_L g2725 ( 
.A(n_2437),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2411),
.B(n_1926),
.Y(n_2726)
);

AND2x4_ASAP7_75t_L g2727 ( 
.A(n_2303),
.B(n_2315),
.Y(n_2727)
);

BUFx12f_ASAP7_75t_L g2728 ( 
.A(n_2380),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2331),
.Y(n_2729)
);

HB1xp67_ASAP7_75t_L g2730 ( 
.A(n_2465),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2245),
.Y(n_2731)
);

INVx6_ASAP7_75t_L g2732 ( 
.A(n_2331),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2281),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2481),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2480),
.Y(n_2735)
);

AOI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2392),
.A2(n_2162),
.B1(n_1977),
.B2(n_2116),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2480),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2287),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2246),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2392),
.A2(n_2529),
.B1(n_2548),
.B2(n_2361),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2320),
.Y(n_2741)
);

INVx6_ASAP7_75t_L g2742 ( 
.A(n_2331),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2264),
.B(n_2298),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2491),
.Y(n_2744)
);

OAI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2438),
.A2(n_2160),
.B(n_2153),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2491),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2500),
.Y(n_2747)
);

CKINVDCx5p33_ASAP7_75t_R g2748 ( 
.A(n_2413),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2320),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2451),
.Y(n_2750)
);

BUFx4f_ASAP7_75t_SL g2751 ( 
.A(n_2477),
.Y(n_2751)
);

HB1xp67_ASAP7_75t_L g2752 ( 
.A(n_2379),
.Y(n_2752)
);

INVx11_ASAP7_75t_L g2753 ( 
.A(n_2496),
.Y(n_2753)
);

OAI21x1_ASAP7_75t_SL g2754 ( 
.A1(n_2540),
.A2(n_1962),
.B(n_1961),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2500),
.Y(n_2755)
);

BUFx2_ASAP7_75t_L g2756 ( 
.A(n_2303),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2323),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2506),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2397),
.B(n_2326),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2270),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2451),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2323),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2352),
.Y(n_2763)
);

BUFx12f_ASAP7_75t_L g2764 ( 
.A(n_2380),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2385),
.B(n_2014),
.Y(n_2765)
);

AO21x1_ASAP7_75t_L g2766 ( 
.A1(n_2468),
.A2(n_1962),
.B(n_2095),
.Y(n_2766)
);

HB1xp67_ASAP7_75t_L g2767 ( 
.A(n_2247),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2315),
.A2(n_2061),
.B1(n_2010),
.B2(n_1962),
.Y(n_2768)
);

BUFx12f_ASAP7_75t_L g2769 ( 
.A(n_2455),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2449),
.B(n_2157),
.Y(n_2770)
);

BUFx10_ASAP7_75t_L g2771 ( 
.A(n_2455),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2397),
.B(n_2173),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2352),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2365),
.Y(n_2774)
);

NAND2x1_ASAP7_75t_L g2775 ( 
.A(n_2442),
.B(n_2095),
.Y(n_2775)
);

BUFx3_ASAP7_75t_L g2776 ( 
.A(n_2377),
.Y(n_2776)
);

CKINVDCx11_ASAP7_75t_R g2777 ( 
.A(n_2413),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2477),
.Y(n_2778)
);

AOI22xp33_ASAP7_75t_SL g2779 ( 
.A1(n_2383),
.A2(n_2173),
.B1(n_2386),
.B2(n_2410),
.Y(n_2779)
);

CKINVDCx11_ASAP7_75t_R g2780 ( 
.A(n_2434),
.Y(n_2780)
);

OAI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2315),
.A2(n_2173),
.B1(n_2399),
.B2(n_2266),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2369),
.Y(n_2782)
);

BUFx2_ASAP7_75t_R g2783 ( 
.A(n_2322),
.Y(n_2783)
);

OAI21x1_ASAP7_75t_SL g2784 ( 
.A1(n_2274),
.A2(n_2295),
.B(n_2356),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_L g2785 ( 
.A1(n_2529),
.A2(n_2548),
.B1(n_2549),
.B2(n_2516),
.Y(n_2785)
);

NAND2x1p5_ASAP7_75t_L g2786 ( 
.A(n_2444),
.B(n_2474),
.Y(n_2786)
);

INVx1_ASAP7_75t_SL g2787 ( 
.A(n_2399),
.Y(n_2787)
);

HB1xp67_ASAP7_75t_L g2788 ( 
.A(n_2420),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2388),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2377),
.Y(n_2790)
);

AND2x4_ASAP7_75t_L g2791 ( 
.A(n_2272),
.B(n_2291),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2394),
.Y(n_2792)
);

CKINVDCx8_ASAP7_75t_R g2793 ( 
.A(n_2267),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2278),
.Y(n_2794)
);

BUFx3_ASAP7_75t_L g2795 ( 
.A(n_2377),
.Y(n_2795)
);

BUFx2_ASAP7_75t_R g2796 ( 
.A(n_2307),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2526),
.B(n_2509),
.Y(n_2797)
);

INVx5_ASAP7_75t_L g2798 ( 
.A(n_2489),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2378),
.B(n_2473),
.Y(n_2799)
);

AOI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2549),
.A2(n_2434),
.B1(n_2452),
.B2(n_2426),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2516),
.B(n_2398),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2546),
.A2(n_2426),
.B1(n_2407),
.B2(n_2403),
.Y(n_2802)
);

CKINVDCx11_ASAP7_75t_R g2803 ( 
.A(n_2452),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2278),
.Y(n_2804)
);

OA21x2_ASAP7_75t_L g2805 ( 
.A1(n_2262),
.A2(n_2290),
.B(n_2546),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2248),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2248),
.Y(n_2807)
);

AOI22xp33_ASAP7_75t_L g2808 ( 
.A1(n_2549),
.A2(n_2522),
.B1(n_2542),
.B2(n_2489),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2274),
.Y(n_2809)
);

INVx1_ASAP7_75t_SL g2810 ( 
.A(n_2353),
.Y(n_2810)
);

AOI22xp33_ASAP7_75t_L g2811 ( 
.A1(n_2544),
.A2(n_2541),
.B1(n_2407),
.B2(n_2403),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2395),
.Y(n_2812)
);

BUFx2_ASAP7_75t_SL g2813 ( 
.A(n_2472),
.Y(n_2813)
);

AOI22xp33_ASAP7_75t_L g2814 ( 
.A1(n_2501),
.A2(n_2502),
.B1(n_2503),
.B2(n_2498),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_2387),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2289),
.Y(n_2816)
);

OR2x6_ASAP7_75t_L g2817 ( 
.A(n_2721),
.B(n_2284),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2743),
.B(n_2321),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2706),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2669),
.B(n_2797),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2799),
.B(n_2321),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2759),
.B(n_2414),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2706),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2633),
.A2(n_2301),
.B1(n_2309),
.B2(n_2414),
.Y(n_2824)
);

AO31x2_ASAP7_75t_L g2825 ( 
.A1(n_2766),
.A2(n_2350),
.A3(n_2299),
.B(n_2314),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2670),
.B(n_2513),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2590),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2624),
.Y(n_2828)
);

CKINVDCx16_ASAP7_75t_R g2829 ( 
.A(n_2641),
.Y(n_2829)
);

CKINVDCx16_ASAP7_75t_R g2830 ( 
.A(n_2674),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2730),
.B(n_2301),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2588),
.B(n_2814),
.Y(n_2832)
);

OAI22xp33_ASAP7_75t_L g2833 ( 
.A1(n_2590),
.A2(n_2798),
.B1(n_2769),
.B2(n_2636),
.Y(n_2833)
);

HB1xp67_ASAP7_75t_L g2834 ( 
.A(n_2666),
.Y(n_2834)
);

CKINVDCx5p33_ASAP7_75t_R g2835 ( 
.A(n_2571),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_R g2836 ( 
.A(n_2731),
.B(n_2335),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2625),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2798),
.B(n_2525),
.Y(n_2838)
);

NAND2xp33_ASAP7_75t_R g2839 ( 
.A(n_2739),
.B(n_2301),
.Y(n_2839)
);

INVxp67_ASAP7_75t_L g2840 ( 
.A(n_2608),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2627),
.Y(n_2841)
);

OR2x2_ASAP7_75t_L g2842 ( 
.A(n_2587),
.B(n_2309),
.Y(n_2842)
);

OAI22xp33_ASAP7_75t_L g2843 ( 
.A1(n_2798),
.A2(n_2297),
.B1(n_2421),
.B2(n_2415),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2594),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2630),
.B(n_2309),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2606),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2690),
.B(n_2488),
.Y(n_2847)
);

BUFx2_ASAP7_75t_L g2848 ( 
.A(n_2750),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2613),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2556),
.B(n_2511),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_R g2851 ( 
.A(n_2577),
.B(n_2335),
.Y(n_2851)
);

OAI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2664),
.A2(n_2421),
.B1(n_2415),
.B2(n_2297),
.Y(n_2852)
);

HB1xp67_ASAP7_75t_L g2853 ( 
.A(n_2561),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2614),
.Y(n_2854)
);

NAND2xp33_ASAP7_75t_R g2855 ( 
.A(n_2815),
.B(n_2467),
.Y(n_2855)
);

AND2x4_ASAP7_75t_L g2856 ( 
.A(n_2691),
.B(n_2272),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2695),
.B(n_2715),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_R g2858 ( 
.A(n_2577),
.B(n_2751),
.Y(n_2858)
);

BUFx3_ASAP7_75t_L g2859 ( 
.A(n_2562),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_R g2860 ( 
.A(n_2577),
.B(n_2591),
.Y(n_2860)
);

INVxp67_ASAP7_75t_SL g2861 ( 
.A(n_2556),
.Y(n_2861)
);

INVxp67_ASAP7_75t_L g2862 ( 
.A(n_2611),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2633),
.B(n_2496),
.Y(n_2863)
);

NOR2x1_ASAP7_75t_L g2864 ( 
.A(n_2646),
.B(n_2291),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2717),
.B(n_2494),
.Y(n_2865)
);

AND2x4_ASAP7_75t_L g2866 ( 
.A(n_2691),
.B(n_2292),
.Y(n_2866)
);

INVx5_ASAP7_75t_L g2867 ( 
.A(n_2584),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2761),
.Y(n_2868)
);

INVxp67_ASAP7_75t_SL g2869 ( 
.A(n_2558),
.Y(n_2869)
);

INVxp67_ASAP7_75t_L g2870 ( 
.A(n_2733),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2626),
.Y(n_2871)
);

AND2x4_ASAP7_75t_L g2872 ( 
.A(n_2691),
.B(n_2292),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2727),
.B(n_2558),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2682),
.A2(n_2458),
.B1(n_2518),
.B2(n_2554),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2628),
.B(n_2466),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_R g2876 ( 
.A(n_2568),
.B(n_2300),
.Y(n_2876)
);

HB1xp67_ASAP7_75t_L g2877 ( 
.A(n_2573),
.Y(n_2877)
);

NOR3xp33_ASAP7_75t_SL g2878 ( 
.A(n_2596),
.B(n_2295),
.C(n_2336),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2584),
.Y(n_2879)
);

INVx6_ASAP7_75t_L g2880 ( 
.A(n_2584),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2727),
.B(n_2300),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2722),
.B(n_2504),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2734),
.B(n_2517),
.Y(n_2883)
);

NOR2xp33_ASAP7_75t_R g2884 ( 
.A(n_2574),
.B(n_2472),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2708),
.Y(n_2885)
);

CKINVDCx12_ASAP7_75t_R g2886 ( 
.A(n_2656),
.Y(n_2886)
);

OR2x6_ASAP7_75t_L g2887 ( 
.A(n_2592),
.B(n_2305),
.Y(n_2887)
);

AOI22xp5_ASAP7_75t_SL g2888 ( 
.A1(n_2578),
.A2(n_2381),
.B1(n_2432),
.B2(n_2553),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2632),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2634),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2704),
.B(n_2467),
.Y(n_2891)
);

AND2x4_ASAP7_75t_L g2892 ( 
.A(n_2565),
.B(n_2518),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2705),
.B(n_2518),
.Y(n_2893)
);

AND2x2_ASAP7_75t_L g2894 ( 
.A(n_2642),
.B(n_2511),
.Y(n_2894)
);

AO31x2_ASAP7_75t_L g2895 ( 
.A1(n_2741),
.A2(n_2757),
.A3(n_2762),
.B(n_2749),
.Y(n_2895)
);

INVx2_ASAP7_75t_SL g2896 ( 
.A(n_2576),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2576),
.Y(n_2897)
);

NAND2x1p5_ASAP7_75t_L g2898 ( 
.A(n_2646),
.B(n_2616),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2647),
.Y(n_2899)
);

NOR3xp33_ASAP7_75t_SL g2900 ( 
.A(n_2748),
.B(n_2336),
.C(n_2357),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2649),
.Y(n_2901)
);

AOI22xp33_ASAP7_75t_L g2902 ( 
.A1(n_2682),
.A2(n_2458),
.B1(n_2312),
.B2(n_2448),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2752),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_L g2904 ( 
.A(n_2572),
.B(n_2643),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2657),
.A2(n_2482),
.B1(n_2499),
.B2(n_2485),
.Y(n_2905)
);

NAND2xp33_ASAP7_75t_R g2906 ( 
.A(n_2565),
.B(n_2538),
.Y(n_2906)
);

HB1xp67_ASAP7_75t_L g2907 ( 
.A(n_2767),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2650),
.B(n_2466),
.Y(n_2908)
);

INVx4_ASAP7_75t_L g2909 ( 
.A(n_2753),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2651),
.B(n_2515),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2710),
.B(n_2360),
.Y(n_2911)
);

INVx8_ASAP7_75t_L g2912 ( 
.A(n_2680),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2652),
.B(n_2305),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2655),
.B(n_2344),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2656),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2567),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2660),
.Y(n_2917)
);

BUFx6f_ASAP7_75t_L g2918 ( 
.A(n_2609),
.Y(n_2918)
);

NAND3xp33_ASAP7_75t_SL g2919 ( 
.A(n_2629),
.B(n_2523),
.C(n_2530),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2661),
.B(n_2344),
.Y(n_2920)
);

CKINVDCx14_ASAP7_75t_R g2921 ( 
.A(n_2580),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2671),
.B(n_2360),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2672),
.Y(n_2923)
);

NOR2x1p5_ASAP7_75t_L g2924 ( 
.A(n_2569),
.B(n_2477),
.Y(n_2924)
);

INVxp67_ASAP7_75t_L g2925 ( 
.A(n_2685),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2673),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2569),
.B(n_2532),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2667),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2684),
.B(n_2289),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2776),
.B(n_2395),
.Y(n_2930)
);

INVx3_ASAP7_75t_L g2931 ( 
.A(n_2812),
.Y(n_2931)
);

INVx8_ASAP7_75t_L g2932 ( 
.A(n_2692),
.Y(n_2932)
);

CKINVDCx5p33_ASAP7_75t_R g2933 ( 
.A(n_2712),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2795),
.B(n_2602),
.Y(n_2934)
);

HB1xp67_ASAP7_75t_L g2935 ( 
.A(n_2648),
.Y(n_2935)
);

NOR3xp33_ASAP7_75t_SL g2936 ( 
.A(n_2714),
.B(n_2357),
.C(n_2376),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2603),
.A2(n_2439),
.B1(n_2543),
.B2(n_2493),
.Y(n_2937)
);

INVxp33_ASAP7_75t_SL g2938 ( 
.A(n_2777),
.Y(n_2938)
);

CKINVDCx5p33_ASAP7_75t_R g2939 ( 
.A(n_2780),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2583),
.Y(n_2940)
);

HB1xp67_ASAP7_75t_L g2941 ( 
.A(n_2788),
.Y(n_2941)
);

INVx1_ASAP7_75t_SL g2942 ( 
.A(n_2810),
.Y(n_2942)
);

BUFx2_ASAP7_75t_L g2943 ( 
.A(n_2812),
.Y(n_2943)
);

NAND2xp33_ASAP7_75t_R g2944 ( 
.A(n_2778),
.B(n_2756),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2729),
.B(n_2395),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2791),
.B(n_2532),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2790),
.B(n_2338),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2653),
.B(n_2338),
.Y(n_2948)
);

CKINVDCx16_ASAP7_75t_R g2949 ( 
.A(n_2728),
.Y(n_2949)
);

BUFx3_ASAP7_75t_L g2950 ( 
.A(n_2711),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2593),
.A2(n_2520),
.B1(n_2471),
.B2(n_2409),
.Y(n_2951)
);

NOR3xp33_ASAP7_75t_SL g2952 ( 
.A(n_2801),
.B(n_2376),
.C(n_2387),
.Y(n_2952)
);

CKINVDCx16_ASAP7_75t_R g2953 ( 
.A(n_2764),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2589),
.Y(n_2954)
);

OAI21x1_ASAP7_75t_L g2955 ( 
.A1(n_2600),
.A2(n_2251),
.B(n_2318),
.Y(n_2955)
);

OAI22xp5_ASAP7_75t_L g2956 ( 
.A1(n_2740),
.A2(n_2490),
.B1(n_2487),
.B2(n_2530),
.Y(n_2956)
);

NAND2xp33_ASAP7_75t_R g2957 ( 
.A(n_2622),
.B(n_2390),
.Y(n_2957)
);

AOI21xp33_ASAP7_75t_L g2958 ( 
.A1(n_2581),
.A2(n_2552),
.B(n_2519),
.Y(n_2958)
);

BUFx6f_ASAP7_75t_L g2959 ( 
.A(n_2667),
.Y(n_2959)
);

OR2x2_ASAP7_75t_L g2960 ( 
.A(n_2694),
.B(n_2306),
.Y(n_2960)
);

CKINVDCx11_ASAP7_75t_R g2961 ( 
.A(n_2564),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2816),
.B(n_2306),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2698),
.B(n_2308),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_2803),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2662),
.A2(n_2527),
.B1(n_2519),
.B2(n_2550),
.Y(n_2965)
);

CKINVDCx5p33_ASAP7_75t_R g2966 ( 
.A(n_2564),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_2711),
.Y(n_2967)
);

AO31x2_ASAP7_75t_L g2968 ( 
.A1(n_2741),
.A2(n_2327),
.A3(n_2341),
.B(n_2314),
.Y(n_2968)
);

AND2x4_ASAP7_75t_L g2969 ( 
.A(n_2791),
.B(n_2450),
.Y(n_2969)
);

INVx3_ASAP7_75t_L g2970 ( 
.A(n_2640),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2698),
.B(n_2308),
.Y(n_2971)
);

AOI21x1_ASAP7_75t_L g2972 ( 
.A1(n_2775),
.A2(n_2354),
.B(n_2393),
.Y(n_2972)
);

INVx3_ASAP7_75t_L g2973 ( 
.A(n_2640),
.Y(n_2973)
);

OAI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2557),
.A2(n_2487),
.B1(n_2490),
.B2(n_2523),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_SL g2975 ( 
.A1(n_2793),
.A2(n_2547),
.B1(n_2422),
.B2(n_2427),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_L g2976 ( 
.A1(n_2654),
.A2(n_2639),
.B1(n_2597),
.B2(n_2598),
.Y(n_2976)
);

CKINVDCx16_ASAP7_75t_R g2977 ( 
.A(n_2813),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2676),
.B(n_2343),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2595),
.B(n_2343),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_R g2980 ( 
.A(n_2771),
.B(n_2547),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2702),
.B(n_2424),
.Y(n_2981)
);

HB1xp67_ASAP7_75t_L g2982 ( 
.A(n_2697),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2595),
.B(n_2351),
.Y(n_2983)
);

BUFx2_ASAP7_75t_R g2984 ( 
.A(n_2610),
.Y(n_2984)
);

NOR2x1_ASAP7_75t_SL g2985 ( 
.A(n_2707),
.B(n_2324),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2585),
.A2(n_2505),
.B(n_2537),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2601),
.B(n_2351),
.Y(n_2987)
);

CKINVDCx14_ASAP7_75t_R g2988 ( 
.A(n_2771),
.Y(n_2988)
);

NOR2xp33_ASAP7_75t_R g2989 ( 
.A(n_2709),
.B(n_2349),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2744),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2746),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_R g2992 ( 
.A(n_2709),
.B(n_2349),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2605),
.A2(n_2505),
.B(n_2471),
.Y(n_2993)
);

CKINVDCx5p33_ASAP7_75t_R g2994 ( 
.A(n_2696),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2747),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2755),
.Y(n_2996)
);

AO31x2_ASAP7_75t_L g2997 ( 
.A1(n_2749),
.A2(n_2762),
.A3(n_2763),
.B(n_2757),
.Y(n_2997)
);

CKINVDCx16_ASAP7_75t_R g2998 ( 
.A(n_2796),
.Y(n_2998)
);

OR2x6_ASAP7_75t_L g2999 ( 
.A(n_2707),
.B(n_2429),
.Y(n_2999)
);

AO31x2_ASAP7_75t_L g3000 ( 
.A1(n_2763),
.A2(n_2327),
.A3(n_2341),
.B(n_2299),
.Y(n_3000)
);

AOI22xp33_ASAP7_75t_L g3001 ( 
.A1(n_2808),
.A2(n_2409),
.B1(n_2408),
.B2(n_2364),
.Y(n_3001)
);

AOI21xp33_ASAP7_75t_L g3002 ( 
.A1(n_2687),
.A2(n_2527),
.B(n_2507),
.Y(n_3002)
);

BUFx3_ASAP7_75t_L g3003 ( 
.A(n_2732),
.Y(n_3003)
);

CKINVDCx20_ASAP7_75t_R g3004 ( 
.A(n_2787),
.Y(n_3004)
);

NOR2xp33_ASAP7_75t_R g3005 ( 
.A(n_2601),
.B(n_2362),
.Y(n_3005)
);

OAI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2621),
.A2(n_2464),
.B1(n_2445),
.B2(n_2364),
.Y(n_3006)
);

AO31x2_ASAP7_75t_L g3007 ( 
.A1(n_2773),
.A2(n_2350),
.A3(n_2282),
.B(n_2288),
.Y(n_3007)
);

BUFx6f_ASAP7_75t_L g3008 ( 
.A(n_2686),
.Y(n_3008)
);

NAND2xp33_ASAP7_75t_R g3009 ( 
.A(n_2663),
.B(n_2390),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2686),
.B(n_2324),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2758),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2686),
.B(n_2324),
.Y(n_3012)
);

OR2x6_ASAP7_75t_L g3013 ( 
.A(n_2675),
.B(n_2429),
.Y(n_3013)
);

NOR3xp33_ASAP7_75t_SL g3014 ( 
.A(n_2688),
.B(n_2408),
.C(n_2424),
.Y(n_3014)
);

OR2x2_ASAP7_75t_L g3015 ( 
.A(n_2735),
.B(n_2737),
.Y(n_3015)
);

NOR3xp33_ASAP7_75t_SL g3016 ( 
.A(n_2586),
.B(n_2521),
.C(n_2436),
.Y(n_3016)
);

INVx4_ASAP7_75t_L g3017 ( 
.A(n_2675),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_R g3018 ( 
.A(n_2618),
.B(n_2362),
.Y(n_3018)
);

BUFx2_ASAP7_75t_SL g3019 ( 
.A(n_2618),
.Y(n_3019)
);

HB1xp67_ASAP7_75t_L g3020 ( 
.A(n_2644),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_R g3021 ( 
.A(n_2620),
.B(n_2725),
.Y(n_3021)
);

CKINVDCx5p33_ASAP7_75t_R g3022 ( 
.A(n_2783),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2604),
.A2(n_2555),
.B1(n_2550),
.B2(n_2293),
.Y(n_3023)
);

AOI21xp33_ASAP7_75t_L g3024 ( 
.A1(n_2784),
.A2(n_2768),
.B(n_2701),
.Y(n_3024)
);

CKINVDCx11_ASAP7_75t_R g3025 ( 
.A(n_2679),
.Y(n_3025)
);

OAI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2635),
.A2(n_2366),
.B1(n_2337),
.B2(n_2358),
.Y(n_3026)
);

CKINVDCx5p33_ASAP7_75t_R g3027 ( 
.A(n_2800),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2726),
.B(n_2531),
.Y(n_3028)
);

INVxp33_ASAP7_75t_SL g3029 ( 
.A(n_2785),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2668),
.Y(n_3030)
);

NAND2xp33_ASAP7_75t_SL g3031 ( 
.A(n_2725),
.B(n_2443),
.Y(n_3031)
);

AO31x2_ASAP7_75t_L g3032 ( 
.A1(n_2774),
.A2(n_2425),
.A3(n_2404),
.B(n_2390),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_2732),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_3020),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2876),
.Y(n_3035)
);

AO21x2_ASAP7_75t_L g3036 ( 
.A1(n_3002),
.A2(n_2781),
.B(n_2754),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_3021),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2844),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2820),
.B(n_2772),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2846),
.Y(n_3040)
);

AND2x4_ASAP7_75t_L g3041 ( 
.A(n_2861),
.B(n_2559),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2850),
.Y(n_3042)
);

AND2x2_ASAP7_75t_L g3043 ( 
.A(n_2818),
.B(n_2811),
.Y(n_3043)
);

HB1xp67_ASAP7_75t_L g3044 ( 
.A(n_2869),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2849),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2854),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2885),
.Y(n_3047)
);

BUFx3_ASAP7_75t_L g3048 ( 
.A(n_2859),
.Y(n_3048)
);

INVx2_ASAP7_75t_SL g3049 ( 
.A(n_2817),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2821),
.B(n_2563),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_3029),
.B(n_2765),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2873),
.B(n_2559),
.Y(n_3052)
);

INVxp67_ASAP7_75t_SL g3053 ( 
.A(n_2982),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2934),
.B(n_2689),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2871),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2894),
.B(n_2693),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2889),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2822),
.B(n_2678),
.Y(n_3058)
);

BUFx3_ASAP7_75t_L g3059 ( 
.A(n_2817),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2890),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2847),
.B(n_2904),
.Y(n_3061)
);

OAI211xp5_ASAP7_75t_SL g3062 ( 
.A1(n_2976),
.A2(n_2716),
.B(n_2638),
.C(n_2582),
.Y(n_3062)
);

INVxp67_ASAP7_75t_SL g3063 ( 
.A(n_2834),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2865),
.B(n_2882),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2828),
.Y(n_3065)
);

NAND2x1p5_ASAP7_75t_SL g3066 ( 
.A(n_2864),
.B(n_2637),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2883),
.B(n_2678),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2837),
.Y(n_3068)
);

OR2x2_ASAP7_75t_L g3069 ( 
.A(n_2941),
.B(n_2802),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2841),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2899),
.Y(n_3071)
);

OR2x2_ASAP7_75t_L g3072 ( 
.A(n_2853),
.B(n_2566),
.Y(n_3072)
);

AND2x4_ASAP7_75t_L g3073 ( 
.A(n_2873),
.B(n_2969),
.Y(n_3073)
);

INVx4_ASAP7_75t_L g3074 ( 
.A(n_2867),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2845),
.B(n_2683),
.Y(n_3075)
);

OR2x2_ASAP7_75t_L g3076 ( 
.A(n_2903),
.B(n_2566),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_3028),
.B(n_2794),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2901),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2917),
.Y(n_3079)
);

OR2x2_ASAP7_75t_L g3080 ( 
.A(n_2907),
.B(n_2575),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2927),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2923),
.Y(n_3082)
);

INVx4_ASAP7_75t_L g3083 ( 
.A(n_2867),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2910),
.B(n_2683),
.Y(n_3084)
);

INVx3_ASAP7_75t_L g3085 ( 
.A(n_2927),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_2968),
.Y(n_3086)
);

OR2x2_ASAP7_75t_L g3087 ( 
.A(n_2877),
.B(n_2575),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_2826),
.B(n_2579),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2926),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_2968),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2819),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_2831),
.B(n_2713),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2823),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2848),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2940),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2954),
.Y(n_3096)
);

INVx3_ASAP7_75t_SL g3097 ( 
.A(n_2909),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_2905),
.A2(n_2681),
.B1(n_2699),
.B2(n_2631),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2857),
.B(n_2713),
.Y(n_3099)
);

HB1xp67_ASAP7_75t_L g3100 ( 
.A(n_2968),
.Y(n_3100)
);

HB1xp67_ASAP7_75t_L g3101 ( 
.A(n_3000),
.Y(n_3101)
);

INVx2_ASAP7_75t_SL g3102 ( 
.A(n_2858),
.Y(n_3102)
);

HB1xp67_ASAP7_75t_L g3103 ( 
.A(n_3000),
.Y(n_3103)
);

NOR2x1_ASAP7_75t_L g3104 ( 
.A(n_2919),
.B(n_2760),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_2969),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2892),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_3015),
.B(n_2760),
.Y(n_3107)
);

OR2x2_ASAP7_75t_L g3108 ( 
.A(n_2870),
.B(n_2579),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2935),
.Y(n_3109)
);

OAI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2993),
.A2(n_2779),
.B(n_2745),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_SL g3111 ( 
.A1(n_2852),
.A2(n_2809),
.B1(n_2619),
.B2(n_2805),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2978),
.B(n_2832),
.Y(n_3112)
);

AND2x4_ASAP7_75t_L g3113 ( 
.A(n_2924),
.B(n_2946),
.Y(n_3113)
);

OR2x2_ASAP7_75t_L g3114 ( 
.A(n_2842),
.B(n_2942),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2963),
.B(n_2804),
.Y(n_3115)
);

AOI22xp33_ASAP7_75t_L g3116 ( 
.A1(n_3006),
.A2(n_2902),
.B1(n_2958),
.B2(n_2951),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2971),
.B(n_2809),
.Y(n_3117)
);

NOR2x1_ASAP7_75t_L g3118 ( 
.A(n_2843),
.B(n_2495),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2990),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2991),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2893),
.B(n_2645),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2995),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2996),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_3011),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2891),
.B(n_2484),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_3001),
.A2(n_2703),
.B1(n_2665),
.B2(n_2677),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_2943),
.B(n_2484),
.Y(n_3127)
);

AND2x4_ASAP7_75t_L g3128 ( 
.A(n_2946),
.B(n_2719),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2981),
.B(n_2720),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2827),
.B(n_2725),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2913),
.B(n_2443),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_3000),
.Y(n_3132)
);

HB1xp67_ASAP7_75t_L g3133 ( 
.A(n_3007),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2914),
.B(n_2460),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3030),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2920),
.Y(n_3136)
);

OAI22xp33_ASAP7_75t_L g3137 ( 
.A1(n_2839),
.A2(n_2723),
.B1(n_2724),
.B2(n_2770),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2911),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2960),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2929),
.Y(n_3140)
);

BUFx2_ASAP7_75t_L g3141 ( 
.A(n_3005),
.Y(n_3141)
);

BUFx3_ASAP7_75t_L g3142 ( 
.A(n_2868),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_3027),
.B(n_2700),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2979),
.B(n_2738),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2983),
.B(n_2806),
.Y(n_3145)
);

BUFx2_ASAP7_75t_L g3146 ( 
.A(n_3018),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2947),
.B(n_2460),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2987),
.B(n_2806),
.Y(n_3148)
);

INVx4_ASAP7_75t_R g3149 ( 
.A(n_2916),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2922),
.B(n_2786),
.Y(n_3150)
);

OR2x2_ASAP7_75t_L g3151 ( 
.A(n_2875),
.B(n_2807),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2908),
.Y(n_3152)
);

INVx4_ASAP7_75t_L g3153 ( 
.A(n_2867),
.Y(n_3153)
);

INVxp67_ASAP7_75t_L g3154 ( 
.A(n_2957),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_3019),
.B(n_2807),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2948),
.B(n_2495),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_2892),
.B(n_2782),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2881),
.B(n_2277),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2881),
.B(n_2277),
.Y(n_3159)
);

OR2x2_ASAP7_75t_L g3160 ( 
.A(n_2840),
.B(n_2389),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2962),
.Y(n_3161)
);

INVxp67_ASAP7_75t_L g3162 ( 
.A(n_3031),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2895),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2895),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_3044),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_3039),
.B(n_2862),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3044),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3112),
.B(n_2997),
.Y(n_3168)
);

AND2x4_ASAP7_75t_L g3169 ( 
.A(n_3053),
.B(n_2825),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_3112),
.B(n_2997),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3063),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3138),
.B(n_3139),
.Y(n_3172)
);

INVx3_ASAP7_75t_R g3173 ( 
.A(n_3035),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_3077),
.B(n_3117),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3061),
.B(n_2945),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3063),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3038),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3064),
.B(n_2930),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3040),
.Y(n_3179)
);

HB1xp67_ASAP7_75t_L g3180 ( 
.A(n_3053),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3045),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_3074),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_3050),
.B(n_2988),
.Y(n_3183)
);

BUFx3_ASAP7_75t_L g3184 ( 
.A(n_3048),
.Y(n_3184)
);

OAI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_3116),
.A2(n_2824),
.B1(n_2874),
.B2(n_3023),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_3077),
.B(n_2997),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_3117),
.B(n_3024),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3140),
.B(n_2825),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_3042),
.B(n_3092),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3075),
.B(n_2898),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3046),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_3034),
.B(n_2931),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_3073),
.B(n_2925),
.Y(n_3193)
);

NAND2x1_ASAP7_75t_L g3194 ( 
.A(n_3149),
.B(n_2880),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3152),
.B(n_3032),
.Y(n_3195)
);

OR2x2_ASAP7_75t_L g3196 ( 
.A(n_3072),
.B(n_2977),
.Y(n_3196)
);

INVxp67_ASAP7_75t_SL g3197 ( 
.A(n_3086),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_3041),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3055),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_3041),
.Y(n_3200)
);

AND2x4_ASAP7_75t_L g3201 ( 
.A(n_3157),
.B(n_3128),
.Y(n_3201)
);

INVx3_ASAP7_75t_L g3202 ( 
.A(n_3074),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3057),
.Y(n_3203)
);

INVxp67_ASAP7_75t_L g3204 ( 
.A(n_3160),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3147),
.B(n_3032),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_3073),
.B(n_2896),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_3065),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3060),
.Y(n_3208)
);

OR2x2_ASAP7_75t_L g3209 ( 
.A(n_3076),
.B(n_2829),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3071),
.Y(n_3210)
);

AND2x4_ASAP7_75t_SL g3211 ( 
.A(n_3113),
.B(n_3004),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_3067),
.B(n_2897),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3078),
.Y(n_3213)
);

INVxp67_ASAP7_75t_SL g3214 ( 
.A(n_3086),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_3079),
.Y(n_3215)
);

NAND2x1_ASAP7_75t_L g3216 ( 
.A(n_3149),
.B(n_2880),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_3068),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_3094),
.B(n_2938),
.Y(n_3218)
);

OAI211xp5_ASAP7_75t_L g3219 ( 
.A1(n_3116),
.A2(n_2860),
.B(n_2980),
.C(n_2851),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3114),
.B(n_3003),
.Y(n_3220)
);

NAND3xp33_ASAP7_75t_L g3221 ( 
.A(n_3110),
.B(n_2900),
.C(n_2878),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3052),
.B(n_2888),
.Y(n_3222)
);

OR2x2_ASAP7_75t_L g3223 ( 
.A(n_3080),
.B(n_2830),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3156),
.B(n_3032),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3070),
.Y(n_3225)
);

INVx1_ASAP7_75t_SL g3226 ( 
.A(n_3142),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_3082),
.Y(n_3227)
);

OR2x2_ASAP7_75t_L g3228 ( 
.A(n_3087),
.B(n_3088),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_3089),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3091),
.Y(n_3230)
);

OA21x2_ASAP7_75t_L g3231 ( 
.A1(n_3154),
.A2(n_2955),
.B(n_2986),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_3052),
.B(n_2970),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3115),
.B(n_3014),
.Y(n_3233)
);

HB1xp67_ASAP7_75t_L g3234 ( 
.A(n_3054),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3136),
.B(n_2973),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3093),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3058),
.B(n_2950),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3108),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3109),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_3037),
.Y(n_3240)
);

AND2x4_ASAP7_75t_L g3241 ( 
.A(n_3157),
.B(n_2838),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3095),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3096),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_3084),
.B(n_2998),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_3097),
.Y(n_3245)
);

HB1xp67_ASAP7_75t_L g3246 ( 
.A(n_3047),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_3245),
.B(n_3059),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3207),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3187),
.B(n_3161),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3171),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_3217),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3176),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_3201),
.B(n_3154),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3189),
.B(n_3131),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3177),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3205),
.B(n_3134),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_3205),
.B(n_3224),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_3225),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3224),
.B(n_3090),
.Y(n_3259)
);

AND2x2_ASAP7_75t_SL g3260 ( 
.A(n_3201),
.B(n_3141),
.Y(n_3260)
);

HB1xp67_ASAP7_75t_L g3261 ( 
.A(n_3165),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_3168),
.B(n_3090),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3179),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3181),
.Y(n_3264)
);

INVxp67_ASAP7_75t_L g3265 ( 
.A(n_3240),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3187),
.B(n_3145),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3168),
.B(n_3100),
.Y(n_3267)
);

BUFx2_ASAP7_75t_L g3268 ( 
.A(n_3165),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_3182),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3170),
.B(n_3100),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_3246),
.Y(n_3271)
);

NOR2x1_ASAP7_75t_L g3272 ( 
.A(n_3184),
.B(n_3146),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3170),
.B(n_3174),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3233),
.B(n_3145),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_3174),
.B(n_3101),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3191),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3234),
.B(n_3101),
.Y(n_3277)
);

AND2x4_ASAP7_75t_L g3278 ( 
.A(n_3204),
.B(n_3162),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3180),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3199),
.Y(n_3280)
);

AND2x2_ASAP7_75t_L g3281 ( 
.A(n_3198),
.B(n_3103),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_3226),
.B(n_3118),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3200),
.B(n_3103),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3203),
.Y(n_3284)
);

CKINVDCx16_ASAP7_75t_R g3285 ( 
.A(n_3183),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3204),
.B(n_3162),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3208),
.Y(n_3287)
);

CKINVDCx5p33_ASAP7_75t_R g3288 ( 
.A(n_3226),
.Y(n_3288)
);

AND2x2_ASAP7_75t_L g3289 ( 
.A(n_3166),
.B(n_3132),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3246),
.Y(n_3290)
);

INVx3_ASAP7_75t_L g3291 ( 
.A(n_3182),
.Y(n_3291)
);

AND2x4_ASAP7_75t_L g3292 ( 
.A(n_3241),
.B(n_3128),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3180),
.Y(n_3293)
);

INVxp67_ASAP7_75t_SL g3294 ( 
.A(n_3167),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3233),
.B(n_3238),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3195),
.B(n_3132),
.Y(n_3296)
);

HB1xp67_ASAP7_75t_L g3297 ( 
.A(n_3228),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3210),
.Y(n_3298)
);

AND2x4_ASAP7_75t_L g3299 ( 
.A(n_3241),
.B(n_3163),
.Y(n_3299)
);

INVx1_ASAP7_75t_SL g3300 ( 
.A(n_3211),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_3195),
.B(n_3186),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3239),
.B(n_3148),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3172),
.B(n_3148),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3186),
.B(n_3133),
.Y(n_3304)
);

HB1xp67_ASAP7_75t_L g3305 ( 
.A(n_3178),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3230),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3172),
.B(n_3110),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_3236),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3213),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_SL g3310 ( 
.A(n_3202),
.B(n_3111),
.Y(n_3310)
);

NAND4xp25_ASAP7_75t_L g3311 ( 
.A(n_3221),
.B(n_3126),
.C(n_3098),
.D(n_3051),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3268),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3306),
.Y(n_3313)
);

OR2x2_ASAP7_75t_L g3314 ( 
.A(n_3297),
.B(n_3257),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_3288),
.Y(n_3315)
);

OR2x2_ASAP7_75t_L g3316 ( 
.A(n_3257),
.B(n_3188),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3273),
.B(n_3301),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3306),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3308),
.Y(n_3319)
);

INVx1_ASAP7_75t_SL g3320 ( 
.A(n_3288),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3308),
.Y(n_3321)
);

INVxp67_ASAP7_75t_SL g3322 ( 
.A(n_3261),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_3305),
.B(n_3188),
.Y(n_3323)
);

OR2x2_ASAP7_75t_L g3324 ( 
.A(n_3274),
.B(n_3144),
.Y(n_3324)
);

OA222x2_ASAP7_75t_L g3325 ( 
.A1(n_3269),
.A2(n_3173),
.B1(n_3196),
.B2(n_3202),
.C1(n_3069),
.C2(n_3209),
.Y(n_3325)
);

NAND4xp75_ASAP7_75t_L g3326 ( 
.A(n_3260),
.B(n_3272),
.C(n_3310),
.D(n_3282),
.Y(n_3326)
);

HB1xp67_ASAP7_75t_L g3327 ( 
.A(n_3268),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3273),
.B(n_3215),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3295),
.Y(n_3329)
);

OAI32xp33_ASAP7_75t_L g3330 ( 
.A1(n_3285),
.A2(n_3223),
.A3(n_3218),
.B1(n_3222),
.B2(n_2944),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3250),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_3253),
.B(n_3175),
.Y(n_3332)
);

AND2x2_ASAP7_75t_L g3333 ( 
.A(n_3253),
.B(n_3193),
.Y(n_3333)
);

NAND3xp33_ASAP7_75t_L g3334 ( 
.A(n_3311),
.B(n_3126),
.C(n_3219),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_3253),
.B(n_3206),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3252),
.Y(n_3336)
);

OR2x2_ASAP7_75t_L g3337 ( 
.A(n_3275),
.B(n_3144),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3289),
.B(n_3232),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3255),
.Y(n_3339)
);

OAI32xp33_ASAP7_75t_L g3340 ( 
.A1(n_3300),
.A2(n_2855),
.A3(n_3083),
.B1(n_3153),
.B2(n_2906),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3263),
.Y(n_3341)
);

NAND2x1_ASAP7_75t_L g3342 ( 
.A(n_3269),
.B(n_3169),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3301),
.B(n_3227),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3264),
.Y(n_3344)
);

INVx2_ASAP7_75t_SL g3345 ( 
.A(n_3260),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3276),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3271),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3271),
.Y(n_3348)
);

NOR2x1p5_ASAP7_75t_SL g3349 ( 
.A(n_3279),
.B(n_3164),
.Y(n_3349)
);

INVx1_ASAP7_75t_SL g3350 ( 
.A(n_3269),
.Y(n_3350)
);

NOR2x1_ASAP7_75t_L g3351 ( 
.A(n_3282),
.B(n_3219),
.Y(n_3351)
);

AND2x2_ASAP7_75t_L g3352 ( 
.A(n_3289),
.B(n_3220),
.Y(n_3352)
);

AND2x4_ASAP7_75t_L g3353 ( 
.A(n_3278),
.B(n_3169),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3275),
.B(n_3229),
.Y(n_3354)
);

AOI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_3307),
.A2(n_3185),
.B1(n_3051),
.B2(n_3062),
.Y(n_3355)
);

AOI32xp33_ASAP7_75t_L g3356 ( 
.A1(n_3310),
.A2(n_3185),
.A3(n_3137),
.B1(n_3049),
.B2(n_3104),
.Y(n_3356)
);

AOI22xp5_ASAP7_75t_L g3357 ( 
.A1(n_3249),
.A2(n_3062),
.B1(n_3098),
.B2(n_3143),
.Y(n_3357)
);

AND2x4_ASAP7_75t_L g3358 ( 
.A(n_3278),
.B(n_3197),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_3254),
.B(n_3212),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3280),
.Y(n_3360)
);

AO22x1_ASAP7_75t_L g3361 ( 
.A1(n_3265),
.A2(n_3097),
.B1(n_2994),
.B2(n_3113),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3256),
.B(n_3242),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_L g3363 ( 
.A1(n_3247),
.A2(n_3102),
.B(n_3216),
.C(n_3194),
.Y(n_3363)
);

AO221x1_ASAP7_75t_L g3364 ( 
.A1(n_3291),
.A2(n_3137),
.B1(n_2833),
.B2(n_3066),
.C(n_3085),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3290),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3254),
.B(n_3244),
.Y(n_3366)
);

AOI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3334),
.A2(n_3259),
.B1(n_3286),
.B2(n_3278),
.Y(n_3367)
);

XNOR2xp5_ASAP7_75t_L g3368 ( 
.A(n_3361),
.B(n_2915),
.Y(n_3368)
);

XNOR2xp5_ASAP7_75t_L g3369 ( 
.A(n_3315),
.B(n_2835),
.Y(n_3369)
);

XNOR2x1_ASAP7_75t_L g3370 ( 
.A(n_3326),
.B(n_2939),
.Y(n_3370)
);

OAI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3334),
.A2(n_3111),
.B(n_3286),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3329),
.B(n_3304),
.Y(n_3372)
);

OAI21xp33_ASAP7_75t_SL g3373 ( 
.A1(n_3364),
.A2(n_3291),
.B(n_3277),
.Y(n_3373)
);

OR2x6_ASAP7_75t_L g3374 ( 
.A(n_3363),
.B(n_2912),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3351),
.A2(n_3345),
.B1(n_3355),
.B2(n_3353),
.Y(n_3375)
);

INVxp67_ASAP7_75t_L g3376 ( 
.A(n_3320),
.Y(n_3376)
);

OAI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_3351),
.A2(n_3291),
.B1(n_3292),
.B2(n_3266),
.Y(n_3377)
);

OAI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_3314),
.A2(n_3085),
.B1(n_3081),
.B2(n_3105),
.Y(n_3378)
);

AND2x4_ASAP7_75t_L g3379 ( 
.A(n_3353),
.B(n_3286),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_3317),
.B(n_3304),
.Y(n_3380)
);

XOR2x2_ASAP7_75t_L g3381 ( 
.A(n_3355),
.B(n_2886),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3354),
.Y(n_3382)
);

OAI31xp33_ASAP7_75t_SL g3383 ( 
.A1(n_3325),
.A2(n_3292),
.A3(n_3277),
.B(n_3190),
.Y(n_3383)
);

BUFx2_ASAP7_75t_L g3384 ( 
.A(n_3322),
.Y(n_3384)
);

NAND3xp33_ASAP7_75t_L g3385 ( 
.A(n_3356),
.B(n_3293),
.C(n_3279),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3323),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3328),
.Y(n_3387)
);

NOR3xp33_ASAP7_75t_L g3388 ( 
.A(n_3340),
.B(n_2953),
.C(n_2949),
.Y(n_3388)
);

OAI21xp33_ASAP7_75t_L g3389 ( 
.A1(n_3330),
.A2(n_3259),
.B(n_3262),
.Y(n_3389)
);

OAI221xp5_ASAP7_75t_SL g3390 ( 
.A1(n_3357),
.A2(n_3143),
.B1(n_3303),
.B2(n_3270),
.C(n_3262),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3332),
.A2(n_3292),
.B1(n_3299),
.B2(n_3081),
.Y(n_3391)
);

OAI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3357),
.A2(n_3327),
.B(n_3350),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3343),
.Y(n_3393)
);

OAI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3350),
.A2(n_3105),
.B1(n_3153),
.B2(n_3083),
.Y(n_3394)
);

AO22x1_ASAP7_75t_L g3395 ( 
.A1(n_3325),
.A2(n_3022),
.B1(n_2967),
.B2(n_3294),
.Y(n_3395)
);

AOI21xp33_ASAP7_75t_SL g3396 ( 
.A1(n_3358),
.A2(n_2912),
.B(n_2932),
.Y(n_3396)
);

NAND2xp33_ASAP7_75t_SL g3397 ( 
.A(n_3342),
.B(n_2884),
.Y(n_3397)
);

XOR2xp5_ASAP7_75t_L g3398 ( 
.A(n_3324),
.B(n_2933),
.Y(n_3398)
);

AOI21xp33_ASAP7_75t_L g3399 ( 
.A1(n_3339),
.A2(n_3150),
.B(n_3231),
.Y(n_3399)
);

O2A1O1Ixp33_ASAP7_75t_SL g3400 ( 
.A1(n_3362),
.A2(n_2863),
.B(n_3293),
.C(n_2961),
.Y(n_3400)
);

AOI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3358),
.A2(n_3267),
.B1(n_3270),
.B2(n_3299),
.Y(n_3401)
);

AOI321xp33_ASAP7_75t_L g3402 ( 
.A1(n_3375),
.A2(n_3366),
.A3(n_3043),
.B1(n_3312),
.B2(n_3267),
.C(n_3296),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_3388),
.B(n_3333),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3384),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3372),
.Y(n_3405)
);

INVxp67_ASAP7_75t_L g3406 ( 
.A(n_3381),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3387),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3393),
.Y(n_3408)
);

AND2x2_ASAP7_75t_SL g3409 ( 
.A(n_3383),
.B(n_3192),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3373),
.B(n_3290),
.Y(n_3410)
);

OAI221xp5_ASAP7_75t_L g3411 ( 
.A1(n_3371),
.A2(n_3341),
.B1(n_3360),
.B2(n_3344),
.C(n_3346),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3395),
.A2(n_2921),
.B(n_2932),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3374),
.A2(n_3359),
.B1(n_3335),
.B2(n_3316),
.Y(n_3413)
);

OAI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_3374),
.A2(n_3352),
.B1(n_3337),
.B2(n_3338),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3382),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3386),
.B(n_3296),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3380),
.B(n_3256),
.Y(n_3417)
);

AOI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3397),
.A2(n_3299),
.B1(n_3235),
.B2(n_3331),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3376),
.Y(n_3419)
);

AOI32xp33_ASAP7_75t_L g3420 ( 
.A1(n_3377),
.A2(n_3389),
.A3(n_3370),
.B1(n_3378),
.B2(n_3379),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3385),
.Y(n_3421)
);

INVx2_ASAP7_75t_SL g3422 ( 
.A(n_3368),
.Y(n_3422)
);

OAI221xp5_ASAP7_75t_L g3423 ( 
.A1(n_3392),
.A2(n_3302),
.B1(n_3336),
.B2(n_2952),
.C(n_3284),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3367),
.B(n_3287),
.Y(n_3424)
);

AND2x2_ASAP7_75t_L g3425 ( 
.A(n_3379),
.B(n_3237),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3401),
.Y(n_3426)
);

OAI32xp33_ASAP7_75t_L g3427 ( 
.A1(n_3391),
.A2(n_3309),
.A3(n_3298),
.B1(n_3348),
.B2(n_3347),
.Y(n_3427)
);

AO22x2_ASAP7_75t_L g3428 ( 
.A1(n_3398),
.A2(n_3365),
.B1(n_3318),
.B2(n_3319),
.Y(n_3428)
);

NAND2xp33_ASAP7_75t_SL g3429 ( 
.A(n_3396),
.B(n_2989),
.Y(n_3429)
);

OR2x2_ASAP7_75t_L g3430 ( 
.A(n_3390),
.B(n_3313),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3369),
.Y(n_3431)
);

AOI22xp5_ASAP7_75t_L g3432 ( 
.A1(n_3400),
.A2(n_3283),
.B1(n_3281),
.B2(n_3121),
.Y(n_3432)
);

OR2x6_ASAP7_75t_L g3433 ( 
.A(n_3394),
.B(n_2887),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3399),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_3383),
.A2(n_3349),
.B(n_3016),
.C(n_2966),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3384),
.Y(n_3436)
);

OAI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3374),
.A2(n_3106),
.B1(n_3009),
.B2(n_3197),
.Y(n_3437)
);

XNOR2x1_ASAP7_75t_L g3438 ( 
.A(n_3431),
.B(n_2964),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_3404),
.B(n_3321),
.Y(n_3439)
);

NOR3x1_ASAP7_75t_L g3440 ( 
.A(n_3422),
.B(n_3423),
.C(n_3421),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3403),
.B(n_3409),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3406),
.B(n_3281),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3436),
.B(n_3283),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3419),
.B(n_3231),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3407),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3412),
.B(n_2984),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3435),
.A2(n_2887),
.B(n_2975),
.Y(n_3447)
);

NOR2x1_ASAP7_75t_L g3448 ( 
.A(n_3433),
.B(n_2879),
.Y(n_3448)
);

NAND3xp33_ASAP7_75t_L g3449 ( 
.A(n_3420),
.B(n_2936),
.C(n_2658),
.Y(n_3449)
);

AOI211xp5_ASAP7_75t_L g3450 ( 
.A1(n_3429),
.A2(n_2992),
.B(n_2836),
.C(n_2974),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_3402),
.B(n_3258),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3408),
.Y(n_3452)
);

OR2x2_ASAP7_75t_L g3453 ( 
.A(n_3430),
.B(n_3248),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3410),
.A2(n_2985),
.B(n_2956),
.Y(n_3454)
);

AND2x2_ASAP7_75t_L g3455 ( 
.A(n_3433),
.B(n_3130),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3428),
.B(n_3405),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3428),
.B(n_3248),
.Y(n_3457)
);

NOR3x1_ASAP7_75t_L g3458 ( 
.A(n_3411),
.B(n_3214),
.C(n_3025),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_SL g3459 ( 
.A(n_3437),
.B(n_3033),
.Y(n_3459)
);

OR2x2_ASAP7_75t_L g3460 ( 
.A(n_3415),
.B(n_3426),
.Y(n_3460)
);

A2O1A1Ixp33_ASAP7_75t_L g3461 ( 
.A1(n_3413),
.A2(n_3414),
.B(n_3418),
.C(n_3427),
.Y(n_3461)
);

NAND3xp33_ASAP7_75t_SL g3462 ( 
.A(n_3434),
.B(n_2965),
.C(n_2937),
.Y(n_3462)
);

NOR3xp33_ASAP7_75t_L g3463 ( 
.A(n_3449),
.B(n_3424),
.C(n_2469),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3447),
.A2(n_3416),
.B(n_3425),
.Y(n_3464)
);

OA211x2_ASAP7_75t_L g3465 ( 
.A1(n_3446),
.A2(n_3417),
.B(n_2736),
.C(n_3432),
.Y(n_3465)
);

OAI211xp5_ASAP7_75t_SL g3466 ( 
.A1(n_3461),
.A2(n_2718),
.B(n_3026),
.C(n_3243),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_3460),
.Y(n_3467)
);

AOI22xp5_ASAP7_75t_L g3468 ( 
.A1(n_3449),
.A2(n_3159),
.B1(n_3158),
.B2(n_3036),
.Y(n_3468)
);

NOR3xp33_ASAP7_75t_L g3469 ( 
.A(n_3462),
.B(n_3017),
.C(n_2612),
.Y(n_3469)
);

OA22x2_ASAP7_75t_L g3470 ( 
.A1(n_3441),
.A2(n_2999),
.B1(n_3013),
.B2(n_3214),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3438),
.B(n_2742),
.Y(n_3471)
);

OAI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3456),
.A2(n_2560),
.B(n_2659),
.Y(n_3472)
);

NOR3xp33_ASAP7_75t_L g3473 ( 
.A(n_3448),
.B(n_2623),
.C(n_2570),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3442),
.B(n_3099),
.Y(n_3474)
);

NAND4xp75_ASAP7_75t_L g3475 ( 
.A(n_3440),
.B(n_2454),
.C(n_2425),
.D(n_2396),
.Y(n_3475)
);

INVx2_ASAP7_75t_SL g3476 ( 
.A(n_3455),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3439),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3445),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_3452),
.B(n_2742),
.Y(n_3479)
);

AOI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3459),
.A2(n_3036),
.B1(n_3106),
.B2(n_3107),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3451),
.B(n_2521),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_3454),
.A2(n_2999),
.B(n_3115),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3476),
.Y(n_3483)
);

AOI221xp5_ASAP7_75t_L g3484 ( 
.A1(n_3466),
.A2(n_3457),
.B1(n_3459),
.B2(n_3444),
.C(n_3453),
.Y(n_3484)
);

OAI211xp5_ASAP7_75t_SL g3485 ( 
.A1(n_3472),
.A2(n_3450),
.B(n_3443),
.C(n_3458),
.Y(n_3485)
);

AND2x2_ASAP7_75t_L g3486 ( 
.A(n_3471),
.B(n_3450),
.Y(n_3486)
);

OAI21xp33_ASAP7_75t_L g3487 ( 
.A1(n_3470),
.A2(n_2464),
.B(n_2445),
.Y(n_3487)
);

NAND4xp75_ASAP7_75t_L g3488 ( 
.A(n_3465),
.B(n_2454),
.C(n_2436),
.D(n_2404),
.Y(n_3488)
);

AOI221x1_ASAP7_75t_L g3489 ( 
.A1(n_3463),
.A2(n_2872),
.B1(n_2866),
.B2(n_2856),
.C(n_3119),
.Y(n_3489)
);

AO221x1_ASAP7_75t_L g3490 ( 
.A1(n_3477),
.A2(n_2959),
.B1(n_2928),
.B2(n_3008),
.C(n_2918),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3467),
.B(n_3251),
.Y(n_3491)
);

NAND3xp33_ASAP7_75t_L g3492 ( 
.A(n_3469),
.B(n_2433),
.C(n_2310),
.Y(n_3492)
);

O2A1O1Ixp33_ASAP7_75t_L g3493 ( 
.A1(n_3478),
.A2(n_3481),
.B(n_3482),
.C(n_3464),
.Y(n_3493)
);

OAI221xp5_ASAP7_75t_SL g3494 ( 
.A1(n_3480),
.A2(n_3013),
.B1(n_3155),
.B2(n_3151),
.C(n_3127),
.Y(n_3494)
);

AOI211xp5_ASAP7_75t_L g3495 ( 
.A1(n_3479),
.A2(n_2872),
.B(n_2866),
.C(n_2856),
.Y(n_3495)
);

NOR3xp33_ASAP7_75t_L g3496 ( 
.A(n_3475),
.B(n_2512),
.C(n_2528),
.Y(n_3496)
);

AOI31xp33_ASAP7_75t_L g3497 ( 
.A1(n_3468),
.A2(n_3012),
.A3(n_3010),
.B(n_3123),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3474),
.B(n_3251),
.Y(n_3498)
);

INVxp67_ASAP7_75t_L g3499 ( 
.A(n_3483),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3488),
.A2(n_3470),
.B1(n_3473),
.B2(n_3056),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3486),
.B(n_3258),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3484),
.B(n_3125),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3491),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3490),
.Y(n_3504)
);

NOR2x1_ASAP7_75t_L g3505 ( 
.A(n_3485),
.B(n_2389),
.Y(n_3505)
);

AOI22xp5_ASAP7_75t_L g3506 ( 
.A1(n_3487),
.A2(n_2497),
.B1(n_3135),
.B2(n_3120),
.Y(n_3506)
);

AND3x4_ASAP7_75t_L g3507 ( 
.A(n_3496),
.B(n_3012),
.C(n_3010),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3493),
.B(n_3122),
.Y(n_3508)
);

OA22x2_ASAP7_75t_L g3509 ( 
.A1(n_3489),
.A2(n_3498),
.B1(n_3494),
.B2(n_3497),
.Y(n_3509)
);

NOR2x1_ASAP7_75t_L g3510 ( 
.A(n_3492),
.B(n_2412),
.Y(n_3510)
);

NAND4xp75_ASAP7_75t_L g3511 ( 
.A(n_3505),
.B(n_3495),
.C(n_2454),
.D(n_2354),
.Y(n_3511)
);

NAND5xp2_ASAP7_75t_L g3512 ( 
.A(n_3499),
.B(n_2615),
.C(n_2617),
.D(n_2607),
.E(n_2599),
.Y(n_3512)
);

AND2x4_ASAP7_75t_L g3513 ( 
.A(n_3504),
.B(n_3124),
.Y(n_3513)
);

OAI211xp5_ASAP7_75t_L g3514 ( 
.A1(n_3503),
.A2(n_3508),
.B(n_3500),
.C(n_3506),
.Y(n_3514)
);

NOR2x1_ASAP7_75t_L g3515 ( 
.A(n_3507),
.B(n_3501),
.Y(n_3515)
);

NAND5xp2_ASAP7_75t_L g3516 ( 
.A(n_3502),
.B(n_2972),
.C(n_2792),
.D(n_2782),
.E(n_2789),
.Y(n_3516)
);

OR2x2_ASAP7_75t_L g3517 ( 
.A(n_3509),
.B(n_3129),
.Y(n_3517)
);

HB1xp67_ASAP7_75t_L g3518 ( 
.A(n_3510),
.Y(n_3518)
);

NAND3xp33_ASAP7_75t_L g3519 ( 
.A(n_3499),
.B(n_2354),
.C(n_2393),
.Y(n_3519)
);

NAND3xp33_ASAP7_75t_L g3520 ( 
.A(n_3513),
.B(n_2324),
.C(n_2928),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3513),
.Y(n_3521)
);

OA21x2_ASAP7_75t_L g3522 ( 
.A1(n_3514),
.A2(n_2476),
.B(n_2463),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_3517),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3518),
.Y(n_3524)
);

AO22x2_ASAP7_75t_L g3525 ( 
.A1(n_3521),
.A2(n_3511),
.B1(n_3515),
.B2(n_3516),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3525),
.Y(n_3526)
);

HB1xp67_ASAP7_75t_L g3527 ( 
.A(n_3526),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3527),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3528),
.B(n_3523),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3529),
.A2(n_3524),
.B1(n_3522),
.B2(n_3520),
.Y(n_3530)
);

OR2x6_ASAP7_75t_L g3531 ( 
.A(n_3530),
.B(n_3522),
.Y(n_3531)
);

AOI22xp33_ASAP7_75t_L g3532 ( 
.A1(n_3531),
.A2(n_3512),
.B1(n_3519),
.B2(n_2497),
.Y(n_3532)
);


endmodule