module real_aes_16082_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g111 ( .A(n_0), .B(n_112), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_1), .A2(n_31), .B1(n_148), .B2(n_240), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_2), .A2(n_9), .B1(n_545), .B2(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_4), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_5), .A2(n_10), .B1(n_546), .B2(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g107 ( .A(n_6), .B(n_27), .Y(n_107) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_7), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_8), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_11), .B(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_12), .A2(n_97), .B1(n_193), .B2(n_545), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_13), .A2(n_28), .B1(n_563), .B2(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_14), .B(n_163), .Y(n_560) );
OAI21x1_ASAP7_75t_L g143 ( .A1(n_15), .A2(n_46), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_16), .B(n_244), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_17), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_18), .A2(n_35), .B1(n_200), .B2(n_215), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_19), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_20), .A2(n_43), .B1(n_215), .B2(n_545), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_21), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_22), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_23), .B(n_223), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_24), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_25), .B(n_141), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_26), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_29), .A2(n_81), .B1(n_148), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_30), .A2(n_34), .B1(n_148), .B2(n_548), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_32), .A2(n_49), .B1(n_545), .B2(n_600), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_33), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_36), .B(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_37), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_38), .B(n_163), .Y(n_211) );
INVx2_ASAP7_75t_L g119 ( .A(n_39), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_40), .B(n_196), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_41), .Y(n_859) );
BUFx3_ASAP7_75t_L g106 ( .A(n_42), .Y(n_106) );
INVx1_ASAP7_75t_L g836 ( .A(n_42), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_44), .B(n_182), .Y(n_246) );
XOR2x2_ASAP7_75t_L g130 ( .A(n_45), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g274 ( .A(n_47), .B(n_182), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_48), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_50), .B(n_223), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_51), .B(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_52), .A2(n_68), .B1(n_200), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_53), .A2(n_71), .B1(n_148), .B2(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_54), .B(n_304), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_55), .A2(n_152), .B(n_161), .C(n_267), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_56), .A2(n_94), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g144 ( .A(n_57), .Y(n_144) );
AND2x4_ASAP7_75t_L g166 ( .A(n_58), .B(n_167), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_59), .A2(n_60), .B1(n_215), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_61), .B(n_141), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_62), .B(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_63), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_64), .B(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g167 ( .A(n_65), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_66), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_67), .B(n_141), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_69), .B(n_148), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g239 ( .A(n_70), .B(n_196), .C(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_72), .B(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_73), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_74), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_75), .B(n_163), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_76), .B(n_157), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_77), .A2(n_93), .B1(n_161), .B2(n_215), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_78), .A2(n_130), .B1(n_838), .B2(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_78), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_79), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g574 ( .A(n_80), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_82), .A2(n_88), .B1(n_222), .B2(n_223), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_83), .B(n_163), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_84), .Y(n_854) );
NAND2xp33_ASAP7_75t_SL g180 ( .A(n_85), .B(n_151), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_86), .B(n_194), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_87), .B(n_141), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_89), .Y(n_585) );
INVx1_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_90), .B(n_835), .Y(n_834) );
NAND2xp33_ASAP7_75t_L g564 ( .A(n_91), .B(n_163), .Y(n_564) );
NAND2xp33_ASAP7_75t_L g150 ( .A(n_92), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_95), .B(n_182), .Y(n_306) );
NAND3xp33_ASAP7_75t_L g176 ( .A(n_96), .B(n_151), .C(n_175), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_98), .B(n_148), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_99), .B(n_223), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_113), .B(n_858), .Y(n_100) );
CKINVDCx6p67_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
BUFx12f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_SL g861 ( .A(n_103), .Y(n_861) );
OR2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_108), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g846 ( .A(n_105), .B(n_129), .Y(n_846) );
NOR2x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_107), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND3x2_ASAP7_75t_L g856 ( .A(n_109), .B(n_122), .C(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_853), .Y(n_113) );
OAI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_123), .B(n_830), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
BUFx12f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x6_ASAP7_75t_SL g117 ( .A(n_118), .B(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g831 ( .A(n_119), .B(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_119), .B(n_845), .Y(n_844) );
INVx3_ASAP7_75t_L g851 ( .A(n_119), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x6_ASAP7_75t_SL g833 ( .A(n_122), .B(n_834), .Y(n_833) );
AOI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_519), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g519 ( .A(n_126), .B(n_520), .Y(n_519) );
INVx8_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx12f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g838 ( .A(n_130), .Y(n_838) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_451), .Y(n_131) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_326), .C(n_366), .D(n_415), .Y(n_132) );
NOR2xp67_ASAP7_75t_L g133 ( .A(n_134), .B(n_275), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_185), .B1(n_247), .B2(n_256), .Y(n_134) );
INVx1_ASAP7_75t_L g447 ( .A(n_135), .Y(n_447) );
INVx1_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_136), .B(n_294), .Y(n_363) );
AND2x2_ASAP7_75t_L g394 ( .A(n_136), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_168), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_137), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g318 ( .A(n_137), .Y(n_318) );
AND2x2_ASAP7_75t_L g493 ( .A(n_137), .B(n_361), .Y(n_493) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx2_ASAP7_75t_L g258 ( .A(n_138), .Y(n_258) );
AND2x2_ASAP7_75t_L g346 ( .A(n_138), .B(n_308), .Y(n_346) );
AND2x2_ASAP7_75t_L g390 ( .A(n_138), .B(n_295), .Y(n_390) );
OR2x2_ASAP7_75t_L g408 ( .A(n_138), .B(n_409), .Y(n_408) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g312 ( .A(n_139), .B(n_295), .Y(n_312) );
BUFx2_ASAP7_75t_L g369 ( .A(n_139), .Y(n_369) );
OR2x2_ASAP7_75t_L g377 ( .A(n_139), .B(n_335), .Y(n_377) );
INVx1_ASAP7_75t_L g432 ( .A(n_139), .Y(n_432) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
INVx2_ASAP7_75t_L g572 ( .A(n_141), .Y(n_572) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_SL g164 ( .A(n_142), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g171 ( .A(n_142), .Y(n_171) );
INVx2_ASAP7_75t_L g207 ( .A(n_142), .Y(n_207) );
BUFx3_ASAP7_75t_L g528 ( .A(n_142), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_142), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g556 ( .A(n_142), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_142), .B(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_142), .B(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_155), .B(n_164), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_150), .B(n_152), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_148), .A2(n_215), .B1(n_272), .B2(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g546 ( .A(n_148), .Y(n_546) );
INVx4_ASAP7_75t_L g548 ( .A(n_148), .Y(n_548) );
INVx1_ASAP7_75t_L g600 ( .A(n_148), .Y(n_600) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_149), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
INVx1_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g224 ( .A(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_149), .Y(n_240) );
INVx2_ASAP7_75t_L g269 ( .A(n_149), .Y(n_269) );
INVx2_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
INVx1_ASAP7_75t_L g563 ( .A(n_151), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_178), .B(n_180), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_152), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_152), .A2(n_299), .B(n_300), .Y(n_298) );
BUFx4f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g159 ( .A(n_154), .Y(n_159) );
INVx1_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
BUFx8_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B1(n_160), .B2(n_162), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_157), .A2(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_163), .A2(n_174), .B(n_176), .Y(n_173) );
INVx1_ASAP7_75t_L g244 ( .A(n_163), .Y(n_244) );
INVx3_ASAP7_75t_L g545 ( .A(n_163), .Y(n_545) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_165), .A2(n_173), .B(n_177), .Y(n_172) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_191), .B(n_197), .Y(n_190) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_165), .A2(n_209), .B(n_212), .Y(n_208) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_165), .A2(n_237), .B(n_241), .Y(n_236) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_165), .A2(n_298), .B(n_301), .Y(n_297) );
BUFx10_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx10_ASAP7_75t_L g231 ( .A(n_166), .Y(n_231) );
INVx1_ASAP7_75t_L g535 ( .A(n_166), .Y(n_535) );
AND2x2_ASAP7_75t_L g259 ( .A(n_168), .B(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g371 ( .A(n_168), .B(n_348), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_168), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g409 ( .A(n_169), .Y(n_409) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_169), .Y(n_414) );
AND2x2_ASAP7_75t_L g431 ( .A(n_169), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g321 ( .A(n_170), .B(n_261), .Y(n_321) );
INVx1_ASAP7_75t_L g335 ( .A(n_170), .Y(n_335) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_181), .Y(n_170) );
INVx1_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
INVx1_ASAP7_75t_L g533 ( .A(n_175), .Y(n_533) );
INVx1_ASAP7_75t_SL g549 ( .A(n_175), .Y(n_549) );
INVx1_ASAP7_75t_L g591 ( .A(n_179), .Y(n_591) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g189 ( .A(n_183), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_183), .B(n_603), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_183), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g230 ( .A(n_184), .Y(n_230) );
INVx2_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
NAND2x1_ASAP7_75t_L g185 ( .A(n_186), .B(n_202), .Y(n_185) );
AND2x4_ASAP7_75t_L g496 ( .A(n_186), .B(n_424), .Y(n_496) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_187), .Y(n_255) );
BUFx3_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
INVx1_ASAP7_75t_L g356 ( .A(n_187), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_187), .B(n_205), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_187), .B(n_235), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_187), .Y(n_387) );
AND2x2_ASAP7_75t_L g419 ( .A(n_187), .B(n_284), .Y(n_419) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_201), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_189), .A2(n_190), .B(n_201), .Y(n_285) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_189), .A2(n_297), .B(n_306), .Y(n_296) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_189), .A2(n_297), .B(n_306), .Y(n_324) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_196), .A2(n_213), .B(n_214), .Y(n_212) );
INVx6_ASAP7_75t_L g225 ( .A(n_196), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g558 ( .A1(n_196), .A2(n_548), .B(n_559), .C(n_560), .Y(n_558) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g328 ( .A(n_204), .B(n_314), .Y(n_328) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g354 ( .A(n_206), .B(n_341), .Y(n_354) );
AND2x2_ASAP7_75t_L g383 ( .A(n_206), .B(n_219), .Y(n_383) );
OR2x2_ASAP7_75t_L g479 ( .A(n_206), .B(n_219), .Y(n_479) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_216), .Y(n_206) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_207), .A2(n_236), .B(n_246), .Y(n_235) );
OAI21x1_ASAP7_75t_L g253 ( .A1(n_207), .A2(n_208), .B(n_216), .Y(n_253) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_207), .A2(n_236), .B(n_246), .Y(n_284) );
INVx2_ASAP7_75t_L g222 ( .A(n_215), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g358 ( .A(n_217), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g507 ( .A(n_217), .Y(n_507) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
OR2x2_ASAP7_75t_L g441 ( .A(n_218), .B(n_251), .Y(n_441) );
INVx1_ASAP7_75t_L g463 ( .A(n_218), .Y(n_463) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_235), .Y(n_218) );
AND2x2_ASAP7_75t_L g279 ( .A(n_219), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g314 ( .A(n_219), .B(n_284), .Y(n_314) );
INVx1_ASAP7_75t_L g341 ( .A(n_219), .Y(n_341) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_219), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_219), .B(n_235), .Y(n_428) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_230), .A3(n_231), .B(n_232), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_225), .B1(n_226), .B2(n_228), .Y(n_220) );
INVx1_ASAP7_75t_L g582 ( .A(n_223), .Y(n_582) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_225), .A2(n_530), .B1(n_532), .B2(n_533), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_225), .A2(n_544), .B1(n_547), .B2(n_549), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_225), .A2(n_562), .B(n_564), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_225), .A2(n_228), .B1(n_570), .B2(n_571), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_225), .A2(n_549), .B1(n_581), .B2(n_583), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_225), .A2(n_228), .B1(n_590), .B2(n_592), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_225), .A2(n_228), .B1(n_599), .B2(n_601), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_225), .A2(n_228), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g593 ( .A(n_227), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_228), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g305 ( .A(n_229), .Y(n_305) );
INVx2_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_230), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_SL g584 ( .A(n_230), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
AO31x2_ASAP7_75t_L g568 ( .A1(n_231), .A2(n_569), .A3(n_572), .B(n_573), .Y(n_568) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_231), .A2(n_542), .A3(n_580), .B(n_584), .Y(n_579) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_231), .A2(n_528), .A3(n_589), .B(n_594), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
BUFx2_ASAP7_75t_L g542 ( .A(n_234), .Y(n_542) );
AND2x2_ASAP7_75t_L g365 ( .A(n_235), .B(n_285), .Y(n_365) );
INVx2_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
AOI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .Y(n_241) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR3x1_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .C(n_254), .Y(n_248) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_251), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g313 ( .A(n_251), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g364 ( .A(n_251), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g404 ( .A(n_251), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_251), .B(n_427), .Y(n_459) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_252), .B(n_340), .Y(n_400) );
AND2x2_ASAP7_75t_L g424 ( .A(n_252), .B(n_284), .Y(n_424) );
BUFx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g280 ( .A(n_253), .Y(n_280) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g435 ( .A(n_255), .B(n_314), .Y(n_435) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_258), .B(n_321), .Y(n_500) );
AND2x4_ASAP7_75t_L g492 ( .A(n_259), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_259), .B(n_312), .Y(n_506) );
INVx2_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
INVx2_ASAP7_75t_L g396 ( .A(n_260), .Y(n_396) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g380 ( .A(n_261), .Y(n_380) );
AOI21x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_274), .Y(n_261) );
NOR2xp67_ASAP7_75t_SL g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g597 ( .A(n_263), .Y(n_597) );
INVx1_ASAP7_75t_L g550 ( .A(n_264), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_270), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_SL g531 ( .A(n_269), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_315), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_291), .B1(n_309), .B2(n_313), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_286), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g343 ( .A(n_279), .B(n_290), .Y(n_343) );
AND2x2_ASAP7_75t_L g503 ( .A(n_279), .B(n_384), .Y(n_503) );
BUFx2_ASAP7_75t_L g374 ( .A(n_280), .Y(n_374) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g373 ( .A(n_283), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g288 ( .A(n_284), .Y(n_288) );
INVx1_ASAP7_75t_L g340 ( .A(n_284), .Y(n_340) );
INVx1_ASAP7_75t_L g465 ( .A(n_285), .Y(n_465) );
AOI31xp33_ASAP7_75t_L g483 ( .A1(n_286), .A2(n_484), .A3(n_485), .B(n_486), .Y(n_483) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_288), .B(n_383), .Y(n_482) );
INVx2_ASAP7_75t_L g510 ( .A(n_288), .Y(n_510) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_289), .Y(n_325) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g338 ( .A(n_290), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_290), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g468 ( .A(n_290), .B(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_307), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g379 ( .A(n_295), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g348 ( .A(n_296), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_305), .Y(n_301) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_311), .Y(n_332) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx1_ASAP7_75t_L g352 ( .A(n_312), .Y(n_352) );
AND2x2_ASAP7_75t_L g413 ( .A(n_312), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g469 ( .A(n_312), .B(n_396), .Y(n_469) );
OAI21xp5_ASAP7_75t_L g385 ( .A1(n_313), .A2(n_386), .B(n_388), .Y(n_385) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_325), .Y(n_315) );
NAND3x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .C(n_322), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g487 ( .A(n_318), .B(n_407), .Y(n_487) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2x1_ASAP7_75t_SL g440 ( .A(n_320), .B(n_352), .Y(n_440) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g360 ( .A(n_321), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_322), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_322), .B(n_431), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_322), .B(n_431), .Y(n_504) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g407 ( .A(n_324), .B(n_380), .Y(n_407) );
AND2x2_ASAP7_75t_L g327 ( .A(n_325), .B(n_328), .Y(n_327) );
AOI221x1_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B1(n_336), .B2(n_345), .C(n_349), .Y(n_326) );
AOI32xp33_ASAP7_75t_L g508 ( .A1(n_328), .A2(n_509), .A3(n_514), .B1(n_515), .B2(n_517), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_333), .B(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g347 ( .A(n_335), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_335), .Y(n_351) );
OR2x2_ASAP7_75t_L g464 ( .A(n_335), .B(n_465), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_342), .C(n_344), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g386 ( .A(n_339), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g403 ( .A(n_339), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_342), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_438) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g516 ( .A(n_346), .Y(n_516) );
INVx2_ASAP7_75t_L g361 ( .A(n_348), .Y(n_361) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B(n_357), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g485 ( .A(n_354), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_355), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_364), .Y(n_357) );
AND2x4_ASAP7_75t_L g454 ( .A(n_360), .B(n_369), .Y(n_454) );
INVx1_ASAP7_75t_L g513 ( .A(n_361), .Y(n_513) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g392 ( .A(n_365), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_365), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_365), .B(n_393), .Y(n_484) );
AOI211x1_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_373), .B(n_375), .C(n_401), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR3x2_ASAP7_75t_L g476 ( .A(n_369), .B(n_371), .C(n_372), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_370), .A2(n_392), .B1(n_394), .B2(n_397), .Y(n_391) );
NOR2x1p5_ASAP7_75t_SL g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_371), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx2_ASAP7_75t_L g393 ( .A(n_374), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_381), .B(n_385), .C(n_391), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_383), .B(n_387), .Y(n_398) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_383), .B(n_490), .Y(n_498) );
OAI32xp33_ASAP7_75t_L g473 ( .A1(n_384), .A2(n_429), .A3(n_474), .B1(n_476), .B2(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g490 ( .A(n_384), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_384), .B(n_404), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_387), .B(n_421), .Y(n_456) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g434 ( .A(n_393), .B(n_419), .Y(n_434) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g443 ( .A(n_396), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g411 ( .A(n_399), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B1(n_410), .B2(n_412), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g449 ( .A(n_406), .Y(n_449) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g430 ( .A(n_407), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_407), .B(n_414), .Y(n_518) );
INVx1_ASAP7_75t_SL g444 ( .A(n_408), .Y(n_444) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_438), .C(n_445), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_429), .B(n_433), .Y(n_416) );
NOR2xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_422), .Y(n_417) );
INVxp67_ASAP7_75t_L g450 ( .A(n_418), .Y(n_450) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .C(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g437 ( .A(n_431), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g446 ( .A(n_434), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_439), .A2(n_490), .B1(n_491), .B2(n_494), .C(n_495), .Y(n_489) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI32xp33_ASAP7_75t_L g445 ( .A1(n_442), .A2(n_446), .A3(n_447), .B1(n_448), .B2(n_450), .Y(n_445) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_448), .A2(n_458), .B1(n_459), .B2(n_460), .C(n_466), .Y(n_457) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_470), .C(n_488), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B(n_457), .Y(n_452) );
AOI211x1_ASAP7_75t_L g470 ( .A1(n_453), .A2(n_471), .B(n_473), .C(n_480), .Y(n_470) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2x1_ASAP7_75t_SL g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g472 ( .A(n_463), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AO21x1_ASAP7_75t_L g480 ( .A1(n_469), .A2(n_481), .B(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g514 ( .A(n_485), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_501), .Y(n_488) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_497), .B(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_505), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g511 ( .A(n_510), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND4xp75_ASAP7_75t_L g520 ( .A(n_521), .B(n_670), .C(n_746), .D(n_798), .Y(n_520) );
AND3x1_ASAP7_75t_L g521 ( .A(n_522), .B(n_643), .C(n_656), .Y(n_521) );
AOI221x1_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_575), .B1(n_604), .B2(n_608), .C(n_620), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_523), .A2(n_644), .B(n_646), .C(n_647), .Y(n_643) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_538), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g607 ( .A(n_527), .Y(n_607) );
BUFx2_ASAP7_75t_L g625 ( .A(n_527), .Y(n_625) );
OR2x2_ASAP7_75t_L g667 ( .A(n_527), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g674 ( .A(n_527), .B(n_541), .Y(n_674) );
AND2x4_ASAP7_75t_L g709 ( .A(n_527), .B(n_540), .Y(n_709) );
OR2x2_ASAP7_75t_L g752 ( .A(n_527), .B(n_568), .Y(n_752) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_529), .A3(n_534), .B(n_536), .Y(n_527) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_534), .A2(n_597), .A3(n_598), .B(n_602), .Y(n_596) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g565 ( .A(n_535), .Y(n_565) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_553), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_540), .B(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_540), .Y(n_639) );
INVx2_ASAP7_75t_L g666 ( .A(n_540), .Y(n_666) );
INVx3_ASAP7_75t_L g679 ( .A(n_540), .Y(n_679) );
AND2x2_ASAP7_75t_L g797 ( .A(n_540), .B(n_626), .Y(n_797) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g606 ( .A(n_541), .B(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g662 ( .A(n_541), .Y(n_662) );
AO31x2_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .A3(n_550), .B(n_551), .Y(n_541) );
AO31x2_ASAP7_75t_L g613 ( .A1(n_550), .A2(n_597), .A3(n_614), .B(n_617), .Y(n_613) );
INVxp67_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g682 ( .A(n_554), .Y(n_682) );
INVx1_ASAP7_75t_L g809 ( .A(n_554), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_567), .Y(n_554) );
AND2x2_ASAP7_75t_L g605 ( .A(n_555), .B(n_568), .Y(n_605) );
INVx1_ASAP7_75t_L g668 ( .A(n_555), .Y(n_668) );
OAI21x1_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_566), .Y(n_555) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_556), .A2(n_557), .B(n_566), .Y(n_627) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_565), .Y(n_557) );
INVx2_ASAP7_75t_L g623 ( .A(n_567), .Y(n_623) );
AND2x2_ASAP7_75t_L g675 ( .A(n_567), .B(n_626), .Y(n_675) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_568), .Y(n_697) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_577), .A2(n_669), .B1(n_673), .B2(n_676), .Y(n_672) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_586), .Y(n_577) );
INVx1_ASAP7_75t_L g690 ( .A(n_578), .Y(n_690) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g610 ( .A(n_579), .B(n_588), .Y(n_610) );
AND2x2_ASAP7_75t_L g641 ( .A(n_579), .B(n_596), .Y(n_641) );
INVx4_ASAP7_75t_SL g652 ( .A(n_579), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_579), .B(n_686), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_579), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g723 ( .A(n_587), .B(n_701), .Y(n_723) );
OR2x2_ASAP7_75t_L g756 ( .A(n_587), .B(n_738), .Y(n_756) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_596), .Y(n_587) );
INVx2_ASAP7_75t_L g630 ( .A(n_588), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_588), .Y(n_635) );
AND2x2_ASAP7_75t_L g642 ( .A(n_588), .B(n_612), .Y(n_642) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_588), .Y(n_658) );
INVx1_ASAP7_75t_L g686 ( .A(n_588), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_588), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g619 ( .A(n_596), .Y(n_619) );
AND2x4_ASAP7_75t_L g629 ( .A(n_596), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g655 ( .A(n_596), .Y(n_655) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_596), .Y(n_732) );
INVx1_ASAP7_75t_L g825 ( .A(n_596), .Y(n_825) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_605), .B(n_678), .Y(n_745) );
AND2x2_ASAP7_75t_L g758 ( .A(n_605), .B(n_674), .Y(n_758) );
AND2x2_ASAP7_75t_L g828 ( .A(n_605), .B(n_679), .Y(n_828) );
AND2x4_ASAP7_75t_L g663 ( .A(n_607), .B(n_626), .Y(n_663) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g730 ( .A(n_610), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g744 ( .A(n_610), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_610), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g646 ( .A(n_611), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_611), .B(n_684), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_611), .A2(n_741), .B(n_744), .C(n_745), .Y(n_740) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_619), .Y(n_611) );
AND2x2_ASAP7_75t_L g711 ( .A(n_612), .B(n_652), .Y(n_711) );
INVx3_ASAP7_75t_L g738 ( .A(n_612), .Y(n_738) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g633 ( .A(n_613), .Y(n_633) );
AND2x4_ASAP7_75t_L g659 ( .A(n_613), .B(n_619), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_619), .B(n_652), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_628), .B1(n_636), .B2(n_640), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g777 ( .A(n_622), .Y(n_777) );
AND2x4_ASAP7_75t_L g688 ( .A(n_623), .B(n_668), .Y(n_688) );
INVx1_ASAP7_75t_L g708 ( .A(n_623), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_625), .A2(n_681), .B1(n_691), .B2(n_693), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_625), .B(n_682), .Y(n_739) );
NAND2x1_ASAP7_75t_L g796 ( .A(n_625), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g811 ( .A(n_625), .Y(n_811) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g750 ( .A(n_627), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
AND2x2_ASAP7_75t_L g669 ( .A(n_629), .B(n_651), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_629), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g710 ( .A(n_629), .B(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_629), .Y(n_784) );
NAND2x1p5_ASAP7_75t_L g791 ( .A(n_629), .B(n_692), .Y(n_791) );
AND2x4_ASAP7_75t_L g814 ( .A(n_629), .B(n_742), .Y(n_814) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx3_ASAP7_75t_L g692 ( .A(n_632), .Y(n_692) );
AND2x2_ASAP7_75t_L g704 ( .A(n_632), .B(n_697), .Y(n_704) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g654 ( .A(n_633), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g702 ( .A(n_633), .Y(n_702) );
INVx1_ASAP7_75t_L g645 ( .A(n_634), .Y(n_645) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g802 ( .A(n_635), .B(n_652), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g728 ( .A(n_637), .B(n_709), .Y(n_728) );
INVx2_ASAP7_75t_L g769 ( .A(n_637), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_637), .B(n_663), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_638), .B(n_688), .Y(n_818) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_641), .B(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g713 ( .A(n_641), .B(n_658), .Y(n_713) );
INVx1_ASAP7_75t_L g805 ( .A(n_641), .Y(n_805) );
AND2x2_ASAP7_75t_L g804 ( .A(n_642), .B(n_731), .Y(n_804) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g775 ( .A1(n_646), .A2(n_776), .B1(n_778), .B2(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g684 ( .A(n_652), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g720 ( .A(n_652), .Y(n_720) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_652), .Y(n_726) );
INVx2_ASAP7_75t_L g743 ( .A(n_652), .Y(n_743) );
OR2x2_ASAP7_75t_L g764 ( .A(n_652), .B(n_727), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_652), .B(n_722), .Y(n_774) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g741 ( .A(n_654), .B(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_654), .Y(n_795) );
INVx1_ASAP7_75t_L g722 ( .A(n_655), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .B(n_664), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_659), .B(n_690), .Y(n_689) );
INVx3_ASAP7_75t_L g727 ( .A(n_659), .Y(n_727) );
AND2x2_ASAP7_75t_L g801 ( .A(n_659), .B(n_802), .Y(n_801) );
AOI211x1_ASAP7_75t_SL g729 ( .A1(n_660), .A2(n_730), .B(n_733), .C(n_740), .Y(n_729) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g786 ( .A(n_662), .B(n_663), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_663), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g779 ( .A(n_663), .Y(n_779) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_669), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g694 ( .A(n_666), .Y(n_694) );
NOR2x1p5_ASAP7_75t_L g751 ( .A(n_666), .B(n_752), .Y(n_751) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_667), .B(n_696), .Y(n_695) );
NOR2xp67_ASAP7_75t_SL g768 ( .A(n_667), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g829 ( .A(n_669), .B(n_737), .Y(n_829) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_714), .Y(n_670) );
NAND3xp33_ASAP7_75t_SL g671 ( .A(n_672), .B(n_680), .C(n_698), .Y(n_671) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_674), .Y(n_705) );
AND2x2_ASAP7_75t_L g712 ( .A(n_674), .B(n_708), .Y(n_712) );
AND2x4_ASAP7_75t_SL g826 ( .A(n_674), .B(n_688), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_675), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_677), .A2(n_719), .B1(n_791), .B2(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_L g808 ( .A(n_679), .B(n_809), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_687), .B2(n_689), .Y(n_681) );
NAND2x1_ASAP7_75t_L g757 ( .A(n_684), .B(n_737), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_684), .B(n_731), .Y(n_767) );
INVx1_ASAP7_75t_L g794 ( .A(n_684), .Y(n_794) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g812 ( .A1(n_687), .A2(n_813), .B(n_816), .Y(n_812) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_688), .A2(n_700), .B(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g773 ( .A(n_692), .Y(n_773) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g717 ( .A(n_695), .Y(n_717) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_705), .B1(n_706), .B2(n_710), .C1(n_712), .C2(n_713), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g733 ( .A1(n_700), .A2(n_734), .B(n_739), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_701), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g815 ( .A(n_701), .Y(n_815) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_702), .Y(n_821) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
AND2x2_ASAP7_75t_L g785 ( .A(n_707), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g778 ( .A(n_708), .B(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_729), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B1(n_724), .B2(n_728), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g735 ( .A(n_721), .Y(n_735) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx4_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g763 ( .A(n_738), .B(n_755), .Y(n_763) );
OR2x2_ASAP7_75t_L g823 ( .A(n_738), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND5xp2_ASAP7_75t_L g799 ( .A(n_744), .B(n_791), .C(n_800), .D(n_803), .E(n_805), .Y(n_799) );
NOR2x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_782), .Y(n_746) );
NAND2xp67_ASAP7_75t_SL g747 ( .A(n_748), .B(n_765), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_753), .B1(n_758), .B2(n_759), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND3xp33_ASAP7_75t_SL g753 ( .A(n_754), .B(n_756), .C(n_757), .Y(n_753) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g788 ( .A(n_757), .Y(n_788) );
NAND3xp33_ASAP7_75t_SL g759 ( .A(n_760), .B(n_763), .C(n_764), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g781 ( .A(n_762), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_SL g793 ( .A1(n_763), .A2(n_794), .B(n_795), .C(n_796), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_770), .B2(n_771), .C(n_775), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_772), .B(n_820), .Y(n_819) );
OR2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g789 ( .A(n_776), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_L g792 ( .A(n_786), .Y(n_792) );
AOI211xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B(n_790), .C(n_793), .Y(n_787) );
AOI211x1_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_806), .B(n_812), .C(n_827), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2x1p5_ASAP7_75t_L g807 ( .A(n_808), .B(n_810), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .B1(n_822), .B2(n_826), .Y(n_816) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_837), .B(n_840), .Y(n_830) );
INVx5_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_836), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_847), .B2(n_852), .Y(n_840) );
INVx6_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx10_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx4_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
CKINVDCx11_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
BUFx6f_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NOR2x1_ASAP7_75t_R g853 ( .A(n_854), .B(n_855), .Y(n_853) );
INVx4_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_SL g858 ( .A(n_859), .B(n_860), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
endmodule