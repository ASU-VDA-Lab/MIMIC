module fake_aes_10922_n_23 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_23);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_23;
wire n_20;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_1), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_3), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_4), .B(n_7), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_2), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_13), .Y(n_15) );
AOI22xp33_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_12), .B1(n_10), .B2(n_11), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NOR3xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_15), .C(n_8), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_20), .B(n_0), .Y(n_21) );
INVxp67_ASAP7_75t_SL g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
endmodule