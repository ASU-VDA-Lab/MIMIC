module fake_jpeg_2514_n_30 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx24_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_9),
.B(n_11),
.C(n_3),
.Y(n_14)
);

A2O1A1Ixp33_ASAP7_75t_SL g18 ( 
.A1(n_14),
.A2(n_10),
.B(n_11),
.C(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_12),
.B1(n_10),
.B2(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_10),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_22),
.A2(n_20),
.B1(n_14),
.B2(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

NAND4xp25_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_21),
.C(n_12),
.D(n_7),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_7),
.B(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_26),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_4),
.B1(n_5),
.B2(n_28),
.Y(n_30)
);


endmodule