module fake_jpeg_13820_n_347 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_18),
.A2(n_9),
.B(n_2),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_19),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_68),
.Y(n_108)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_71),
.B(n_79),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_83),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_35),
.C(n_33),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_74),
.B(n_6),
.C(n_7),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_31),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_39),
.B1(n_33),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_85),
.A2(n_107),
.B1(n_112),
.B2(n_40),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_88),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_43),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_96),
.A2(n_2),
.B(n_6),
.C(n_7),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_41),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_18),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_41),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_27),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_106),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_39),
.B1(n_33),
.B2(n_26),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_48),
.Y(n_111)
);

NAND2x1_ASAP7_75t_SL g150 ( 
.A(n_111),
.B(n_17),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_33),
.B1(n_39),
.B2(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_23),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_25),
.Y(n_129)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_117),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_19),
.B1(n_38),
.B2(n_40),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_152),
.B1(n_78),
.B2(n_72),
.Y(n_158)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_0),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_128),
.A2(n_134),
.B1(n_144),
.B2(n_108),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_132),
.Y(n_155)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_130),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_37),
.B1(n_38),
.B2(n_19),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_30),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_39),
.B1(n_37),
.B2(n_34),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_36),
.B(n_38),
.C(n_21),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_99),
.B(n_114),
.Y(n_181)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_138),
.Y(n_173)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_74),
.A2(n_25),
.B1(n_36),
.B2(n_31),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_80),
.B(n_93),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_0),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_72),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_75),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_143),
.Y(n_180)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_36),
.B1(n_21),
.B2(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_21),
.B1(n_3),
.B2(n_5),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_108),
.B1(n_99),
.B2(n_81),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_99),
.B1(n_92),
.B2(n_89),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_10),
.C(n_11),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_89),
.A2(n_95),
.B1(n_73),
.B2(n_78),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_84),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_8),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_95),
.B1(n_93),
.B2(n_102),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_156),
.A2(n_185),
.B1(n_181),
.B2(n_183),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_164),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_166),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_87),
.B(n_75),
.C(n_103),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_179),
.B(n_141),
.C(n_149),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_91),
.B1(n_72),
.B2(n_78),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_167),
.B(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_84),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_176),
.B1(n_177),
.B2(n_143),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_150),
.B(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_189),
.C(n_145),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_108),
.B1(n_104),
.B2(n_103),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_129),
.B(n_87),
.CI(n_104),
.CON(n_179),
.SN(n_179)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_181),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_117),
.B1(n_116),
.B2(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_102),
.B1(n_81),
.B2(n_114),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_171),
.A2(n_140),
.B1(n_151),
.B2(n_153),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_192),
.A2(n_194),
.B1(n_206),
.B2(n_162),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_190),
.B1(n_155),
.B2(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_126),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_127),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_119),
.C(n_138),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_213),
.C(n_178),
.Y(n_233)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_214),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_122),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_130),
.B1(n_144),
.B2(n_148),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_223),
.B1(n_181),
.B2(n_173),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_208),
.B(n_186),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_123),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_136),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_160),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_238),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_218),
.A2(n_178),
.B1(n_181),
.B2(n_185),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_225),
.A2(n_226),
.B1(n_242),
.B2(n_246),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_233),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_221),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_234),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_205),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_193),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_197),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_249),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_156),
.B1(n_162),
.B2(n_159),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_195),
.B1(n_222),
.B2(n_207),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_189),
.B1(n_173),
.B2(n_182),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_191),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_182),
.B1(n_183),
.B2(n_170),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_220),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_270),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_236),
.A2(n_202),
.B(n_222),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_267),
.B(n_242),
.Y(n_274)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_195),
.B(n_194),
.C(n_196),
.D(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_257),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_213),
.C(n_192),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.C(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_228),
.C(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_199),
.C(n_198),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_183),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_201),
.B1(n_216),
.B2(n_211),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_170),
.C(n_172),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_273),
.C(n_250),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_238),
.B(n_225),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_172),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_272),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_214),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_121),
.C(n_14),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_286),
.B(n_13),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_231),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_259),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_237),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_235),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_262),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_284),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_287),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_241),
.B(n_239),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_241),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_239),
.C(n_227),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_258),
.C(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_245),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_248),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_300),
.C(n_303),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_252),
.B1(n_271),
.B2(n_270),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_257),
.B1(n_254),
.B2(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_248),
.C(n_247),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_277),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_13),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_280),
.C(n_283),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_285),
.B(n_275),
.C(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_14),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_15),
.Y(n_311)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_297),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_317),
.Y(n_325)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_294),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_274),
.B1(n_286),
.B2(n_281),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_318),
.A2(n_313),
.B1(n_312),
.B2(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_300),
.C(n_292),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_296),
.C(n_278),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_303),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_308),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_313),
.B1(n_312),
.B2(n_287),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_329),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_299),
.B(n_307),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_331),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_298),
.B(n_315),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_321),
.B(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_304),
.B(n_291),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_338),
.B(n_334),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_339),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_340),
.B(n_341),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_323),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_336),
.C(n_332),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_331),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_342),
.B1(n_333),
.B2(n_16),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_16),
.Y(n_347)
);


endmodule