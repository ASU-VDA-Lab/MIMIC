module fake_jpeg_1343_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_19),
.B(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_50),
.A2(n_46),
.B1(n_37),
.B2(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_46),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_71),
.Y(n_79)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_37),
.B1(n_51),
.B2(n_35),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_18),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_15),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_59),
.B1(n_38),
.B2(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_81),
.B1(n_87),
.B2(n_84),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_59),
.B1(n_38),
.B2(n_2),
.Y(n_81)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_13),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_5),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_12),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_76),
.B1(n_72),
.B2(n_8),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_27),
.B(n_29),
.C(n_28),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_16),
.B(n_32),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_109),
.B(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_117),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_99),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_116),
.C(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_7),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_115),
.B(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.C(n_109),
.Y(n_123)
);

OAI31xp33_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_120),
.A3(n_114),
.B(n_11),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_124),
.B(n_9),
.C(n_10),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_8),
.C(n_9),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_34),
.Y(n_129)
);


endmodule