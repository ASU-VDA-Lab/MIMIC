module fake_jpeg_30982_n_528 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_15),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_14),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_59),
.B(n_93),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_14),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_65),
.B(n_74),
.Y(n_139)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_66),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_26),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_77),
.B(n_89),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_79),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_41),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_85),
.Y(n_171)
);

CKINVDCx10_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_86),
.Y(n_129)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_26),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_91),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_34),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx2_ASAP7_75t_R g93 ( 
.A(n_17),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_23),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_95),
.B(n_106),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_28),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_28),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_30),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_93),
.B(n_49),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_59),
.A2(n_19),
.B(n_12),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_142),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_45),
.B1(n_19),
.B2(n_52),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_137),
.A2(n_144),
.B1(n_146),
.B2(n_73),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_77),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_100),
.A2(n_45),
.B1(n_19),
.B2(n_52),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_45),
.B1(n_54),
.B2(n_43),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g149 ( 
.A(n_83),
.Y(n_149)
);

CKINVDCx12_ASAP7_75t_R g213 ( 
.A(n_149),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_29),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_31),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g223 ( 
.A(n_153),
.Y(n_223)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_66),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_132),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_190),
.Y(n_245)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_197),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_64),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_182),
.B(n_183),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_108),
.C(n_104),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_117),
.A2(n_96),
.B1(n_56),
.B2(n_78),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g255 ( 
.A1(n_187),
.A2(n_191),
.B1(n_214),
.B2(n_120),
.Y(n_255)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_112),
.A2(n_67),
.B1(n_70),
.B2(n_63),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_164),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_196),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_113),
.B(n_139),
.Y(n_196)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_103),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_97),
.B1(n_62),
.B2(n_72),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_139),
.B(n_17),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_39),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_218),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_207),
.Y(n_233)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_76),
.B1(n_102),
.B2(n_39),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_225),
.B1(n_138),
.B2(n_129),
.Y(n_239)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_133),
.A2(n_71),
.B1(n_105),
.B2(n_92),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_33),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_110),
.B(n_32),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_110),
.B(n_38),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_144),
.A2(n_32),
.B1(n_51),
.B2(n_50),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_151),
.Y(n_237)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_222),
.Y(n_253)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_116),
.A2(n_43),
.B1(n_38),
.B2(n_94),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_237),
.A2(n_185),
.B1(n_188),
.B2(n_204),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_162),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_246),
.B(n_256),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_198),
.A2(n_146),
.B(n_137),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_254),
.A2(n_138),
.B(n_130),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_255),
.A2(n_178),
.B1(n_210),
.B2(n_208),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_181),
.B(n_140),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_218),
.B(n_140),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_260),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_162),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_141),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_177),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_175),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_290),
.C(n_264),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_267),
.B(n_270),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_238),
.A2(n_198),
.B1(n_191),
.B2(n_187),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_274),
.B1(n_295),
.B2(n_233),
.Y(n_301)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_173),
.Y(n_270)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_261),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_275),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_250),
.B1(n_229),
.B2(n_255),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_273),
.A2(n_298),
.B1(n_255),
.B2(n_207),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_238),
.A2(n_214),
.B1(n_145),
.B2(n_141),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_173),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_292),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_234),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_281),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_223),
.Y(n_281)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_213),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_294),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_205),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_287),
.Y(n_319)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_226),
.B(n_184),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_288),
.A2(n_253),
.B(n_232),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_226),
.B(n_259),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_248),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_291),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_293),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_222),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_246),
.A2(n_145),
.B1(n_116),
.B2(n_118),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_233),
.B(n_180),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_258),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_301),
.A2(n_284),
.B1(n_292),
.B2(n_274),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_276),
.A2(n_229),
.B1(n_255),
.B2(n_233),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_320),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_276),
.A2(n_293),
.B1(n_288),
.B2(n_269),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_308),
.A2(n_322),
.B(n_247),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_243),
.B(n_253),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_309),
.A2(n_314),
.B(n_312),
.Y(n_356)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_253),
.B(n_244),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_316),
.A2(n_323),
.B1(n_295),
.B2(n_268),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

AOI32xp33_ASAP7_75t_L g321 ( 
.A1(n_281),
.A2(n_193),
.A3(n_257),
.B1(n_161),
.B2(n_168),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_219),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_289),
.A2(n_220),
.B1(n_263),
.B2(n_172),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_241),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_266),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_231),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_327),
.Y(n_345)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_336),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_303),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_332),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_357),
.B1(n_318),
.B2(n_300),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_287),
.B1(n_285),
.B2(n_283),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_334),
.A2(n_346),
.B1(n_309),
.B2(n_345),
.Y(n_367)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_325),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_358),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_310),
.B(n_291),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_340),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_282),
.B1(n_286),
.B2(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_359),
.Y(n_372)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_323),
.A2(n_252),
.B1(n_251),
.B2(n_277),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_311),
.B(n_51),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_347),
.B(n_25),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_348),
.A2(n_349),
.B(n_353),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_329),
.A2(n_247),
.B(n_265),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_320),
.A2(n_265),
.B(n_176),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_212),
.B(n_216),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_354),
.Y(n_364)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_355),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_314),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_313),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_302),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_301),
.A2(n_134),
.B1(n_189),
.B2(n_147),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_342),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_306),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_365),
.B(n_385),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_367),
.B(n_374),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_327),
.C(n_319),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_386),
.C(n_388),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_319),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_369),
.B(n_368),
.Y(n_393)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_376),
.C(n_381),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_333),
.A2(n_334),
.B1(n_337),
.B2(n_339),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_373),
.A2(n_387),
.B1(n_344),
.B2(n_338),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_340),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_332),
.B(n_313),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_391),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_380),
.A2(n_342),
.B1(n_360),
.B2(n_354),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_SL g381 ( 
.A(n_347),
.B(n_315),
.C(n_326),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_359),
.B(n_307),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_328),
.Y(n_384)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_384),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_315),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_324),
.C(n_300),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_318),
.C(n_299),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_299),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_349),
.B(n_50),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_416),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_357),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_394),
.B(n_406),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_341),
.Y(n_395)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_395),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_379),
.A2(n_348),
.B(n_364),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_372),
.A2(n_341),
.B1(n_342),
.B2(n_346),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_399),
.A2(n_400),
.B1(n_414),
.B2(n_419),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_389),
.Y(n_401)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_364),
.A2(n_342),
.B(n_353),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_404),
.A2(n_417),
.B(n_352),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_355),
.C(n_335),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_410),
.C(n_411),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_385),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_383),
.Y(n_408)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_373),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_409),
.B(n_415),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_363),
.C(n_386),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_351),
.C(n_350),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_350),
.Y(n_412)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_412),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_413),
.A2(n_230),
.B1(n_236),
.B2(n_211),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_359),
.B1(n_307),
.B2(n_352),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_366),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_379),
.B(n_271),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_371),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_420),
.A2(n_224),
.B1(n_174),
.B2(n_160),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_372),
.C(n_390),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_426),
.C(n_429),
.Y(n_448)
);

FAx1_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_381),
.CI(n_361),
.CON(n_424),
.SN(n_424)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_433),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_R g425 ( 
.A(n_408),
.B(n_361),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_425),
.A2(n_430),
.B(n_126),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_390),
.C(n_371),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_248),
.C(n_240),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_240),
.C(n_236),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_443),
.C(n_412),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_227),
.Y(n_433)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_413),
.A2(n_230),
.B1(n_192),
.B2(n_36),
.Y(n_436)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_416),
.B(n_199),
.Y(n_439)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_143),
.C(n_121),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_442),
.A2(n_428),
.B1(n_402),
.B2(n_427),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_444),
.B(n_454),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_441),
.Y(n_446)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_397),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_449),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_425),
.A2(n_403),
.B1(n_395),
.B2(n_418),
.Y(n_450)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_393),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_431),
.Y(n_473)
);

AOI321xp33_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_394),
.A3(n_404),
.B1(n_411),
.B2(n_399),
.C(n_407),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_452),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g455 ( 
.A(n_424),
.B(n_396),
.C(n_417),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_455),
.A2(n_432),
.B1(n_29),
.B2(n_31),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_435),
.A2(n_219),
.B(n_174),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_460),
.B(n_439),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_440),
.B(n_126),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_429),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_435),
.A2(n_114),
.B1(n_118),
.B2(n_36),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_25),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_467),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_437),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_466),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_457),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_440),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_426),
.C(n_423),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_468),
.B(n_478),
.C(n_479),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_443),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_477),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_473),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_42),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_80),
.C(n_79),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_82),
.C(n_84),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_476),
.A2(n_453),
.B(n_455),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_481),
.B(n_486),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_475),
.A2(n_460),
.B1(n_445),
.B2(n_461),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_482),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_462),
.B1(n_452),
.B2(n_454),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_485),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_465),
.B(n_468),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_451),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_492),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_488),
.A2(n_480),
.B1(n_484),
.B2(n_482),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_114),
.B1(n_42),
.B2(n_69),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_479),
.B(n_0),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_148),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_1),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_495),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_473),
.C(n_478),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_500),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_494),
.B(n_467),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_498),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_491),
.A2(n_148),
.B(n_3),
.Y(n_498)
);

AOI321xp33_ASAP7_75t_L g500 ( 
.A1(n_494),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_504),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_493),
.B1(n_490),
.B2(n_9),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_4),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_506),
.A2(n_6),
.B(n_8),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_513),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_511),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_490),
.B1(n_9),
.B2(n_10),
.Y(n_513)
);

OAI211xp5_ASAP7_75t_L g514 ( 
.A1(n_499),
.A2(n_8),
.B(n_10),
.C(n_501),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_514),
.A2(n_506),
.B(n_502),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_518),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_503),
.B(n_505),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_504),
.C(n_8),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_514),
.Y(n_520)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_515),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_508),
.B(n_512),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_523),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_524),
.B(n_522),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_517),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_527),
.Y(n_528)
);


endmodule