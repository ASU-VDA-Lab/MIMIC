module fake_jpeg_27259_n_93 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_24),
.B(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_45),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_55),
.B(n_56),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_4),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_12),
.B(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_6),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_76),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_64),
.B(n_48),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_77),
.B1(n_68),
.B2(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_40),
.B1(n_34),
.B2(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_69),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_66),
.B(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_80),
.B(n_81),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_72),
.A3(n_46),
.B1(n_33),
.B2(n_43),
.C1(n_44),
.C2(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_23),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_72),
.B(n_38),
.Y(n_93)
);


endmodule