module real_jpeg_25501_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_61),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_38),
.B1(n_42),
.B2(n_61),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_79),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_38),
.B1(n_42),
.B2(n_79),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_3),
.B(n_52),
.C(n_54),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_99),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_77),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_99),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_3),
.B(n_38),
.C(n_85),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_37),
.B(n_153),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_58),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_38),
.B1(n_42),
.B2(n_58),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_38),
.B1(n_42),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_38),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_14),
.A2(n_36),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_128),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_105),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_72),
.B2(n_73),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_48),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

AOI32xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.A3(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_23),
.A2(n_24),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_24),
.B(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_93)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_37),
.A2(n_41),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_37),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_37),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_42),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_39),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_42),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_45),
.A2(n_167),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_65),
.C(n_68),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_49),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_59),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_52),
.B1(n_84),
.B2(n_85),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_52),
.B(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_60),
.B(n_77),
.Y(n_138)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_91),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_87),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_87),
.B(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_83),
.B(n_99),
.Y(n_173)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_113),
.B1(n_115),
.B2(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_101),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_102),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_99),
.B(n_100),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_155),
.Y(n_178)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_107),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_116),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_114),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_111),
.A2(n_114),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_119),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.Y(n_119)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_142),
.B(n_189),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_139),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.C(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_183),
.B(n_188),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_163),
.B(n_182),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_157),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_157),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_171),
.B(n_181),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_169),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_180),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_187),
.Y(n_188)
);


endmodule