module real_jpeg_11148_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_3),
.A2(n_19),
.B1(n_20),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_33),
.B(n_35),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_19),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_4),
.B(n_19),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_49),
.B1(n_54),
.B2(n_86),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_11),
.A2(n_19),
.B1(n_20),
.B2(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_42),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_65),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_58),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_58),
.Y(n_65)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_16),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_31),
.CI(n_43),
.CON(n_16),
.SN(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_18),
.A2(n_22),
.B1(n_25),
.B2(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_23),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_19),
.A2(n_20),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_22),
.A2(n_25),
.B1(n_60),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_25),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_26),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_26),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_37),
.Y(n_38)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_62),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_54),
.B1(n_71),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_51),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_62),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_63),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_61),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_94),
.B(n_98),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_83),
.B(n_93),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_82),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_77),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_88),
.B(n_92),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);


endmodule