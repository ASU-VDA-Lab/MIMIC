module fake_jpeg_21480_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_15),
.B1(n_20),
.B2(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_16),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_48),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_31),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_14),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_54),
.B1(n_40),
.B2(n_17),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_66),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_35),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_36),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_36),
.B(n_30),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_40),
.B(n_18),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_14),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_18),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_49),
.C(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_87),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_63),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_67),
.B(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_70),
.B1(n_65),
.B2(n_64),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_26),
.C(n_25),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_55),
.C(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_77),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_96),
.B(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_67),
.B(n_13),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_61),
.B1(n_59),
.B2(n_86),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_61),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_75),
.C(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_83),
.B1(n_79),
.B2(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_25),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_0),
.C(n_2),
.Y(n_114)
);

OAI321xp33_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_89),
.A3(n_93),
.B1(n_96),
.B2(n_90),
.C(n_88),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_114),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_101),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_110),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_123),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_107),
.A3(n_105),
.B1(n_5),
.B2(n_8),
.C1(n_10),
.C2(n_11),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_4),
.C(n_8),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_121),
.C(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_0),
.Y(n_129)
);


endmodule