module fake_netlist_5_1241_n_938 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_938);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_938;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_615;
wire n_469;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_928;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_525;
wire n_493;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_929;
wire n_804;
wire n_867;
wire n_186;
wire n_537;
wire n_902;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_570;
wire n_457;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_185;
wire n_243;
wire n_183;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_632;
wire n_489;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_917;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_911;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_679;
wire n_407;
wire n_527;
wire n_513;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_832;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_70),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_59),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_54),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_73),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_90),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_48),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_76),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_120),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_49),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_109),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_45),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_65),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_53),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_97),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_27),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_79),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_177),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_169),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_87),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_135),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_118),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_71),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_46),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_117),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_61),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_62),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_108),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_18),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_43),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_107),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_153),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_72),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_114),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_35),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_75),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_128),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_174),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_91),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_121),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_4),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_181),
.B(n_0),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_0),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_181),
.B(n_197),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_212),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_176),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_1),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_1),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_178),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_206),
.B(n_2),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_2),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_244),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_185),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_3),
.Y(n_287)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_180),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_179),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_210),
.B(n_3),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_210),
.B(n_5),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_183),
.B(n_175),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_210),
.B(n_5),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_186),
.B(n_6),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_191),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_182),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_212),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_241),
.B(n_6),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_222),
.B(n_7),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g306 ( 
.A(n_187),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_279),
.A2(n_211),
.B1(n_201),
.B2(n_213),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_250),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_223),
.B1(n_245),
.B2(n_231),
.Y(n_309)
);

NAND3x1_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_237),
.C(n_236),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_220),
.B1(n_188),
.B2(n_221),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_258),
.A2(n_238),
.B1(n_252),
.B2(n_251),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_240),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_258),
.A2(n_247),
.B1(n_249),
.B2(n_248),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_215),
.B1(n_246),
.B2(n_242),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_287),
.A2(n_254),
.B1(n_234),
.B2(n_233),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_232),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_292),
.A2(n_230),
.B1(n_229),
.B2(n_228),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_276),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_227),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_288),
.A2(n_224),
.B1(n_219),
.B2(n_216),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_288),
.A2(n_287),
.B1(n_259),
.B2(n_275),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_189),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_190),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_271),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_284),
.B(n_193),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_293),
.A2(n_214),
.B1(n_208),
.B2(n_207),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_203),
.B1(n_202),
.B2(n_199),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_204),
.B1(n_196),
.B2(n_195),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_194),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_293),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_283),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_265),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_10),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

AO22x2_ASAP7_75t_L g342 ( 
.A1(n_295),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_342)
);

BUFx6f_ASAP7_75t_SL g343 ( 
.A(n_268),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_31),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_L g346 ( 
.A1(n_297),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_17),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_R g349 ( 
.A1(n_269),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_273),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_304),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_291),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_265),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_259),
.A2(n_275),
.B1(n_265),
.B2(n_288),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_290),
.B(n_32),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_304),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_271),
.B(n_268),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_272),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_290),
.B(n_33),
.Y(n_361)
);

OA22x2_ASAP7_75t_L g362 ( 
.A1(n_269),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_271),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_312),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_268),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_314),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_307),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_324),
.B(n_294),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_272),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_268),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_257),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_345),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_307),
.B(n_272),
.Y(n_387)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_351),
.B(n_272),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_356),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_325),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_294),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_342),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_311),
.B(n_257),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_299),
.Y(n_406)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_339),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_318),
.B(n_294),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_257),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_299),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_357),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_359),
.B(n_281),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_359),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_309),
.B(n_334),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_355),
.B(n_294),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_313),
.B(n_281),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_315),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_346),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_349),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_330),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_358),
.B(n_299),
.Y(n_432)
);

AND2x6_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_281),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_312),
.Y(n_435)
);

BUFx6f_ASAP7_75t_SL g436 ( 
.A(n_341),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_365),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_282),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_282),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_282),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_377),
.A2(n_282),
.B(n_256),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_365),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_383),
.B(n_286),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_286),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_429),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_306),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_390),
.B(n_298),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_430),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_431),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_298),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

NAND2x1p5_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_298),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_403),
.B(n_298),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_364),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_378),
.B(n_301),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_375),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_386),
.B(n_301),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_366),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_399),
.A2(n_305),
.B1(n_301),
.B2(n_296),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_363),
.B(n_301),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_410),
.B(n_306),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_368),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_305),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_306),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_430),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_433),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_385),
.B(n_363),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_374),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_411),
.B(n_305),
.Y(n_480)
);

AND2x2_ASAP7_75t_SL g481 ( 
.A(n_388),
.B(n_283),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_388),
.B(n_305),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_283),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_256),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_256),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_392),
.B(n_402),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_380),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_414),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_426),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_408),
.A2(n_422),
.B(n_404),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_296),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_270),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_433),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_418),
.B(n_270),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_270),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_399),
.A2(n_296),
.B1(n_300),
.B2(n_303),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_410),
.B(n_37),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_277),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_394),
.B(n_38),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_277),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_277),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_396),
.B(n_416),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_406),
.B(n_266),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_416),
.B(n_280),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_413),
.B(n_296),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_421),
.A2(n_303),
.B(n_300),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_399),
.B(n_296),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_296),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_400),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_432),
.B(n_266),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_417),
.B(n_280),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_417),
.B(n_280),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_511),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_481),
.B(n_425),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_508),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_447),
.B(n_381),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_401),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_465),
.Y(n_529)
);

BUFx8_ASAP7_75t_L g530 ( 
.A(n_508),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_384),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_371),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_447),
.B(n_425),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_407),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_520),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_260),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_458),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_518),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_510),
.B(n_436),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_468),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_450),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_437),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_521),
.Y(n_549)
);

NAND2x1p5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_428),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_458),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_437),
.Y(n_552)
);

BUFx8_ASAP7_75t_SL g553 ( 
.A(n_468),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_452),
.B(n_39),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_445),
.B(n_407),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_515),
.B(n_436),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_521),
.B(n_387),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_296),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_452),
.B(n_40),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_484),
.B(n_439),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_514),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_466),
.B(n_41),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_437),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_285),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_466),
.B(n_42),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_454),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_471),
.B(n_285),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_515),
.B(n_424),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_454),
.B(n_47),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_450),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_471),
.B(n_285),
.Y(n_574)
);

OR2x6_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_424),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_476),
.Y(n_576)
);

NOR2x1_ASAP7_75t_L g577 ( 
.A(n_477),
.B(n_300),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_454),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_488),
.B(n_303),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_454),
.B(n_50),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_505),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

NOR2x1_ASAP7_75t_L g584 ( 
.A(n_477),
.B(n_267),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_477),
.B(n_494),
.Y(n_585)
);

BUFx8_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_570),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_557),
.A2(n_481),
.B1(n_472),
.B2(n_512),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_579),
.Y(n_590)
);

BUFx4_ASAP7_75t_SL g591 ( 
.A(n_561),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_530),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_555),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_536),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_538),
.Y(n_595)
);

BUFx2_ASAP7_75t_SL g596 ( 
.A(n_536),
.Y(n_596)
);

BUFx6f_ASAP7_75t_SL g597 ( 
.A(n_575),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_523),
.B(n_481),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_529),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_478),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_525),
.B(n_456),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

INVxp67_ASAP7_75t_SL g604 ( 
.A(n_536),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

INVx3_ASAP7_75t_SL g606 ( 
.A(n_556),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_548),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_548),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_546),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_548),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_564),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_547),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_SL g615 ( 
.A1(n_575),
.A2(n_445),
.B1(n_492),
.B2(n_453),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_585),
.Y(n_616)
);

CKINVDCx14_ASAP7_75t_R g617 ( 
.A(n_535),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_585),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_549),
.B(n_478),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_552),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_522),
.Y(n_621)
);

BUFx12f_ASAP7_75t_L g622 ( 
.A(n_556),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_526),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_499),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_552),
.Y(n_625)
);

BUFx2_ASAP7_75t_SL g626 ( 
.A(n_544),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_531),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_537),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_543),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_531),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_553),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_552),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_556),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_563),
.B(n_494),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_582),
.B(n_502),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_537),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_527),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_589),
.A2(n_524),
.B1(n_493),
.B2(n_575),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_619),
.A2(n_524),
.B1(n_501),
.B2(n_464),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_SL g642 ( 
.A1(n_617),
.A2(n_505),
.B1(n_527),
.B2(n_566),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_621),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_586),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_602),
.A2(n_583),
.B1(n_502),
.B2(n_482),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_602),
.A2(n_502),
.B1(n_482),
.B2(n_505),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_590),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_600),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_593),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_624),
.A2(n_493),
.B(n_560),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_632),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_599),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_591),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_601),
.A2(n_501),
.B1(n_464),
.B2(n_545),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_603),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_595),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_617),
.A2(n_545),
.B1(n_562),
.B2(n_566),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_623),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_622),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_607),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_607),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_621),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_607),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_627),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_607),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_637),
.A2(n_562),
.B1(n_554),
.B2(n_559),
.Y(n_667)
);

BUFx2_ASAP7_75t_SL g668 ( 
.A(n_592),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_597),
.A2(n_559),
.B1(n_554),
.B2(n_581),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_614),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_586),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_627),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_630),
.Y(n_673)
);

INVx6_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_630),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_632),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_634),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_629),
.B(n_638),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_588),
.A2(n_490),
.B1(n_456),
.B2(n_571),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_598),
.A2(n_490),
.B1(n_581),
.B2(n_571),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_637),
.A2(n_528),
.B1(n_560),
.B2(n_488),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_597),
.A2(n_443),
.B1(n_468),
.B2(n_516),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_607),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_605),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_598),
.A2(n_441),
.B1(n_454),
.B2(n_499),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_637),
.B(n_500),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_605),
.A2(n_441),
.B1(n_500),
.B2(n_528),
.Y(n_689)
);

OAI22x1_ASAP7_75t_SL g690 ( 
.A1(n_592),
.A2(n_518),
.B1(n_463),
.B2(n_459),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_597),
.A2(n_468),
.B1(n_480),
.B2(n_507),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_648),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_657),
.B(n_639),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_650),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_653),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_678),
.B(n_506),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_647),
.A2(n_615),
.B1(n_608),
.B2(n_468),
.Y(n_698)
);

BUFx4f_ASAP7_75t_SL g699 ( 
.A(n_660),
.Y(n_699)
);

BUFx2_ASAP7_75t_L g700 ( 
.A(n_659),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_669),
.A2(n_611),
.B1(n_608),
.B2(n_626),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_643),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_L g703 ( 
.A1(n_667),
.A2(n_611),
.B1(n_610),
.B2(n_448),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_649),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_685),
.Y(n_705)
);

OAI222xp33_ASAP7_75t_L g706 ( 
.A1(n_669),
.A2(n_448),
.B1(n_463),
.B2(n_509),
.C1(n_572),
.C2(n_446),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_656),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_658),
.A2(n_681),
.B1(n_640),
.B2(n_642),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_640),
.A2(n_476),
.B1(n_446),
.B2(n_442),
.Y(n_709)
);

BUFx12f_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_644),
.A2(n_587),
.B1(n_448),
.B2(n_613),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_670),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_674),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_658),
.A2(n_606),
.B1(n_613),
.B2(n_448),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_691),
.A2(n_517),
.B(n_507),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_672),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_SL g718 ( 
.A1(n_644),
.A2(n_668),
.B1(n_645),
.B2(n_674),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_690),
.Y(n_719)
);

INVx5_ASAP7_75t_SL g720 ( 
.A(n_661),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_646),
.A2(n_606),
.B1(n_613),
.B2(n_448),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_677),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_691),
.A2(n_476),
.B1(n_442),
.B2(n_504),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_673),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_676),
.B(n_587),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_675),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_SL g728 ( 
.A1(n_683),
.A2(n_506),
.B(n_504),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_679),
.A2(n_613),
.B1(n_563),
.B2(n_497),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_689),
.A2(n_469),
.B1(n_474),
.B2(n_513),
.Y(n_730)
);

INVx3_ASAP7_75t_SL g731 ( 
.A(n_644),
.Y(n_731)
);

CKINVDCx11_ASAP7_75t_R g732 ( 
.A(n_652),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_688),
.A2(n_469),
.B1(n_474),
.B2(n_513),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_665),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_688),
.A2(n_470),
.B1(n_489),
.B2(n_498),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_674),
.A2(n_671),
.B1(n_641),
.B2(n_680),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_683),
.A2(n_470),
.B1(n_489),
.B2(n_498),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_682),
.A2(n_503),
.B1(n_460),
.B2(n_462),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_662),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_686),
.A2(n_613),
.B1(n_569),
.B2(n_574),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_641),
.A2(n_574),
.B1(n_569),
.B2(n_558),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_682),
.B(n_487),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_SL g744 ( 
.A1(n_655),
.A2(n_534),
.B(n_495),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_651),
.B(n_449),
.C(n_519),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_651),
.A2(n_503),
.B1(n_460),
.B2(n_487),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_655),
.A2(n_475),
.B1(n_479),
.B2(n_485),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_684),
.A2(n_475),
.B1(n_479),
.B2(n_485),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_684),
.A2(n_618),
.B1(n_616),
.B2(n_596),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_708),
.A2(n_494),
.B1(n_573),
.B2(n_577),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_708),
.A2(n_618),
.B1(n_616),
.B2(n_596),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_697),
.B(n_662),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_695),
.B(n_662),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_736),
.A2(n_467),
.B1(n_558),
.B2(n_551),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_696),
.Y(n_755)
);

OAI222xp33_ASAP7_75t_L g756 ( 
.A1(n_714),
.A2(n_635),
.B1(n_631),
.B2(n_628),
.C1(n_580),
.C2(n_633),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_703),
.A2(n_577),
.B1(n_568),
.B2(n_578),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_698),
.A2(n_568),
.B1(n_578),
.B2(n_565),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_712),
.B(n_705),
.Y(n_759)
);

AOI221xp5_ASAP7_75t_L g760 ( 
.A1(n_728),
.A2(n_580),
.B1(n_483),
.B2(n_461),
.C(n_635),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_721),
.A2(n_616),
.B1(n_618),
.B2(n_564),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_SL g762 ( 
.A(n_731),
.B(n_565),
.Y(n_762)
);

AOI222xp33_ASAP7_75t_L g763 ( 
.A1(n_715),
.A2(n_564),
.B1(n_604),
.B2(n_578),
.C1(n_568),
.C2(n_565),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_719),
.A2(n_564),
.B1(n_455),
.B2(n_567),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_719),
.A2(n_455),
.B1(n_576),
.B2(n_631),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_711),
.B(n_666),
.C(n_664),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_718),
.A2(n_636),
.B1(n_576),
.B2(n_625),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_702),
.B(n_664),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_700),
.B(n_694),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_709),
.B1(n_737),
.B2(n_724),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_723),
.A2(n_636),
.B1(n_625),
.B2(n_633),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_743),
.A2(n_628),
.B1(n_635),
.B2(n_631),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_740),
.A2(n_666),
.B1(n_664),
.B2(n_594),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_740),
.A2(n_666),
.B1(n_612),
.B2(n_609),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_729),
.A2(n_455),
.B1(n_584),
.B2(n_594),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_699),
.A2(n_612),
.B1(n_609),
.B2(n_636),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_692),
.A2(n_620),
.B1(n_594),
.B2(n_609),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_704),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_730),
.A2(n_733),
.B1(n_744),
.B2(n_747),
.C(n_735),
.Y(n_779)
);

OAI222xp33_ASAP7_75t_L g780 ( 
.A1(n_749),
.A2(n_620),
.B1(n_584),
.B2(n_542),
.C1(n_440),
.C2(n_451),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_707),
.A2(n_713),
.B1(n_717),
.B2(n_727),
.Y(n_781)
);

AOI222xp33_ASAP7_75t_L g782 ( 
.A1(n_706),
.A2(n_473),
.B1(n_260),
.B2(n_267),
.C1(n_261),
.C2(n_262),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_748),
.B(n_612),
.C(n_609),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_710),
.A2(n_620),
.B1(n_612),
.B2(n_609),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_726),
.A2(n_612),
.B1(n_440),
.B2(n_542),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_741),
.A2(n_264),
.B1(n_261),
.B2(n_267),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_734),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_732),
.A2(n_440),
.B1(n_457),
.B2(n_267),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_716),
.B(n_52),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_741),
.A2(n_457),
.B1(n_267),
.B2(n_264),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_742),
.B(n_55),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_738),
.A2(n_457),
.B1(n_267),
.B2(n_264),
.Y(n_792)
);

OA21x2_ASAP7_75t_L g793 ( 
.A1(n_745),
.A2(n_457),
.B(n_267),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_457),
.B1(n_264),
.B2(n_263),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_759),
.B(n_725),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_778),
.B(n_787),
.Y(n_796)
);

OAI221xp5_ASAP7_75t_SL g797 ( 
.A1(n_751),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.C(n_60),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_754),
.B(n_739),
.C(n_693),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_770),
.A2(n_720),
.B1(n_722),
.B2(n_693),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_725),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_752),
.B(n_725),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_779),
.A2(n_766),
.B1(n_782),
.B2(n_750),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_755),
.B(n_725),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_753),
.B(n_725),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_774),
.B(n_725),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_768),
.B(n_722),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_773),
.B(n_720),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_781),
.B(n_720),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_781),
.B(n_64),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_772),
.B(n_66),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_763),
.B(n_260),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_772),
.B(n_68),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_L g813 ( 
.A(n_791),
.B(n_69),
.C(n_77),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_767),
.B(n_771),
.C(n_776),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_SL g815 ( 
.A1(n_758),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.C(n_82),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_789),
.B(n_84),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_754),
.A2(n_264),
.B1(n_263),
.B2(n_262),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_773),
.B(n_85),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_SL g819 ( 
.A1(n_761),
.A2(n_86),
.B(n_88),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_793),
.B(n_260),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_793),
.B(n_260),
.Y(n_821)
);

NAND3xp33_ASAP7_75t_L g822 ( 
.A(n_765),
.B(n_264),
.C(n_263),
.Y(n_822)
);

OAI22xp5_ASAP7_75t_L g823 ( 
.A1(n_757),
.A2(n_788),
.B1(n_764),
.B2(n_784),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_777),
.B(n_785),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_777),
.B(n_89),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_796),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_815),
.B(n_756),
.C(n_783),
.Y(n_827)
);

NAND4xp75_ASAP7_75t_L g828 ( 
.A(n_809),
.B(n_790),
.C(n_793),
.D(n_794),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_813),
.B(n_814),
.C(n_799),
.Y(n_829)
);

NOR2x1_ASAP7_75t_L g830 ( 
.A(n_803),
.B(n_780),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_796),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_800),
.B(n_786),
.Y(n_833)
);

NAND4xp75_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_760),
.C(n_762),
.D(n_94),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_802),
.B(n_798),
.C(n_824),
.Y(n_835)
);

NAND4xp75_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_92),
.C(n_93),
.D(n_96),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_801),
.B(n_775),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_797),
.B(n_792),
.C(n_264),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_804),
.Y(n_839)
);

INVx2_ASAP7_75t_SL g840 ( 
.A(n_806),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_801),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_L g842 ( 
.A(n_819),
.B(n_98),
.C(n_100),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_808),
.B(n_263),
.C(n_262),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_835),
.B(n_818),
.Y(n_844)
);

NAND4xp75_ASAP7_75t_L g845 ( 
.A(n_830),
.B(n_811),
.C(n_807),
.D(n_805),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_841),
.B(n_805),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_826),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_831),
.Y(n_848)
);

NOR2x1_ASAP7_75t_L g849 ( 
.A(n_839),
.B(n_822),
.Y(n_849)
);

NAND4xp75_ASAP7_75t_SL g850 ( 
.A(n_837),
.B(n_807),
.C(n_821),
.D(n_820),
.Y(n_850)
);

NAND4xp75_ASAP7_75t_SL g851 ( 
.A(n_829),
.B(n_821),
.C(n_820),
.D(n_823),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_840),
.Y(n_852)
);

NAND4xp75_ASAP7_75t_L g853 ( 
.A(n_833),
.B(n_825),
.C(n_810),
.D(n_812),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_842),
.A2(n_817),
.B1(n_816),
.B2(n_263),
.Y(n_854)
);

NAND4xp75_ASAP7_75t_L g855 ( 
.A(n_833),
.B(n_101),
.C(n_102),
.D(n_103),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_832),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_843),
.B(n_104),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_828),
.Y(n_858)
);

XNOR2xp5_ASAP7_75t_L g859 ( 
.A(n_853),
.B(n_842),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_858),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_847),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_844),
.B(n_834),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_856),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_846),
.B(n_827),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_856),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_852),
.B(n_836),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_861),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_862),
.B(n_844),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_863),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_860),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_865),
.Y(n_871)
);

AOI22x1_ASAP7_75t_L g872 ( 
.A1(n_859),
.A2(n_857),
.B1(n_851),
.B2(n_846),
.Y(n_872)
);

XNOR2xp5_ASAP7_75t_L g873 ( 
.A(n_864),
.B(n_845),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_862),
.A2(n_866),
.B1(n_860),
.B2(n_854),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_861),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_870),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_875),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_867),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_870),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_873),
.Y(n_880)
);

AOI322xp5_ASAP7_75t_L g881 ( 
.A1(n_868),
.A2(n_849),
.A3(n_827),
.B1(n_848),
.B2(n_852),
.C1(n_850),
.C2(n_838),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_880),
.A2(n_868),
.B1(n_874),
.B2(n_872),
.Y(n_882)
);

AOI31xp33_ASAP7_75t_L g883 ( 
.A1(n_879),
.A2(n_871),
.A3(n_857),
.B(n_869),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_877),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_878),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_882),
.A2(n_880),
.B1(n_876),
.B2(n_881),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_885),
.A2(n_876),
.B1(n_869),
.B2(n_855),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_884),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_883),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_886),
.A2(n_263),
.B1(n_262),
.B2(n_261),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_888),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_889),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_887),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_886),
.A2(n_263),
.B1(n_262),
.B2(n_261),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_889),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_888),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_896),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_892),
.B(n_895),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_891),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_893),
.B(n_105),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_890),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_894),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_896),
.Y(n_903)
);

AND4x1_ASAP7_75t_L g904 ( 
.A(n_900),
.B(n_106),
.C(n_110),
.D(n_111),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_899),
.B(n_112),
.C(n_115),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_898),
.Y(n_906)
);

NOR2xp67_ASAP7_75t_L g907 ( 
.A(n_897),
.B(n_119),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_903),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_908)
);

AND4x1_ASAP7_75t_L g909 ( 
.A(n_901),
.B(n_122),
.C(n_123),
.D(n_124),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_906),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_907),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_909),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_908),
.Y(n_913)
);

XOR2xp5_ASAP7_75t_L g914 ( 
.A(n_904),
.B(n_902),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_905),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_906),
.A2(n_902),
.B1(n_262),
.B2(n_261),
.Y(n_916)
);

AOI211xp5_ASAP7_75t_SL g917 ( 
.A1(n_911),
.A2(n_127),
.B(n_129),
.C(n_130),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_SL g918 ( 
.A1(n_914),
.A2(n_261),
.B1(n_260),
.B2(n_137),
.Y(n_918)
);

AOI211xp5_ASAP7_75t_SL g919 ( 
.A1(n_912),
.A2(n_134),
.B(n_136),
.C(n_138),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_910),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_915),
.A2(n_266),
.B1(n_140),
.B2(n_142),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_916),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_913),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_910),
.A2(n_266),
.B1(n_144),
.B2(n_145),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_920),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_923),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_918),
.Y(n_927)
);

NAND4xp25_ASAP7_75t_L g928 ( 
.A(n_927),
.B(n_922),
.C(n_919),
.D(n_917),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_926),
.A2(n_921),
.B1(n_924),
.B2(n_266),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_925),
.A2(n_266),
.B1(n_146),
.B2(n_147),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_928),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_930),
.Y(n_932)
);

AOI211xp5_ASAP7_75t_L g933 ( 
.A1(n_931),
.A2(n_929),
.B(n_149),
.C(n_150),
.Y(n_933)
);

AOI31xp33_ASAP7_75t_L g934 ( 
.A1(n_932),
.A2(n_139),
.A3(n_151),
.B(n_154),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_933),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_934),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_936),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.C(n_161),
.Y(n_937)
);

AOI211xp5_ASAP7_75t_L g938 ( 
.A1(n_937),
.A2(n_935),
.B(n_163),
.C(n_166),
.Y(n_938)
);


endmodule