module fake_jpeg_5415_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_12),
.B1(n_20),
.B2(n_16),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_37),
.B1(n_18),
.B2(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_12),
.B1(n_19),
.B2(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_18),
.B1(n_10),
.B2(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_21),
.A2(n_20),
.B1(n_19),
.B2(n_12),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_43),
.B1(n_30),
.B2(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_35),
.B1(n_32),
.B2(n_37),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_26),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_29),
.B(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_29),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.C(n_57),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_28),
.C(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_46),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_30),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_27),
.B(n_26),
.Y(n_75)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_55),
.B1(n_51),
.B2(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_15),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_65),
.C(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_72),
.C(n_75),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_77),
.B1(n_14),
.B2(n_17),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_47),
.C(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_75),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_17),
.B(n_26),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_85),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_61),
.B1(n_17),
.B2(n_14),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_89)
);

OAI322xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_27),
.A3(n_26),
.B1(n_14),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_83)
);

OA21x2_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_9),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

OA21x2_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_27),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_2),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_82),
.B(n_9),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_78),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_95),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_96),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_79),
.C(n_85),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_93),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_90),
.B1(n_87),
.B2(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_99),
.B(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_3),
.B(n_5),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_100),
.B1(n_5),
.B2(n_98),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_104),
.Y(n_108)
);


endmodule