module fake_ariane_1950_n_1660 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1660);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1660;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_97),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_24),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

BUFx8_ASAP7_75t_SL g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_25),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_39),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_48),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_73),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_85),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_83),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_79),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_66),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_58),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_25),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_9),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_109),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_42),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_119),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_98),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_61),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_3),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_35),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_50),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_147),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_45),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_19),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_71),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_41),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_52),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_91),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_60),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_67),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_27),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_80),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_42),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_57),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_5),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_30),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_78),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_93),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_26),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_103),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_89),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_130),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_124),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_56),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_21),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_11),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_106),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_59),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_108),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_62),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_0),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_35),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_6),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_105),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_22),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_90),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_111),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_121),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_112),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_47),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_86),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_13),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_96),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_125),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_1),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_127),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_117),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_40),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_81),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_87),
.Y(n_268)
);

BUFx8_ASAP7_75t_SL g269 ( 
.A(n_55),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_31),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_22),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_34),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_145),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_70),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_34),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_69),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_126),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_32),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_33),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_1),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_84),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_134),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_31),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_37),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_17),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_2),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_155),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_155),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_156),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_153),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_156),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_164),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_200),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_164),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_181),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_211),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_203),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_181),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_183),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_184),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_184),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_197),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_197),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_206),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_206),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_228),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_230),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_208),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_223),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_238),
.Y(n_330)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_149),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_239),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_205),
.Y(n_335)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_180),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_203),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_250),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_190),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_180),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_157),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_180),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_158),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_209),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_165),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_174),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_258),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_261),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_175),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_176),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_270),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_189),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_270),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_279),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_193),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_203),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_203),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_241),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_241),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_241),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_241),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_194),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_322),
.A2(n_248),
.B1(n_268),
.B2(n_278),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_248),
.B1(n_268),
.B2(n_278),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_194),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_361),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_370),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_241),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_304),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_309),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

CKINVDCx6p67_ASAP7_75t_R g397 ( 
.A(n_307),
.Y(n_397)
);

BUFx8_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_297),
.B(n_232),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g402 ( 
.A(n_297),
.B(n_190),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_343),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_298),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_298),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_346),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_299),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_299),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_315),
.A2(n_244),
.B1(n_277),
.B2(n_286),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_301),
.B(n_232),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_301),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_312),
.A2(n_296),
.B1(n_294),
.B2(n_186),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_303),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_303),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_306),
.B(n_204),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_324),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_349),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_331),
.B(n_247),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_308),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_308),
.B(n_204),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_311),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_311),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_313),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_313),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_314),
.B(n_207),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_342),
.B(n_224),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_314),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_316),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_198),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_317),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_355),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_347),
.B(n_207),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_318),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_330),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_318),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_418),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_380),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_402),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_421),
.B(n_360),
.Y(n_445)
);

INVx4_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_420),
.B(n_365),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_302),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_394),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_400),
.B(n_412),
.Y(n_450)
);

BUFx4f_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_400),
.B(n_319),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_395),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_418),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_418),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_SL g459 ( 
.A(n_437),
.B(n_199),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g460 ( 
.A1(n_402),
.A2(n_344),
.B1(n_335),
.B2(n_325),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_389),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_319),
.Y(n_463)
);

CKINVDCx6p67_ASAP7_75t_R g464 ( 
.A(n_397),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_412),
.B(n_320),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_320),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_412),
.B(n_323),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_412),
.B(n_402),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_393),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_374),
.B(n_323),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_326),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_408),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_393),
.B(n_326),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_407),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_431),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_393),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_378),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_419),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_393),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_440),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_375),
.A2(n_289),
.B1(n_271),
.B2(n_201),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_431),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_377),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_411),
.A2(n_273),
.B1(n_222),
.B2(n_225),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_426),
.B(n_327),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_327),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_373),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_426),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

BUFx10_ASAP7_75t_L g502 ( 
.A(n_417),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_405),
.B(n_328),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_436),
.B(n_376),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_426),
.B(n_328),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_410),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_373),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_426),
.B(n_329),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_379),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_398),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_379),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_413),
.B(n_329),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_378),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_415),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_409),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_433),
.B(n_332),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_423),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_409),
.B(n_167),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_398),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_429),
.A2(n_333),
.B(n_332),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_382),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_397),
.B(n_166),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_382),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_378),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_383),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_383),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_386),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_416),
.B(n_333),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_378),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_416),
.B(n_334),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_385),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_387),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_378),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_425),
.B(n_334),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_398),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_398),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_391),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_427),
.B(n_348),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_427),
.B(n_195),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_415),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_423),
.B(n_428),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_430),
.B(n_348),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_411),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_386),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_423),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_399),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_401),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_432),
.B(n_435),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_401),
.Y(n_559)
);

NOR2x1p5_ASAP7_75t_L g560 ( 
.A(n_423),
.B(n_151),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_381),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_432),
.Y(n_562)
);

BUFx6f_ASAP7_75t_SL g563 ( 
.A(n_428),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_435),
.B(n_350),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_381),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_422),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_422),
.B(n_350),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_381),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_381),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_381),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_424),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_381),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_403),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_424),
.B(n_351),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_403),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_403),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_434),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_428),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_428),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_403),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_434),
.B(n_351),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_439),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_414),
.B(n_438),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_439),
.B(n_352),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_438),
.B(n_352),
.Y(n_586)
);

INVx8_ASAP7_75t_L g587 ( 
.A(n_403),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_414),
.A2(n_284),
.B1(n_249),
.B2(n_245),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_518),
.B(n_353),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_444),
.A2(n_359),
.B1(n_364),
.B2(n_363),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_444),
.B(n_463),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_463),
.B(n_257),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_L g594 ( 
.A1(n_469),
.A2(n_359),
.B1(n_364),
.B2(n_363),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_531),
.B(n_353),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_484),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_506),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_463),
.B(n_357),
.Y(n_598)
);

AO22x2_ASAP7_75t_L g599 ( 
.A1(n_470),
.A2(n_358),
.B1(n_362),
.B2(n_357),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_499),
.B(n_358),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_542),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_472),
.B(n_362),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_473),
.B(n_151),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_542),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_392),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_443),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_584),
.A2(n_253),
.B1(n_259),
.B2(n_242),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_499),
.B(n_224),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_551),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_473),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_491),
.B(n_169),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_468),
.B(n_255),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_499),
.B(n_287),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_475),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_551),
.B(n_253),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_562),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_441),
.B(n_259),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_481),
.B(n_287),
.Y(n_619)
);

A2O1A1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_450),
.A2(n_296),
.B(n_294),
.C(n_186),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_469),
.B(n_154),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_558),
.A2(n_154),
.B(n_215),
.C(n_219),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_453),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_481),
.B(n_150),
.Y(n_624)
);

A2O1A1Ixp33_ASAP7_75t_L g625 ( 
.A1(n_532),
.A2(n_242),
.B(n_215),
.C(n_219),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_526),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_L g627 ( 
.A(n_445),
.B(n_454),
.C(n_449),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_469),
.A2(n_172),
.B1(n_162),
.B2(n_161),
.Y(n_628)
);

NOR3xp33_ASAP7_75t_L g629 ( 
.A(n_449),
.B(n_221),
.C(n_233),
.Y(n_629)
);

INVx8_ASAP7_75t_L g630 ( 
.A(n_469),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_465),
.A2(n_178),
.B(n_160),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_586),
.B(n_221),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_586),
.Y(n_633)
);

NOR3xp33_ASAP7_75t_L g634 ( 
.A(n_454),
.B(n_488),
.C(n_485),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_233),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_503),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_464),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_481),
.B(n_150),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_513),
.B(n_226),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_513),
.B(n_234),
.Y(n_640)
);

INVxp33_ASAP7_75t_L g641 ( 
.A(n_552),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_243),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_555),
.B(n_243),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_485),
.B(n_272),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_465),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_513),
.B(n_246),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_452),
.B(n_263),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_555),
.B(n_272),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_563),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_567),
.A2(n_281),
.B(n_291),
.C(n_290),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_560),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_466),
.B(n_266),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_474),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_456),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_464),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_578),
.B(n_579),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_504),
.B(n_280),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_490),
.B(n_160),
.Y(n_659)
);

OAI221xp5_ASAP7_75t_L g660 ( 
.A1(n_489),
.A2(n_578),
.B1(n_579),
.B2(n_584),
.C(n_588),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_456),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_494),
.B(n_285),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_494),
.B(n_293),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_488),
.B(n_511),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_493),
.A2(n_212),
.B(n_178),
.C(n_196),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_484),
.A2(n_264),
.B1(n_260),
.B2(n_212),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_479),
.A2(n_152),
.B1(n_282),
.B2(n_276),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_461),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_480),
.B(n_148),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_584),
.B(n_231),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_490),
.B(n_196),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_460),
.B(n_167),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_517),
.A2(n_264),
.B(n_260),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_471),
.B(n_159),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_498),
.B(n_163),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_462),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_523),
.B(n_168),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_563),
.B(n_0),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_451),
.A2(n_210),
.B(n_218),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_170),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_459),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_471),
.B(n_171),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_462),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_482),
.B(n_210),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_547),
.B(n_173),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_524),
.B(n_177),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_482),
.B(n_486),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_502),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_584),
.B(n_2),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_524),
.B(n_179),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_502),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_511),
.Y(n_693)
);

BUFx6f_ASAP7_75t_SL g694 ( 
.A(n_475),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_500),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_527),
.Y(n_696)
);

OAI221xp5_ASAP7_75t_L g697 ( 
.A1(n_549),
.A2(n_167),
.B1(n_283),
.B2(n_231),
.C(n_265),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_486),
.A2(n_288),
.B1(n_182),
.B2(n_274),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_524),
.B(n_229),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_505),
.B(n_227),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_514),
.B(n_236),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_535),
.B(n_220),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_502),
.A2(n_185),
.B1(n_262),
.B2(n_254),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_492),
.A2(n_283),
.B1(n_195),
.B2(n_235),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_455),
.B(n_187),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_447),
.B(n_188),
.C(n_252),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_539),
.B(n_237),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_529),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_550),
.B(n_214),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_467),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_549),
.B(n_240),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_500),
.B(n_202),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_530),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_530),
.Y(n_715)
);

AND2x4_ASAP7_75t_SL g716 ( 
.A(n_519),
.B(n_195),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_476),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_500),
.B(n_251),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_451),
.B(n_195),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_509),
.B(n_446),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_446),
.B(n_3),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_476),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_446),
.B(n_4),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_521),
.B(n_191),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_451),
.A2(n_192),
.B(n_235),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_448),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_477),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_501),
.B(n_283),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_501),
.B(n_4),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_564),
.B(n_540),
.C(n_521),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_501),
.B(n_235),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_507),
.B(n_7),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_507),
.B(n_8),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_507),
.B(n_522),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_522),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_536),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_477),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_522),
.B(n_235),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_566),
.B(n_9),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_455),
.B(n_235),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_455),
.B(n_10),
.Y(n_743)
);

OAI21xp33_ASAP7_75t_L g744 ( 
.A1(n_537),
.A2(n_195),
.B(n_11),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_554),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_487),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_566),
.B(n_10),
.Y(n_747)
);

BUFx6f_ASAP7_75t_SL g748 ( 
.A(n_637),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_705),
.A2(n_571),
.B1(n_577),
.B2(n_582),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_615),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_611),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_745),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_602),
.B(n_540),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_740),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_617),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_695),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_637),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_660),
.A2(n_541),
.B1(n_571),
.B2(n_582),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_677),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_656),
.B(n_633),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_630),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_594),
.B(n_483),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_594),
.B(n_483),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_656),
.B(n_653),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_746),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_693),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_689),
.B(n_517),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

BUFx8_ASAP7_75t_SL g771 ( 
.A(n_694),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_595),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_644),
.B(n_574),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_693),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_746),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_589),
.B(n_543),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_592),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_641),
.B(n_543),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_591),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_630),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_702),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_709),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_734),
.A2(n_553),
.B(n_548),
.Y(n_783)
);

NOR2x1_ASAP7_75t_R g784 ( 
.A(n_651),
.B(n_581),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_649),
.B(n_585),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_692),
.B(n_603),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_726),
.B(n_548),
.Y(n_787)
);

NOR2x2_ASAP7_75t_L g788 ( 
.A(n_670),
.B(n_495),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_604),
.B(n_496),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_607),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_654),
.Y(n_791)
);

OAI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_670),
.A2(n_553),
.B1(n_556),
.B2(n_508),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_714),
.B(n_715),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_636),
.B(n_556),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_731),
.B(n_496),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_694),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_737),
.B(n_544),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_670),
.B(n_621),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_654),
.B(n_544),
.Y(n_799)
);

INVx3_ASAP7_75t_SL g800 ( 
.A(n_693),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_719),
.A2(n_442),
.B(n_458),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_590),
.B(n_510),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_590),
.B(n_510),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_645),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_649),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_735),
.A2(n_442),
.B(n_457),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_616),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_658),
.A2(n_457),
.B1(n_458),
.B2(n_508),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_654),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_599),
.B(n_613),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_599),
.B(n_591),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_690),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_599),
.B(n_559),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_598),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_608),
.A2(n_559),
.B1(n_512),
.B2(n_534),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_692),
.B(n_533),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_608),
.A2(n_557),
.B1(n_512),
.B2(n_534),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_672),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_598),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_705),
.A2(n_557),
.B1(n_478),
.B2(n_520),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_634),
.B(n_478),
.Y(n_821)
);

CKINVDCx11_ASAP7_75t_R g822 ( 
.A(n_627),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_639),
.B(n_483),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_716),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_597),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_601),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_679),
.B(n_565),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_596),
.Y(n_828)
);

OAI21xp33_ASAP7_75t_L g829 ( 
.A1(n_639),
.A2(n_576),
.B(n_533),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_736),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_623),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_626),
.B(n_576),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_716),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_606),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_605),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_736),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_610),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_655),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_632),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_679),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_682),
.B(n_576),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_730),
.B(n_573),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_635),
.Y(n_844)
);

O2A1O1Ixp5_ASAP7_75t_L g845 ( 
.A1(n_734),
.A2(n_533),
.B(n_538),
.C(n_573),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_593),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_668),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_676),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_684),
.Y(n_849)
);

BUFx4f_ASAP7_75t_L g850 ( 
.A(n_711),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_717),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_722),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_629),
.B(n_520),
.Y(n_853)
);

BUFx8_ASAP7_75t_SL g854 ( 
.A(n_662),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_612),
.B(n_538),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_657),
.B(n_538),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_727),
.B(n_573),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_738),
.B(n_565),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_643),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_663),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_618),
.B(n_600),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_741),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_721),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_640),
.B(n_483),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_648),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_600),
.A2(n_587),
.B(n_583),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_640),
.B(n_568),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_646),
.B(n_568),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_593),
.B(n_570),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_747),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_647),
.A2(n_520),
.B1(n_583),
.B2(n_580),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_729),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_642),
.B(n_561),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_646),
.B(n_720),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_647),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_720),
.B(n_561),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_724),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_728),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_733),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_687),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_628),
.B(n_497),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_673),
.B(n_569),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_620),
.B(n_569),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_652),
.A2(n_520),
.B1(n_580),
.B2(n_575),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_707),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_659),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_688),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_659),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_671),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_652),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_620),
.B(n_575),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_691),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_683),
.A2(n_520),
.B1(n_587),
.B2(n_570),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_701),
.B(n_572),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_704),
.B(n_497),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_671),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_703),
.B(n_572),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_712),
.B(n_520),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_674),
.Y(n_899)
);

NAND2x1_ASAP7_75t_L g900 ( 
.A(n_743),
.B(n_497),
.Y(n_900)
);

HB1xp67_ASAP7_75t_SL g901 ( 
.A(n_697),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_624),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_624),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_SL g904 ( 
.A(n_650),
.B(n_12),
.C(n_13),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_638),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_688),
.B(n_515),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_638),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_743),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_631),
.Y(n_909)
);

NAND2x1_ASAP7_75t_L g910 ( 
.A(n_721),
.B(n_497),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_685),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_669),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_R g913 ( 
.A(n_723),
.B(n_546),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_685),
.A2(n_520),
.B1(n_587),
.B2(n_546),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_732),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_622),
.A2(n_528),
.B1(n_515),
.B2(n_587),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_622),
.B(n_528),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_723),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_708),
.B(n_528),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_675),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_875),
.A2(n_650),
.B(n_625),
.C(n_678),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_874),
.A2(n_706),
.B(n_614),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_756),
.Y(n_923)
);

O2A1O1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_875),
.A2(n_625),
.B(n_710),
.C(n_609),
.Y(n_924)
);

INVx3_ASAP7_75t_SL g925 ( 
.A(n_796),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_772),
.B(n_698),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_794),
.B(n_700),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_863),
.A2(n_874),
.B(n_787),
.C(n_912),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_752),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_863),
.A2(n_609),
.B(n_614),
.C(n_619),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_776),
.A2(n_719),
.B(n_718),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_760),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_890),
.B(n_667),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_751),
.Y(n_934)
);

BUFx12f_ASAP7_75t_L g935 ( 
.A(n_809),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_908),
.A2(n_699),
.B(n_739),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_841),
.B(n_681),
.Y(n_937)
);

O2A1O1Ixp5_ASAP7_75t_SL g938 ( 
.A1(n_823),
.A2(n_619),
.B(n_742),
.C(n_739),
.Y(n_938)
);

O2A1O1Ixp5_ASAP7_75t_L g939 ( 
.A1(n_910),
.A2(n_713),
.B(n_732),
.C(n_742),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_776),
.A2(n_744),
.B1(n_666),
.B2(n_686),
.Y(n_940)
);

AOI22x1_ASAP7_75t_L g941 ( 
.A1(n_783),
.A2(n_725),
.B1(n_680),
.B2(n_665),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_778),
.B(n_528),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_768),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_900),
.A2(n_515),
.B(n_54),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_762),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_920),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_783),
.A2(n_515),
.B(n_72),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_762),
.B(n_20),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_793),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_757),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_SL g951 ( 
.A1(n_750),
.A2(n_800),
.B1(n_754),
.B2(n_755),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_867),
.A2(n_868),
.B(n_919),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_777),
.Y(n_953)
);

AOI221xp5_ASAP7_75t_L g954 ( 
.A1(n_904),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_954)
);

BUFx8_ASAP7_75t_L g955 ( 
.A(n_748),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_771),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_790),
.Y(n_957)
);

OR2x6_ASAP7_75t_SL g958 ( 
.A(n_798),
.B(n_38),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_773),
.B(n_40),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_R g960 ( 
.A(n_767),
.B(n_95),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_904),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_786),
.A2(n_43),
.B(n_46),
.C(n_63),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_867),
.A2(n_64),
.B(n_75),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_834),
.B(n_100),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_822),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_901),
.B(n_115),
.Y(n_966)
);

INVx5_ASAP7_75t_L g967 ( 
.A(n_762),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_901),
.A2(n_120),
.B1(n_133),
.B2(n_140),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_806),
.A2(n_143),
.B(n_801),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_864),
.A2(n_868),
.B(n_882),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_758),
.B(n_799),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_774),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_793),
.A2(n_797),
.B1(n_795),
.B2(n_918),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_805),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_870),
.A2(n_860),
.B(n_879),
.C(n_862),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_919),
.A2(n_897),
.B(n_894),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_806),
.A2(n_866),
.B(n_845),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_753),
.Y(n_978)
);

CKINVDCx14_ASAP7_75t_R g979 ( 
.A(n_791),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_791),
.B(n_748),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_799),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_831),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_846),
.A2(n_804),
.B(n_865),
.C(n_859),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_834),
.B(n_807),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_894),
.A2(n_897),
.B(n_829),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_795),
.A2(n_797),
.B(n_866),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_918),
.A2(n_781),
.B1(n_782),
.B2(n_817),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_839),
.B(n_844),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_765),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_789),
.B(n_846),
.Y(n_990)
);

AND2x2_ASAP7_75t_SL g991 ( 
.A(n_810),
.B(n_811),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_847),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_838),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_876),
.A2(n_856),
.B(n_861),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_765),
.B(n_825),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_779),
.B(n_814),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_821),
.A2(n_861),
.B(n_810),
.C(n_792),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_779),
.B(n_819),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_759),
.A2(n_855),
.B(n_869),
.C(n_808),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_876),
.A2(n_856),
.B(n_845),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_854),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_872),
.A2(n_763),
.B(n_764),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_770),
.B(n_791),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_885),
.A2(n_837),
.B(n_826),
.C(n_835),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_770),
.B(n_791),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_780),
.B(n_850),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_761),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_818),
.A2(n_812),
.B1(n_892),
.B2(n_880),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_815),
.A2(n_880),
.B(n_892),
.C(n_898),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_780),
.B(n_832),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_877),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_802),
.B(n_803),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_799),
.B(n_785),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_802),
.B(n_803),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_877),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_832),
.B(n_836),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_828),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_852),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_916),
.A2(n_766),
.B(n_775),
.C(n_842),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_917),
.A2(n_749),
.B1(n_820),
.B2(n_813),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_883),
.A2(n_891),
.B(n_813),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_850),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_785),
.B(n_843),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_878),
.B(n_827),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_827),
.B(n_811),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_916),
.A2(n_917),
.B(n_881),
.C(n_873),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_828),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_882),
.A2(n_909),
.B(n_883),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_827),
.A2(n_853),
.B1(n_843),
.B2(n_917),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_891),
.A2(n_857),
.B(n_907),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_827),
.B(n_848),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_824),
.B(n_833),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_858),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_824),
.B(n_833),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_886),
.Y(n_1036)
);

INVx3_ASAP7_75t_SL g1037 ( 
.A(n_788),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_895),
.A2(n_911),
.B(n_903),
.C(n_902),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_899),
.B(n_784),
.C(n_888),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_896),
.A2(n_905),
.B(n_889),
.C(n_914),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_871),
.B(n_884),
.C(n_830),
.Y(n_1041)
);

CKINVDCx6p67_ASAP7_75t_R g1042 ( 
.A(n_840),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_828),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_816),
.A2(n_893),
.B(n_915),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_887),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_816),
.A2(n_769),
.B(n_906),
.Y(n_1046)
);

AO32x2_ASAP7_75t_L g1047 ( 
.A1(n_913),
.A2(n_887),
.A3(n_840),
.B1(n_851),
.B2(n_769),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_906),
.A2(n_875),
.B(n_874),
.C(n_445),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_928),
.A2(n_840),
.B(n_927),
.Y(n_1049)
);

INVxp67_ASAP7_75t_SL g1050 ( 
.A(n_973),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_976),
.A2(n_994),
.B(n_1000),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_984),
.B(n_937),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_921),
.A2(n_1048),
.B(n_999),
.C(n_924),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_974),
.B(n_990),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_923),
.Y(n_1055)
);

AOI21xp33_ASAP7_75t_SL g1056 ( 
.A1(n_925),
.A2(n_951),
.B(n_949),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_986),
.A2(n_973),
.B(n_985),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_980),
.Y(n_1058)
);

AO32x2_ASAP7_75t_L g1059 ( 
.A1(n_987),
.A2(n_1021),
.A3(n_949),
.B1(n_940),
.B2(n_991),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_984),
.B(n_974),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_970),
.A2(n_936),
.B(n_987),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_932),
.Y(n_1062)
);

AO21x2_ASAP7_75t_L g1063 ( 
.A1(n_1022),
.A2(n_1026),
.B(n_1014),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_SL g1064 ( 
.A(n_956),
.B(n_1001),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_943),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_929),
.B(n_1010),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_969),
.A2(n_977),
.B(n_1029),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_933),
.B(n_1024),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_922),
.A2(n_930),
.B(n_931),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1044),
.A2(n_944),
.B(n_947),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_989),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_959),
.B(n_996),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_967),
.B(n_945),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_998),
.B(n_975),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1024),
.B(n_1013),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_1013),
.B(n_926),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_988),
.B(n_1035),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_954),
.A2(n_940),
.B(n_966),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1027),
.A2(n_1020),
.B(n_1002),
.Y(n_1079)
);

NAND3x1_ASAP7_75t_L g1080 ( 
.A(n_958),
.B(n_968),
.C(n_955),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1012),
.A2(n_963),
.B(n_1031),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_978),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_983),
.B(n_1033),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1033),
.B(n_1007),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_995),
.B(n_1016),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1031),
.A2(n_1046),
.B(n_1009),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_934),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_993),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_981),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_939),
.B(n_1004),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_1022),
.A2(n_1026),
.B(n_1025),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1037),
.B(n_1039),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_955),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1021),
.A2(n_1030),
.B1(n_1011),
.B2(n_981),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1019),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_967),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_967),
.B(n_945),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1023),
.B(n_1008),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_938),
.A2(n_941),
.B(n_1038),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_948),
.B(n_1041),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1006),
.B(n_1045),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1040),
.A2(n_1032),
.B(n_964),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_997),
.A2(n_1036),
.B(n_1034),
.Y(n_1103)
);

BUFx4f_ASAP7_75t_L g1104 ( 
.A(n_935),
.Y(n_1104)
);

AO21x1_ASAP7_75t_L g1105 ( 
.A1(n_961),
.A2(n_962),
.B(n_946),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_953),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_972),
.B(n_992),
.Y(n_1107)
);

AO21x2_ASAP7_75t_L g1108 ( 
.A1(n_950),
.A2(n_957),
.B(n_1018),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_982),
.A2(n_1047),
.A3(n_1042),
.B(n_1043),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1047),
.A2(n_979),
.B(n_1043),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1017),
.A2(n_971),
.A3(n_1028),
.B(n_960),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1017),
.A2(n_971),
.A3(n_1003),
.B(n_1005),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1015),
.B(n_965),
.Y(n_1113)
);

AO21x1_ASAP7_75t_L g1114 ( 
.A1(n_973),
.A2(n_863),
.B(n_874),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_927),
.A2(n_863),
.B1(n_874),
.B2(n_875),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_928),
.A2(n_875),
.B(n_445),
.C(n_421),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_923),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_SL g1121 ( 
.A1(n_927),
.A2(n_874),
.B(n_642),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_936),
.A2(n_976),
.A3(n_952),
.B(n_985),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_959),
.B(n_644),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_923),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_923),
.Y(n_1126)
);

NOR4xp25_ASAP7_75t_L g1127 ( 
.A(n_949),
.B(n_904),
.C(n_921),
.D(n_946),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_921),
.A2(n_421),
.B1(n_588),
.B2(n_375),
.C(n_322),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_952),
.A2(n_874),
.B(n_863),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_923),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_952),
.A2(n_874),
.B(n_863),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_SL g1132 ( 
.A1(n_927),
.A2(n_874),
.B(n_642),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_927),
.A2(n_863),
.B1(n_874),
.B2(n_875),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_967),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_984),
.B(n_449),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_952),
.A2(n_874),
.B(n_863),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_923),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_984),
.B(n_449),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_SL g1144 ( 
.A(n_956),
.B(n_449),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1145)
);

OAI22x1_ASAP7_75t_L g1146 ( 
.A1(n_966),
.A2(n_411),
.B1(n_841),
.B2(n_875),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_974),
.B(n_449),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_959),
.B(n_644),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_921),
.A2(n_875),
.B(n_863),
.C(n_1048),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_921),
.A2(n_875),
.B(n_863),
.C(n_1048),
.Y(n_1151)
);

AND2x6_ASAP7_75t_L g1152 ( 
.A(n_1030),
.B(n_948),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_984),
.B(n_449),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1013),
.B(n_762),
.Y(n_1154)
);

BUFx4f_ASAP7_75t_L g1155 ( 
.A(n_925),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_981),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_936),
.A2(n_976),
.A3(n_952),
.B(n_985),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_927),
.A2(n_863),
.B1(n_874),
.B2(n_875),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_928),
.B(n_874),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_SL g1163 ( 
.A1(n_954),
.A2(n_421),
.B(n_875),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1164)
);

AND2x2_ASAP7_75t_SL g1165 ( 
.A(n_981),
.B(n_966),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_967),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_630),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_981),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_923),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_921),
.A2(n_875),
.B(n_863),
.C(n_1048),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_934),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_969),
.A2(n_977),
.B(n_986),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_928),
.A2(n_874),
.B(n_863),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1013),
.B(n_762),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_973),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_981),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1070),
.A2(n_1067),
.B(n_1117),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1118),
.A2(n_1124),
.B(n_1119),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1083),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1060),
.Y(n_1181)
);

AOI221xp5_ASAP7_75t_L g1182 ( 
.A1(n_1128),
.A2(n_1078),
.B1(n_1127),
.B2(n_1163),
.C(n_1146),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_SL g1183 ( 
.A(n_1166),
.B(n_1094),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1134),
.A2(n_1139),
.B(n_1136),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1155),
.Y(n_1185)
);

BUFx10_ASAP7_75t_L g1186 ( 
.A(n_1093),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_1155),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1074),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1166),
.B(n_1154),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_SL g1191 ( 
.A1(n_1100),
.A2(n_1152),
.B1(n_1165),
.B2(n_1050),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1145),
.A2(n_1158),
.B(n_1147),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1168),
.A2(n_1173),
.B(n_1099),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1112),
.B(n_1152),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1078),
.A2(n_1163),
.B(n_1116),
.C(n_1053),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1052),
.B(n_1137),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1104),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1069),
.A2(n_1051),
.B(n_1057),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1141),
.B(n_1153),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1112),
.B(n_1152),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1123),
.A2(n_1149),
.B1(n_1115),
.B2(n_1160),
.Y(n_1201)
);

OAI221xp5_ASAP7_75t_L g1202 ( 
.A1(n_1127),
.A2(n_1148),
.B1(n_1056),
.B2(n_1151),
.C(n_1171),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1133),
.B(n_1077),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1061),
.A2(n_1102),
.B(n_1081),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1076),
.B(n_1054),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1154),
.B(n_1175),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1089),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1062),
.Y(n_1208)
);

INVx4_ASAP7_75t_SL g1209 ( 
.A(n_1152),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1066),
.B(n_1072),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1176),
.A2(n_1164),
.B(n_1156),
.C(n_1161),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1150),
.A2(n_1162),
.B(n_1143),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1079),
.A2(n_1129),
.B(n_1138),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_1167),
.B(n_1110),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1090),
.A2(n_1086),
.B(n_1131),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1103),
.A2(n_1132),
.B(n_1121),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1065),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1100),
.A2(n_1143),
.B1(n_1174),
.B2(n_1161),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1049),
.A2(n_1156),
.B(n_1174),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1120),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_1092),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1125),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1056),
.A2(n_1080),
.B1(n_1085),
.B2(n_1068),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1105),
.A2(n_1095),
.B1(n_1088),
.B2(n_1098),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1126),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1167),
.B(n_1175),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1075),
.B(n_1071),
.Y(n_1227)
);

OR2x6_ASAP7_75t_L g1228 ( 
.A(n_1089),
.B(n_1177),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1089),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1130),
.A2(n_1140),
.B1(n_1170),
.B2(n_1059),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1106),
.A2(n_1091),
.B1(n_1172),
.B2(n_1087),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1108),
.A2(n_1084),
.B(n_1107),
.Y(n_1232)
);

NAND3xp33_ASAP7_75t_L g1233 ( 
.A(n_1144),
.B(n_1101),
.C(n_1096),
.Y(n_1233)
);

INVx6_ASAP7_75t_L g1234 ( 
.A(n_1157),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1113),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1111),
.B(n_1109),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1157),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1135),
.A2(n_1073),
.B(n_1097),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1064),
.A2(n_1122),
.B(n_1159),
.C(n_1111),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1122),
.A2(n_1159),
.B(n_1109),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1169),
.A2(n_1163),
.B1(n_863),
.B2(n_875),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1169),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1055),
.Y(n_1243)
);

AO21x2_ASAP7_75t_L g1244 ( 
.A1(n_1102),
.A2(n_952),
.B(n_1090),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1058),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_SL g1246 ( 
.A1(n_1142),
.A2(n_1156),
.B(n_1143),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1052),
.B(n_1060),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1052),
.B(n_1060),
.Y(n_1248)
);

INVx5_ASAP7_75t_SL g1249 ( 
.A(n_1089),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1055),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1082),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1091),
.Y(n_1252)
);

OAI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1068),
.A2(n_411),
.B1(n_454),
.B2(n_449),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1083),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1150),
.A2(n_874),
.B(n_1171),
.C(n_1151),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1082),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1078),
.A2(n_414),
.B1(n_1146),
.B2(n_402),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1082),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1089),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1063),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1055),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1070),
.A2(n_1067),
.B(n_1173),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1063),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1055),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1163),
.A2(n_863),
.B1(n_875),
.B2(n_1137),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1082),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_952),
.B(n_1090),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1055),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1055),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1078),
.A2(n_863),
.B(n_874),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1093),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1063),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1051),
.A2(n_1057),
.B(n_1069),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1078),
.A2(n_863),
.B(n_874),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1078),
.A2(n_554),
.B1(n_664),
.B2(n_1128),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1055),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1070),
.A2(n_1067),
.B(n_1173),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1114),
.A2(n_936),
.A3(n_952),
.B(n_1102),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1070),
.A2(n_1067),
.B(n_1173),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1055),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1055),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1078),
.A2(n_863),
.B(n_874),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1070),
.A2(n_1067),
.B(n_1173),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1055),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1195),
.A2(n_1202),
.B(n_1182),
.C(n_1265),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1189),
.B(n_1180),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1195),
.A2(n_1189),
.B(n_1183),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1187),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1180),
.B(n_1254),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1254),
.B(n_1203),
.Y(n_1290)
);

CKINVDCx6p67_ASAP7_75t_R g1291 ( 
.A(n_1197),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1209),
.B(n_1194),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1239),
.A2(n_1274),
.B(n_1270),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1241),
.A2(n_1255),
.B(n_1223),
.C(n_1212),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1255),
.A2(n_1282),
.B(n_1211),
.C(n_1257),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1208),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1275),
.A2(n_1257),
.B1(n_1218),
.B2(n_1201),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1210),
.B(n_1205),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1258),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1271),
.Y(n_1300)
);

NOR3xp33_ASAP7_75t_L g1301 ( 
.A(n_1233),
.B(n_1199),
.C(n_1196),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1211),
.A2(n_1273),
.B(n_1218),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1217),
.Y(n_1303)
);

A2O1A1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1191),
.A2(n_1224),
.B(n_1219),
.C(n_1201),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1191),
.A2(n_1224),
.B1(n_1251),
.B2(n_1221),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1220),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1222),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1271),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_1252),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1247),
.B(n_1248),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1225),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1227),
.B(n_1266),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1181),
.B(n_1230),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1181),
.B(n_1284),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1250),
.B(n_1261),
.Y(n_1316)
);

AOI221x1_ASAP7_75t_SL g1317 ( 
.A1(n_1264),
.A2(n_1281),
.B1(n_1280),
.B2(n_1269),
.C(n_1268),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1215),
.A2(n_1276),
.B1(n_1188),
.B2(n_1197),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1204),
.A2(n_1193),
.B(n_1198),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1209),
.B(n_1226),
.Y(n_1320)
);

AND2x6_ASAP7_75t_L g1321 ( 
.A(n_1194),
.B(n_1200),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1232),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1273),
.A2(n_1267),
.B(n_1244),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1200),
.B(n_1214),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1226),
.B(n_1256),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1188),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1246),
.B(n_1215),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1235),
.A2(n_1256),
.B(n_1186),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1215),
.A2(n_1200),
.B1(n_1245),
.B2(n_1185),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1245),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1240),
.A2(n_1237),
.B(n_1242),
.C(n_1213),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1235),
.A2(n_1206),
.B1(n_1226),
.B2(n_1190),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1229),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1240),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1229),
.B(n_1259),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1178),
.A2(n_1283),
.B(n_1279),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1190),
.A2(n_1234),
.B1(n_1207),
.B2(n_1249),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1259),
.A2(n_1253),
.B(n_1228),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_1186),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1259),
.B(n_1249),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1242),
.A2(n_1236),
.B(n_1216),
.C(n_1231),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1207),
.A2(n_1234),
.B1(n_1231),
.B2(n_1263),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1260),
.A2(n_1272),
.B(n_1263),
.C(n_1278),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1234),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1278),
.A2(n_1238),
.B(n_1277),
.C(n_1262),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1278),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1179),
.A2(n_1078),
.B(n_1182),
.C(n_1275),
.Y(n_1347)
);

AND2x2_ASAP7_75t_SL g1348 ( 
.A(n_1184),
.B(n_1192),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1205),
.B(n_1227),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1189),
.B(n_1180),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1195),
.A2(n_1078),
.B(n_863),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1255),
.A2(n_863),
.B(n_1162),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1205),
.B(n_1227),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1189),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1189),
.Y(n_1355)
);

O2A1O1Ixp5_ASAP7_75t_L g1356 ( 
.A1(n_1195),
.A2(n_1212),
.B(n_1162),
.C(n_1105),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1205),
.B(n_1227),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1205),
.B(n_1227),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1204),
.A2(n_1193),
.B(n_1198),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1255),
.A2(n_863),
.B(n_1162),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1195),
.A2(n_1212),
.B(n_1162),
.C(n_1105),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1195),
.A2(n_1163),
.B(n_1202),
.C(n_1078),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1210),
.B(n_1205),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1199),
.A2(n_1141),
.B(n_1137),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1327),
.B(n_1302),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1327),
.B(n_1323),
.Y(n_1366)
);

OAI221xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1362),
.A2(n_1285),
.B1(n_1351),
.B2(n_1295),
.C(n_1294),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1321),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1336),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1334),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1290),
.B(n_1286),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1348),
.Y(n_1372)
);

BUFx2_ASAP7_75t_SL g1373 ( 
.A(n_1329),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1356),
.A2(n_1361),
.B(n_1347),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1346),
.B(n_1319),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1290),
.B(n_1314),
.Y(n_1376)
);

OR2x6_ASAP7_75t_L g1377 ( 
.A(n_1324),
.B(n_1292),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1321),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1304),
.A2(n_1293),
.B(n_1341),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1359),
.B(n_1329),
.Y(n_1380)
);

OR2x2_ASAP7_75t_SL g1381 ( 
.A(n_1354),
.B(n_1355),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1318),
.A2(n_1331),
.B(n_1322),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1318),
.A2(n_1343),
.B(n_1297),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1286),
.B(n_1350),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1297),
.A2(n_1342),
.B(n_1350),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1309),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1342),
.A2(n_1289),
.B(n_1305),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1317),
.B(n_1315),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1288),
.B(n_1296),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1332),
.A2(n_1337),
.B(n_1360),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1303),
.B(n_1306),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1307),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1311),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1312),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1316),
.B(n_1358),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1310),
.B(n_1287),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1301),
.A2(n_1352),
.B1(n_1333),
.B2(n_1363),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1345),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1299),
.B(n_1298),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1349),
.B(n_1357),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1365),
.B(n_1353),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1402)
);

INVxp67_ASAP7_75t_SL g1403 ( 
.A(n_1386),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1386),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1376),
.B(n_1313),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1370),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1369),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1381),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1409)
);

NAND4xp25_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1364),
.C(n_1330),
.D(n_1325),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1366),
.B(n_1380),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1376),
.B(n_1335),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1376),
.B(n_1344),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1374),
.A2(n_1338),
.B(n_1340),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1380),
.B(n_1333),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1380),
.B(n_1333),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1392),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1380),
.B(n_1320),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1395),
.B(n_1375),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1395),
.B(n_1375),
.Y(n_1420)
);

NOR2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1368),
.B(n_1291),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1375),
.B(n_1326),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1368),
.Y(n_1423)
);

OR2x6_ASAP7_75t_L g1424 ( 
.A(n_1415),
.B(n_1368),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1412),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1411),
.B(n_1400),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1410),
.B(n_1339),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_SL g1428 ( 
.A(n_1423),
.B(n_1377),
.Y(n_1428)
);

OAI322xp33_ASAP7_75t_L g1429 ( 
.A1(n_1411),
.A2(n_1388),
.A3(n_1376),
.B1(n_1371),
.B2(n_1384),
.C1(n_1399),
.C2(n_1398),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1404),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1408),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1404),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1408),
.A2(n_1379),
.B1(n_1383),
.B2(n_1373),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1415),
.A2(n_1379),
.B1(n_1383),
.B2(n_1387),
.Y(n_1434)
);

AOI222xp33_ASAP7_75t_L g1435 ( 
.A1(n_1411),
.A2(n_1374),
.B1(n_1388),
.B2(n_1396),
.C1(n_1371),
.C2(n_1398),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1415),
.B(n_1378),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1408),
.A2(n_1374),
.B1(n_1367),
.B2(n_1388),
.C(n_1396),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1406),
.Y(n_1438)
);

OAI211xp5_ASAP7_75t_L g1439 ( 
.A1(n_1410),
.A2(n_1398),
.B(n_1397),
.C(n_1384),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1411),
.B(n_1402),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1414),
.A2(n_1396),
.B1(n_1373),
.B2(n_1384),
.C(n_1397),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1402),
.A2(n_1383),
.B1(n_1379),
.B2(n_1385),
.C(n_1387),
.Y(n_1442)
);

AOI21xp33_ASAP7_75t_L g1443 ( 
.A1(n_1416),
.A2(n_1379),
.B(n_1383),
.Y(n_1443)
);

AOI33xp33_ASAP7_75t_L g1444 ( 
.A1(n_1402),
.A2(n_1400),
.A3(n_1391),
.B1(n_1389),
.B2(n_1393),
.B3(n_1394),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1402),
.B(n_1399),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1400),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1413),
.A2(n_1381),
.B1(n_1373),
.B2(n_1372),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1409),
.B(n_1399),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1417),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1416),
.A2(n_1379),
.B1(n_1383),
.B2(n_1387),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1417),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_R g1452 ( 
.A(n_1416),
.B(n_1300),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1409),
.B(n_1399),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1423),
.B(n_1378),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1407),
.A2(n_1383),
.B(n_1379),
.Y(n_1455)
);

AOI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1409),
.A2(n_1390),
.B(n_1372),
.C(n_1381),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1417),
.Y(n_1457)
);

AOI211xp5_ASAP7_75t_L g1458 ( 
.A1(n_1414),
.A2(n_1372),
.B(n_1418),
.C(n_1422),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1401),
.B(n_1403),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1419),
.B(n_1385),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1449),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1424),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1431),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1455),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1455),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1455),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1419),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1438),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1427),
.B(n_1401),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1449),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1440),
.B(n_1419),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1431),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_SL g1473 ( 
.A(n_1435),
.B(n_1413),
.C(n_1422),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1444),
.B(n_1403),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1443),
.A2(n_1382),
.B(n_1387),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1451),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1437),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1424),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1454),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1451),
.Y(n_1480)
);

NOR2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1460),
.B(n_1405),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1454),
.Y(n_1482)
);

NOR2x1_ASAP7_75t_L g1483 ( 
.A(n_1429),
.B(n_1421),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1457),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1430),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1432),
.Y(n_1486)
);

CKINVDCx16_ASAP7_75t_R g1487 ( 
.A(n_1452),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1424),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1459),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1441),
.Y(n_1490)
);

NOR2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1460),
.B(n_1405),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1478),
.B(n_1426),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1478),
.B(n_1426),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1461),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1461),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1475),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1474),
.B(n_1445),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1470),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1478),
.B(n_1424),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1470),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1474),
.B(n_1486),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1476),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1490),
.B(n_1439),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1472),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1485),
.B(n_1425),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1488),
.B(n_1420),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1475),
.Y(n_1507)
);

NAND2x1_ASAP7_75t_L g1508 ( 
.A(n_1488),
.B(n_1436),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1486),
.B(n_1489),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1488),
.B(n_1428),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1485),
.B(n_1442),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1462),
.B(n_1428),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1467),
.B(n_1420),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1477),
.B(n_1433),
.C(n_1450),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1463),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1475),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1475),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1480),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1480),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1471),
.B(n_1483),
.Y(n_1521)
);

NAND2x1p5_ASAP7_75t_L g1522 ( 
.A(n_1483),
.B(n_1368),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1490),
.B(n_1445),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1446),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1489),
.B(n_1448),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1464),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1515),
.A2(n_1473),
.B1(n_1434),
.B2(n_1387),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1503),
.Y(n_1530)
);

INVx1_ASAP7_75t_SL g1531 ( 
.A(n_1516),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1522),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1509),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1509),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1516),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1494),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1523),
.B(n_1473),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1515),
.A2(n_1456),
.B(n_1458),
.C(n_1491),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1494),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1524),
.B(n_1463),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1495),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1511),
.A2(n_1464),
.B1(n_1465),
.B2(n_1466),
.C(n_1447),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1523),
.B(n_1448),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1496),
.Y(n_1545)
);

NAND2x1_ASAP7_75t_SL g1546 ( 
.A(n_1521),
.B(n_1479),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1495),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_L g1548 ( 
.A(n_1511),
.B(n_1456),
.C(n_1472),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_SL g1549 ( 
.A(n_1504),
.B(n_1487),
.Y(n_1549)
);

NOR2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1508),
.B(n_1479),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1521),
.B(n_1472),
.Y(n_1551)
);

NOR2x1_ASAP7_75t_L g1552 ( 
.A(n_1504),
.B(n_1482),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1496),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1501),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1498),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1522),
.B(n_1504),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1498),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1508),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1501),
.B(n_1453),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1500),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1492),
.B(n_1493),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1563),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1565)
);

INVx1_ASAP7_75t_SL g1566 ( 
.A(n_1531),
.Y(n_1566)
);

NOR2x1_ASAP7_75t_L g1567 ( 
.A(n_1536),
.B(n_1510),
.Y(n_1567)
);

NOR2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1551),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1533),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1537),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1563),
.B(n_1492),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1548),
.B(n_1510),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1546),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1539),
.A2(n_1458),
.B1(n_1481),
.B2(n_1491),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1505),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1540),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1549),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1493),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1554),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_1538),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1555),
.B(n_1505),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1554),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1497),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1559),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1513),
.Y(n_1587)
);

AND2x2_ASAP7_75t_SL g1588 ( 
.A(n_1529),
.B(n_1510),
.Y(n_1588)
);

CKINVDCx16_ASAP7_75t_R g1589 ( 
.A(n_1566),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1564),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1581),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1587),
.Y(n_1592)
);

AOI221xp5_ASAP7_75t_L g1593 ( 
.A1(n_1574),
.A2(n_1543),
.B1(n_1539),
.B2(n_1526),
.C(n_1518),
.Y(n_1593)
);

AOI22x1_ASAP7_75t_L g1594 ( 
.A1(n_1573),
.A2(n_1560),
.B1(n_1532),
.B2(n_1547),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1572),
.A2(n_1534),
.B(n_1552),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1575),
.A2(n_1534),
.B1(n_1557),
.B2(n_1561),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1575),
.A2(n_1496),
.B1(n_1518),
.B2(n_1526),
.C(n_1517),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1583),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1569),
.A2(n_1582),
.B(n_1577),
.C(n_1578),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1584),
.B(n_1525),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1565),
.B(n_1557),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1570),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1571),
.B(n_1506),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1588),
.A2(n_1517),
.B(n_1518),
.C(n_1507),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1308),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1570),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_L g1609 ( 
.A(n_1601),
.B(n_1567),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1591),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1589),
.B(n_1573),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1586),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1600),
.B(n_1568),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1607),
.B(n_1571),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1592),
.B(n_1587),
.Y(n_1615)
);

NOR2x1_ASAP7_75t_L g1616 ( 
.A(n_1600),
.B(n_1576),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1602),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1605),
.B(n_1584),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1615),
.B(n_1607),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_L g1620 ( 
.A(n_1613),
.B(n_1593),
.C(n_1594),
.Y(n_1620)
);

NOR3x1_ASAP7_75t_L g1621 ( 
.A(n_1611),
.B(n_1599),
.C(n_1603),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1610),
.A2(n_1596),
.B1(n_1590),
.B2(n_1595),
.C(n_1585),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_L g1623 ( 
.A1(n_1616),
.A2(n_1588),
.B1(n_1598),
.B2(n_1606),
.C1(n_1597),
.C2(n_1604),
.Y(n_1623)
);

AOI211xp5_ASAP7_75t_L g1624 ( 
.A1(n_1612),
.A2(n_1585),
.B(n_1608),
.C(n_1565),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1614),
.A2(n_1565),
.B(n_1579),
.C(n_1576),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1618),
.B(n_1579),
.Y(n_1626)
);

AOI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1609),
.A2(n_1558),
.B(n_1556),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1627),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1620),
.A2(n_1617),
.B1(n_1526),
.B2(n_1517),
.C(n_1507),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1623),
.A2(n_1562),
.B(n_1507),
.C(n_1545),
.Y(n_1630)
);

AOI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1626),
.A2(n_1553),
.B(n_1545),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1619),
.Y(n_1632)
);

OAI21xp33_ASAP7_75t_SL g1633 ( 
.A1(n_1628),
.A2(n_1621),
.B(n_1625),
.Y(n_1633)
);

AOI221xp5_ASAP7_75t_L g1634 ( 
.A1(n_1630),
.A2(n_1622),
.B1(n_1624),
.B2(n_1553),
.C(n_1527),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1632),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1631),
.B(n_1482),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1629),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1632),
.B(n_1512),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1633),
.A2(n_1634),
.B1(n_1637),
.B2(n_1636),
.C(n_1635),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1638),
.B(n_1512),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1633),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1633),
.B(n_1512),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1500),
.Y(n_1643)
);

NAND4xp75_ASAP7_75t_L g1644 ( 
.A(n_1642),
.B(n_1506),
.C(n_1525),
.D(n_1527),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1640),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1641),
.B(n_1479),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1645),
.A2(n_1639),
.B1(n_1643),
.B2(n_1528),
.Y(n_1647)
);

OAI322xp33_ASAP7_75t_L g1648 ( 
.A1(n_1647),
.A2(n_1644),
.A3(n_1646),
.B1(n_1527),
.B2(n_1466),
.C1(n_1464),
.C2(n_1465),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1648),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1648),
.A2(n_1512),
.B(n_1502),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1649),
.Y(n_1651)
);

OAI22x1_ASAP7_75t_L g1652 ( 
.A1(n_1650),
.A2(n_1468),
.B1(n_1528),
.B2(n_1514),
.Y(n_1652)
);

AND2x4_ASAP7_75t_SL g1653 ( 
.A(n_1651),
.B(n_1482),
.Y(n_1653)
);

INVx4_ASAP7_75t_L g1654 ( 
.A(n_1652),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1653),
.B1(n_1514),
.B2(n_1520),
.Y(n_1655)
);

AO21x2_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1520),
.B(n_1519),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1656),
.B(n_1502),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1519),
.B1(n_1469),
.B2(n_1479),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1464),
.B1(n_1465),
.B2(n_1466),
.C(n_1469),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1659),
.A2(n_1328),
.B(n_1468),
.C(n_1466),
.Y(n_1660)
);


endmodule