module real_aes_9203_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_0), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_1), .A2(n_161), .B1(n_298), .B2(n_514), .Y(n_513) );
XOR2x2_ASAP7_75t_L g551 ( .A(n_2), .B(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_3), .A2(n_126), .B1(n_263), .B2(n_266), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_4), .A2(n_42), .B1(n_423), .B2(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g238 ( .A(n_5), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_6), .A2(n_178), .B1(n_348), .B2(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_7), .Y(n_452) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_8), .A2(n_20), .B1(n_168), .B2(n_351), .C1(n_568), .C2(n_570), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_9), .A2(n_131), .B1(n_330), .B2(n_448), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_10), .B(n_251), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_11), .A2(n_53), .B1(n_559), .B2(n_561), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_12), .A2(n_576), .B1(n_600), .B2(n_601), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_12), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_13), .A2(n_45), .B1(n_314), .B2(n_316), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_14), .A2(n_303), .B1(n_368), .B2(n_369), .Y(n_302) );
INVx1_ASAP7_75t_L g368 ( .A(n_14), .Y(n_368) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_15), .B(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_16), .A2(n_206), .B1(n_428), .B2(n_470), .Y(n_617) );
INVx1_ASAP7_75t_L g475 ( .A(n_17), .Y(n_475) );
AO22x2_ASAP7_75t_L g227 ( .A1(n_18), .A2(n_60), .B1(n_228), .B2(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g641 ( .A(n_18), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_19), .A2(n_110), .B1(n_315), .B2(n_333), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_21), .Y(n_300) );
AOI222xp33_ASAP7_75t_L g450 ( .A1(n_22), .A2(n_66), .B1(n_189), .B2(n_224), .C1(n_246), .C2(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_23), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_24), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_25), .A2(n_136), .B1(n_246), .B2(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_26), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_27), .A2(n_36), .B1(n_381), .B2(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_28), .A2(n_29), .B1(n_251), .B2(n_468), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_30), .A2(n_156), .B1(n_293), .B2(n_448), .Y(n_456) );
AO22x2_ASAP7_75t_L g231 ( .A1(n_31), .A2(n_62), .B1(n_228), .B2(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g642 ( .A(n_31), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_32), .A2(n_98), .B1(n_295), .B2(n_298), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_33), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_34), .A2(n_52), .B1(n_431), .B2(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_35), .A2(n_149), .B1(n_381), .B2(n_382), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_37), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_38), .B(n_468), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_39), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_40), .A2(n_67), .B1(n_329), .B2(n_331), .Y(n_328) );
AOI22xp5_ASAP7_75t_SL g457 ( .A1(n_41), .A2(n_192), .B1(n_458), .B2(n_460), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_43), .A2(n_174), .B1(n_326), .B2(n_418), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_44), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_46), .B(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_47), .A2(n_195), .B1(n_240), .B2(n_246), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_48), .B(n_257), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_49), .A2(n_190), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_50), .A2(n_155), .B1(n_281), .B2(n_330), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_51), .B(n_423), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_54), .A2(n_137), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_55), .A2(n_114), .B1(n_355), .B2(n_428), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_56), .A2(n_72), .B1(n_311), .B2(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_57), .A2(n_88), .B1(n_415), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_58), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_59), .A2(n_197), .B1(n_252), .B2(n_422), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_61), .A2(n_128), .B1(n_266), .B2(n_426), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_63), .A2(n_194), .B1(n_284), .B2(n_415), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_64), .A2(n_154), .B1(n_413), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_65), .A2(n_163), .B1(n_288), .B2(n_315), .Y(n_658) );
INVx1_ASAP7_75t_L g214 ( .A(n_68), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_69), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_70), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_71), .A2(n_139), .B1(n_311), .B2(n_565), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_73), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g211 ( .A(n_74), .Y(n_211) );
INVx1_ASAP7_75t_L g478 ( .A(n_75), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_76), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_77), .A2(n_105), .B1(n_288), .B2(n_291), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_78), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_79), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_80), .A2(n_125), .B1(n_290), .B2(n_330), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_81), .A2(n_143), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_82), .A2(n_90), .B1(n_311), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_83), .A2(n_175), .B1(n_317), .B2(n_448), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_84), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_85), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_86), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_87), .A2(n_150), .B1(n_514), .B2(n_597), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_89), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_91), .A2(n_95), .B1(n_348), .B2(n_445), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_92), .A2(n_162), .B1(n_331), .B2(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_93), .A2(n_485), .B1(n_486), .B2(n_518), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_93), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_94), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_96), .A2(n_201), .B1(n_288), .B2(n_565), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_97), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_99), .A2(n_124), .B1(n_417), .B2(n_418), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_100), .A2(n_127), .B1(n_157), .B2(n_225), .C1(n_240), .C2(n_399), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_101), .A2(n_188), .B1(n_470), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_102), .A2(n_147), .B1(n_544), .B2(n_545), .Y(n_543) );
AOI22x1_ASAP7_75t_L g373 ( .A1(n_103), .A2(n_374), .B1(n_404), .B2(n_405), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_103), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_104), .A2(n_177), .B1(n_314), .B2(n_460), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_106), .Y(n_349) );
INVx2_ASAP7_75t_L g215 ( .A(n_107), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_108), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_109), .A2(n_179), .B1(n_355), .B2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_111), .A2(n_138), .B1(n_385), .B2(n_465), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_112), .A2(n_645), .B1(n_646), .B2(n_663), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_112), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_113), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_115), .A2(n_180), .B1(n_426), .B2(n_428), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_116), .A2(n_167), .B1(n_434), .B2(n_548), .Y(n_547) );
AND2x6_ASAP7_75t_L g210 ( .A(n_117), .B(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_117), .Y(n_635) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_118), .A2(n_172), .B1(n_228), .B2(n_232), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_119), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_120), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_121), .A2(n_173), .B1(n_593), .B2(n_594), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_122), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_123), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_129), .A2(n_152), .B1(n_501), .B2(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_130), .A2(n_191), .B1(n_463), .B2(n_516), .Y(n_624) );
INVx1_ASAP7_75t_L g673 ( .A(n_132), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_133), .A2(n_198), .B1(n_272), .B2(n_431), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_134), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_135), .A2(n_165), .B1(n_314), .B2(n_316), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_140), .A2(n_169), .B1(n_284), .B2(n_559), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_141), .B(n_251), .Y(n_654) );
AO22x2_ASAP7_75t_L g237 ( .A1(n_142), .A2(n_181), .B1(n_228), .B2(n_229), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g271 ( .A1(n_144), .A2(n_185), .B1(n_272), .B2(n_276), .Y(n_271) );
XOR2x2_ASAP7_75t_L g408 ( .A(n_145), .B(n_409), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_146), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_148), .A2(n_151), .B1(n_281), .B2(n_284), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_153), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_158), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_159), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_160), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_164), .A2(n_204), .B1(n_240), .B2(n_263), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_166), .A2(n_208), .B(n_216), .C(n_643), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_170), .A2(n_203), .B1(n_314), .B2(n_316), .Y(n_313) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_171), .B(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_172), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_176), .A2(n_183), .B1(n_433), .B2(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g638 ( .A(n_181), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_182), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_184), .A2(n_205), .B1(n_421), .B2(n_423), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_186), .Y(n_378) );
INVx1_ASAP7_75t_L g608 ( .A(n_187), .Y(n_608) );
INVx1_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
INVx1_ASAP7_75t_L g230 ( .A(n_193), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_196), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_199), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_200), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_202), .Y(n_491) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_210), .B(n_212), .Y(n_209) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_211), .Y(n_634) );
OA21x2_ASAP7_75t_L g671 ( .A1(n_212), .A2(n_633), .B(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_215), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_481), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_216) );
INVx1_ASAP7_75t_L g628 ( .A(n_217), .Y(n_628) );
XNOR2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_371), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_301), .B1(n_302), .B2(n_370), .Y(n_218) );
INVx3_ASAP7_75t_SL g370 ( .A(n_219), .Y(n_370) );
XOR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_300), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_269), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_249), .Y(n_221) );
OAI21xp5_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_238), .B(n_239), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_225), .Y(n_351) );
INVx4_ASAP7_75t_L g474 ( .A(n_225), .Y(n_474) );
INVx2_ASAP7_75t_SL g525 ( .A(n_225), .Y(n_525) );
INVx2_ASAP7_75t_L g649 ( .A(n_225), .Y(n_649) );
AND2x6_ASAP7_75t_L g225 ( .A(n_226), .B(n_233), .Y(n_225) );
AND2x4_ASAP7_75t_L g266 ( .A(n_226), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g366 ( .A(n_226), .Y(n_366) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
AND2x2_ASAP7_75t_L g245 ( .A(n_227), .B(n_235), .Y(n_245) );
INVx2_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_230), .Y(n_232) );
INVx2_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
AND2x2_ASAP7_75t_L g253 ( .A(n_231), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g261 ( .A(n_231), .B(n_254), .Y(n_261) );
INVx1_ASAP7_75t_L g265 ( .A(n_231), .Y(n_265) );
AND2x6_ASAP7_75t_L g290 ( .A(n_233), .B(n_260), .Y(n_290) );
AND2x4_ASAP7_75t_L g293 ( .A(n_233), .B(n_253), .Y(n_293) );
AND2x2_ASAP7_75t_L g297 ( .A(n_233), .B(n_275), .Y(n_297) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g255 ( .A(n_234), .B(n_237), .Y(n_255) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g274 ( .A(n_235), .B(n_268), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_235), .B(n_237), .Y(n_279) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g243 ( .A(n_237), .Y(n_243) );
INVx1_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
INVx1_ASAP7_75t_L g395 ( .A(n_240), .Y(n_395) );
BUFx4f_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_241), .Y(n_348) );
BUFx2_ASAP7_75t_L g477 ( .A(n_241), .Y(n_477) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_241), .Y(n_536) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_241), .Y(n_612) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g248 ( .A(n_243), .Y(n_248) );
AND2x2_ASAP7_75t_L g275 ( .A(n_244), .B(n_254), .Y(n_275) );
INVx1_ASAP7_75t_L g285 ( .A(n_244), .Y(n_285) );
AND2x4_ASAP7_75t_L g247 ( .A(n_245), .B(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g263 ( .A(n_245), .B(n_264), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_245), .B(n_285), .Y(n_361) );
BUFx4f_ASAP7_75t_SL g399 ( .A(n_246), .Y(n_399) );
INVx2_ASAP7_75t_L g569 ( .A(n_246), .Y(n_569) );
BUFx12f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_247), .Y(n_355) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_247), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_256), .C(n_262), .Y(n_249) );
BUFx4f_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_SL g424 ( .A(n_252), .Y(n_424) );
BUFx2_ASAP7_75t_L g534 ( .A(n_252), .Y(n_534) );
AND2x6_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g283 ( .A(n_253), .B(n_274), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_253), .B(n_255), .Y(n_344) );
AND2x4_ASAP7_75t_L g259 ( .A(n_255), .B(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g299 ( .A(n_255), .B(n_275), .Y(n_299) );
INVx1_ASAP7_75t_L g340 ( .A(n_255), .Y(n_340) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx5_ASAP7_75t_L g422 ( .A(n_258), .Y(n_422) );
INVx2_ASAP7_75t_L g468 ( .A(n_258), .Y(n_468) );
INVx2_ASAP7_75t_L g616 ( .A(n_258), .Y(n_616) );
INVx4_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g339 ( .A(n_261), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g427 ( .A(n_263), .Y(n_427) );
BUFx3_ASAP7_75t_L g445 ( .A(n_263), .Y(n_445) );
BUFx2_ASAP7_75t_L g470 ( .A(n_263), .Y(n_470) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x6_ASAP7_75t_L g318 ( .A(n_265), .B(n_279), .Y(n_318) );
BUFx2_ASAP7_75t_SL g428 ( .A(n_266), .Y(n_428) );
BUFx3_ASAP7_75t_L g451 ( .A(n_266), .Y(n_451) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_266), .Y(n_471) );
BUFx2_ASAP7_75t_SL g570 ( .A(n_266), .Y(n_570) );
INVx1_ASAP7_75t_L g367 ( .A(n_267), .Y(n_367) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_286), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_280), .Y(n_270) );
BUFx2_ASAP7_75t_L g599 ( .A(n_272), .Y(n_599) );
BUFx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx3_ASAP7_75t_L g448 ( .A(n_273), .Y(n_448) );
BUFx3_ASAP7_75t_L g542 ( .A(n_273), .Y(n_542) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_274), .B(n_275), .Y(n_308) );
AND2x4_ASAP7_75t_L g277 ( .A(n_275), .B(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx3_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
BUFx3_ASAP7_75t_L g431 ( .A(n_277), .Y(n_431) );
BUFx2_ASAP7_75t_SL g465 ( .A(n_277), .Y(n_465) );
BUFx3_ASAP7_75t_L g545 ( .A(n_277), .Y(n_545) );
INVx1_ASAP7_75t_L g562 ( .A(n_277), .Y(n_562) );
AND2x2_ASAP7_75t_L g284 ( .A(n_278), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx5_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
INVx4_ASAP7_75t_L g459 ( .A(n_282), .Y(n_459) );
BUFx3_ASAP7_75t_L g549 ( .A(n_282), .Y(n_549) );
INVx3_ASAP7_75t_L g593 ( .A(n_282), .Y(n_593) );
INVx8_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_294), .Y(n_286) );
INVx4_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g510 ( .A(n_289), .Y(n_510) );
INVx11_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx11_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g385 ( .A(n_292), .Y(n_385) );
INVx2_ASAP7_75t_L g434 ( .A(n_292), .Y(n_434) );
INVx2_ASAP7_75t_L g597 ( .A(n_292), .Y(n_597) );
INVx6_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx3_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
BUFx3_ASAP7_75t_L g565 ( .A(n_293), .Y(n_565) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g544 ( .A(n_296), .Y(n_544) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
BUFx2_ASAP7_75t_SL g412 ( .A(n_297), .Y(n_412) );
BUFx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_299), .Y(n_415) );
INVx2_ASAP7_75t_L g560 ( .A(n_299), .Y(n_560) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_334), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_319), .Y(n_304) );
OAI221xp5_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_309), .B1(n_310), .B2(n_312), .C(n_313), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g387 ( .A(n_307), .Y(n_387) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_311), .Y(n_382) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_315), .Y(n_417) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
BUFx2_ASAP7_75t_L g460 ( .A(n_317), .Y(n_460) );
INVx6_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g594 ( .A(n_318), .Y(n_594) );
OAI221xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_323), .B1(n_324), .B2(n_327), .C(n_328), .Y(n_319) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_320), .A2(n_414), .B1(n_590), .B2(n_591), .C(n_592), .Y(n_589) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx1_ASAP7_75t_L g433 ( .A(n_322), .Y(n_433) );
INVx2_ASAP7_75t_SL g540 ( .A(n_322), .Y(n_540) );
OAI221xp5_ASAP7_75t_SL g376 ( .A1(n_324), .A2(n_377), .B1(n_378), .B2(n_379), .C(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_330), .Y(n_463) );
BUFx3_ASAP7_75t_L g514 ( .A(n_330), .Y(n_514) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_345), .C(n_357), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_341), .B2(n_342), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_337), .A2(n_342), .B1(n_392), .B2(n_393), .Y(n_391) );
OAI221xp5_ASAP7_75t_SL g578 ( .A1(n_337), .A2(n_579), .B1(n_580), .B2(n_581), .C(n_582), .Y(n_578) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g490 ( .A(n_338), .Y(n_490) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g580 ( .A(n_343), .Y(n_580) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g494 ( .A(n_344), .Y(n_494) );
OAI222xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_350), .B2(n_352), .C1(n_353), .C2(n_356), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g495 ( .A1(n_346), .A2(n_496), .B1(n_498), .B2(n_499), .C(n_500), .Y(n_495) );
INVx2_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI222xp33_ASAP7_75t_L g394 ( .A1(n_350), .A2(n_395), .B1(n_396), .B2(n_397), .C1(n_398), .C2(n_400), .Y(n_394) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_362), .B2(n_363), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_359), .A2(n_363), .B1(n_402), .B2(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx4_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g504 ( .A(n_361), .Y(n_504) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g506 ( .A(n_364), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_365), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_406), .B2(n_480), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_375), .B(n_390), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_383), .Y(n_375) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_386), .B1(n_387), .B2(n_388), .C(n_389), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_394), .C(n_401), .Y(n_390) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_398), .A2(n_496), .B1(n_584), .B2(n_585), .C1(n_586), .C2(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g480 ( .A(n_406), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_436), .B2(n_479), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND4xp75_ASAP7_75t_L g409 ( .A(n_410), .B(n_419), .C(n_429), .D(n_435), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_416), .Y(n_410) );
INVx4_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_420), .B(n_425), .Y(n_419) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_422), .Y(n_532) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_453), .Y(n_436) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_452), .Y(n_437) );
NAND4xp75_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .C(n_446), .D(n_450), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_443), .B(n_444), .Y(n_442) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g517 ( .A(n_448), .Y(n_517) );
XOR2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_478), .Y(n_453) );
NOR4xp75_ASAP7_75t_L g454 ( .A(n_455), .B(n_461), .C(n_466), .D(n_472), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_456), .B(n_457), .Y(n_455) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx1_ASAP7_75t_SL g529 ( .A(n_471), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_475), .B(n_476), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g497 ( .A(n_474), .Y(n_497) );
INVx1_ASAP7_75t_L g629 ( .A(n_481), .Y(n_629) );
XOR2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_572), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_519), .B1(n_520), .B2(n_571), .Y(n_482) );
INVx1_ASAP7_75t_L g571 ( .A(n_483), .Y(n_571) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_507), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_495), .C(n_502), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_488) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_496), .A2(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
XOR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_551), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_537), .Y(n_522) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_524), .B(n_530), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_525), .A2(n_526), .B(n_527), .Y(n_524) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .C(n_535), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_536), .Y(n_584) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_538), .B(n_546), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
INVx1_ASAP7_75t_L g621 ( .A(n_540), .Y(n_621) );
BUFx4f_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .Y(n_546) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND4xp75_ASAP7_75t_L g552 ( .A(n_553), .B(n_556), .C(n_563), .D(n_567), .Y(n_552) );
AND2x2_ASAP7_75t_SL g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_602), .B1(n_626), .B2(n_627), .Y(n_573) );
INVx1_ASAP7_75t_L g626 ( .A(n_574), .Y(n_626) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g601 ( .A(n_576), .Y(n_601) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_588), .Y(n_576) );
NOR2xp33_ASAP7_75t_SL g577 ( .A(n_578), .B(n_583), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_595), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g627 ( .A(n_602), .Y(n_627) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND3x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_618), .C(n_623), .Y(n_605) );
NOR2x1_ASAP7_75t_SL g606 ( .A(n_607), .B(n_613), .Y(n_606) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx4_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .C(n_617), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NOR2x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
OR2x2_ASAP7_75t_SL g679 ( .A(n_632), .B(n_637), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_633), .Y(n_665) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_634), .B(n_668), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g668 ( .A(n_635), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OAI322xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_664), .A3(n_666), .B1(n_669), .B2(n_673), .C1(n_674), .C2(n_677), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
XOR2x2_ASAP7_75t_L g676 ( .A(n_646), .B(n_673), .Y(n_676) );
NAND2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_656), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .C(n_655), .Y(n_652) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
endmodule