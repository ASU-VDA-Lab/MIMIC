module fake_jpeg_14295_n_188 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_29),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_63),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_41),
.B(n_45),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_9),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_51),
.Y(n_94)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_52),
.B(n_55),
.Y(n_96)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_13),
.B(n_4),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_58),
.Y(n_90)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_20),
.B1(n_33),
.B2(n_27),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_74),
.B1(n_91),
.B2(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_35),
.B1(n_33),
.B2(n_27),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_95),
.B1(n_66),
.B2(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_72)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_87),
.B(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_28),
.B1(n_5),
.B2(n_7),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_36),
.A2(n_28),
.B1(n_4),
.B2(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_99),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_53),
.B(n_36),
.C(n_60),
.Y(n_91)
);

AO21x1_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_79),
.B(n_80),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_65),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_49),
.B1(n_59),
.B2(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_37),
.B(n_38),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_103),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_112),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_61),
.B(n_43),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_111),
.B(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_123),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_122),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_78),
.B(n_95),
.C(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_78),
.B1(n_68),
.B2(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_124),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_86),
.B1(n_69),
.B2(n_89),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_78),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_109),
.B(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.C(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_106),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_114),
.B(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_125),
.B1(n_118),
.B2(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_136),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_111),
.B(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_123),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_153),
.Y(n_165)
);

BUFx12f_ASAP7_75t_SL g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_138),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_138),
.Y(n_155)
);

BUFx12f_ASAP7_75t_SL g156 ( 
.A(n_139),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_135),
.C(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_164),
.C(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_140),
.B1(n_136),
.B2(n_126),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_151),
.C(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_168),
.C(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_155),
.C(n_156),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_150),
.B(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_163),
.B1(n_160),
.B2(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_162),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_177),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_144),
.A3(n_142),
.B1(n_148),
.B2(n_132),
.C1(n_137),
.C2(n_130),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_120),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_177),
.Y(n_182)
);

OAI21x1_ASAP7_75t_SL g185 ( 
.A1(n_182),
.A2(n_184),
.B(n_179),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_175),
.B(n_132),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_186),
.C(n_117),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_132),
.B(n_130),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_108),
.Y(n_188)
);


endmodule