module fake_netlist_5_2254_n_1794 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1794);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1794;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_6),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_28),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_61),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_52),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_36),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_130),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_103),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_94),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_65),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_21),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_51),
.Y(n_195)
);

INVx4_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_39),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_29),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_82),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_90),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_48),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_151),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_25),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_128),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_87),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_44),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_5),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_42),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_20),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_139),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_95),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_4),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_96),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_44),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_93),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_76),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_40),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_9),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_155),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_89),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_117),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_74),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_35),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_72),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_68),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_92),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_125),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_23),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_153),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_75),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_7),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_116),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_42),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_22),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_154),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_83),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_84),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_109),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_160),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_67),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_142),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_50),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_169),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_156),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_49),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_38),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_152),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_73),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_2),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_133),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_108),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_37),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_141),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_26),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_105),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_80),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_1),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_4),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_166),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_144),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_17),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_26),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_122),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_131),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_36),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_33),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_30),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_8),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_140),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_135),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_101),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_104),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_9),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_31),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_137),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_32),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_162),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_23),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_120),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_50),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_17),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_63),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_34),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_98),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_14),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_27),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_7),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_37),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_123),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_148),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_121),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_97),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_159),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_33),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_157),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_43),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_106),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_27),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_40),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_85),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_12),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_10),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_10),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_127),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_32),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_118),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_24),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_39),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_79),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_178),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_236),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_211),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_179),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_179),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_236),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_269),
.B(n_3),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_175),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_179),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_179),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_197),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_179),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_179),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_200),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_253),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_212),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_179),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_260),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_260),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_243),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_182),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_202),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_260),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_205),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_208),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_240),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_209),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_3),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_253),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_260),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_260),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_213),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_262),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_332),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_262),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_271),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_260),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_271),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_260),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_225),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_296),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_182),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_225),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_210),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_177),
.B(n_8),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_319),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_214),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_220),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_225),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_184),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_221),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_225),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_224),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_226),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_227),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_235),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_235),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_233),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_235),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_235),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_263),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_296),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_263),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_263),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_234),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_263),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_239),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_311),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_269),
.B(n_12),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_244),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_184),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_192),
.B(n_13),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_311),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_247),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_311),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_311),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_248),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_250),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_212),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_335),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_251),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_256),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_335),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_177),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_R g435 ( 
.A(n_346),
.B(n_257),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_349),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_406),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_358),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_361),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_369),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_371),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_331),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_192),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_347),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_363),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_355),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_363),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_372),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_374),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_367),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_404),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_363),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_379),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_394),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_395),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_363),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_368),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_426),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_172),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_398),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_400),
.B(n_401),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_426),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_402),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_405),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_412),
.B(n_261),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_427),
.B(n_305),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_414),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_381),
.B(n_391),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_410),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_417),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_421),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_352),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_425),
.B(n_266),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_428),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_420),
.B(n_305),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_353),
.A2(n_306),
.B(n_180),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_422),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_429),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_362),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_422),
.B(n_172),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_430),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_376),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_430),
.Y(n_511)
);

AND3x2_ASAP7_75t_L g512 ( 
.A(n_442),
.B(n_375),
.C(n_419),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_484),
.B(n_373),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_484),
.B(n_418),
.C(n_416),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_472),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_461),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_476),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_316),
.B1(n_337),
.B2(n_199),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

INVx4_ASAP7_75t_SL g527 ( 
.A(n_472),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_448),
.B(n_306),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_454),
.B(n_431),
.Y(n_531)
);

NOR2x1p5_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_439),
.Y(n_532)
);

AND2x2_ASAP7_75t_SL g533 ( 
.A(n_454),
.B(n_212),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_474),
.B(n_373),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_448),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_441),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_SL g537 ( 
.A(n_501),
.B(n_316),
.C(n_199),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_454),
.B(n_431),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_474),
.B(n_424),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_442),
.B(n_424),
.C(n_348),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_432),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_444),
.A2(n_445),
.B1(n_460),
.B2(n_459),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_482),
.B(n_212),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_482),
.B(n_432),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_446),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_503),
.A2(n_195),
.B1(n_270),
.B2(n_281),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_470),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_446),
.B(n_331),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_447),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_447),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_482),
.B(n_457),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_434),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_457),
.B(n_246),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_450),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_451),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_457),
.B(n_507),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_507),
.B(n_350),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_502),
.B(n_246),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_465),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_451),
.B(n_452),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_350),
.Y(n_565)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_502),
.B(n_246),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_494),
.B(n_302),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_453),
.B(n_351),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_503),
.A2(n_281),
.B1(n_313),
.B2(n_270),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_503),
.A2(n_195),
.B1(n_313),
.B2(n_392),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_462),
.B(n_302),
.Y(n_571)
);

AND2x2_ASAP7_75t_SL g572 ( 
.A(n_502),
.B(n_246),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_464),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_440),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_466),
.B(n_279),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_478),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_467),
.B(n_337),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_478),
.B(n_201),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_502),
.B(n_279),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_485),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_475),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_440),
.B(n_215),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_351),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_440),
.B(n_433),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_440),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_486),
.B(n_356),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_511),
.A2(n_259),
.B1(n_217),
.B2(n_249),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_487),
.B(n_356),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_487),
.A2(n_252),
.B1(n_315),
.B2(n_318),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_489),
.B(n_357),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_480),
.B(n_279),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_483),
.B(n_433),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_481),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_492),
.B(n_309),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_511),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_492),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_493),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_493),
.B(n_357),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_477),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_499),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_498),
.B(n_359),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_504),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_508),
.B(n_359),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_SL g619 ( 
.A1(n_508),
.A2(n_364),
.B(n_360),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_434),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_497),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_506),
.B(n_320),
.C(n_204),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_434),
.B(n_324),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_495),
.B(n_279),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_500),
.B(n_173),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_505),
.B(n_183),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_434),
.B(n_360),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_477),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_477),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_477),
.B(n_188),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_449),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_449),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_477),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_456),
.A2(n_272),
.B1(n_329),
.B2(n_254),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_456),
.B(n_273),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_510),
.B(n_365),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_458),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_458),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_458),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_463),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_463),
.B(n_365),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_509),
.A2(n_278),
.B1(n_218),
.B2(n_230),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_463),
.B(n_338),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_468),
.B(n_366),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_468),
.B(n_366),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_477),
.B(n_190),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_468),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_469),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_469),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_469),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_510),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_490),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_490),
.B(n_370),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_491),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_491),
.A2(n_293),
.B1(n_288),
.B2(n_341),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_491),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_438),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_523),
.B(n_191),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_513),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_518),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_517),
.Y(n_663)
);

BUFx12f_ASAP7_75t_SL g664 ( 
.A(n_599),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_520),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_535),
.B(n_183),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_526),
.B(n_185),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_593),
.B(n_185),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_644),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_533),
.B(n_193),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_519),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_533),
.B(n_207),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_608),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_561),
.B(n_216),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_603),
.B(n_380),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_574),
.B(n_289),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_554),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_521),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_534),
.B(n_187),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_544),
.B(n_222),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_544),
.B(n_237),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_531),
.A2(n_370),
.B(n_386),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_534),
.B(n_382),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_636),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_539),
.B(n_187),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_566),
.B(n_572),
.Y(n_686)
);

NOR3xp33_ASAP7_75t_L g687 ( 
.A(n_537),
.B(n_242),
.C(n_255),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_539),
.A2(n_619),
.B(n_571),
.C(n_542),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_570),
.A2(n_241),
.B1(n_342),
.B2(n_328),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_566),
.B(n_258),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_572),
.B(n_265),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_514),
.B(n_189),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_608),
.Y(n_693)
);

AOI221xp5_ASAP7_75t_L g694 ( 
.A1(n_524),
.A2(n_344),
.B1(n_339),
.B2(n_338),
.C(n_298),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_514),
.B(n_515),
.Y(n_695)
);

OR2x6_ASAP7_75t_L g696 ( 
.A(n_595),
.B(n_300),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_549),
.A2(n_343),
.B1(n_386),
.B2(n_384),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_607),
.B(n_268),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_625),
.B(n_548),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_530),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_625),
.B(n_189),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_607),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_549),
.A2(n_377),
.B1(n_384),
.B2(n_378),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_604),
.B(n_336),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_538),
.B(n_274),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_530),
.A2(n_409),
.B1(n_388),
.B2(n_385),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_567),
.B(n_336),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_547),
.B(n_282),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_636),
.Y(n_709)
);

OAI22x1_ASAP7_75t_SL g710 ( 
.A1(n_525),
.A2(n_383),
.B1(n_339),
.B2(n_344),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_528),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_536),
.B(n_297),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_569),
.A2(n_570),
.B1(n_530),
.B2(n_634),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_540),
.B(n_301),
.Y(n_714)
);

A2O1A1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_571),
.A2(n_378),
.B(n_377),
.C(n_303),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_567),
.B(n_340),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_584),
.A2(n_203),
.B1(n_275),
.B2(n_334),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_550),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_546),
.B(n_304),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_552),
.B(n_310),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_553),
.B(n_325),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_575),
.B(n_586),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_555),
.B(n_326),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_569),
.A2(n_340),
.B1(n_345),
.B2(n_330),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_578),
.B(n_174),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_558),
.B(n_277),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_606),
.B(n_211),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_559),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_573),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_280),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_580),
.B(n_285),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_578),
.B(n_176),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_581),
.B(n_286),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_530),
.A2(n_290),
.B1(n_327),
.B2(n_307),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_530),
.A2(n_312),
.B1(n_314),
.B2(n_317),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_649),
.A2(n_333),
.B1(n_186),
.B2(n_231),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_582),
.B(n_194),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_623),
.B(n_186),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_634),
.A2(n_211),
.B1(n_323),
.B2(n_322),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_657),
.A2(n_597),
.B1(n_600),
.B2(n_545),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_198),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_605),
.B(n_206),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_609),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_545),
.A2(n_196),
.B(n_321),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_611),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_623),
.B(n_219),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_602),
.B(n_267),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_643),
.B(n_524),
.C(n_541),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_615),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_613),
.A2(n_276),
.B1(n_308),
.B2(n_299),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_624),
.B(n_245),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_624),
.B(n_333),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_577),
.B(n_223),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_583),
.B(n_228),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_583),
.B(n_283),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_SL g756 ( 
.A(n_599),
.B(n_333),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_295),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_294),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_519),
.B(n_551),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_626),
.B(n_292),
.C(n_287),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_590),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_551),
.B(n_238),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_512),
.B(n_232),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_590),
.B(n_229),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_284),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_616),
.B(n_284),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_L g767 ( 
.A(n_562),
.B(n_284),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_657),
.A2(n_264),
.B1(n_231),
.B2(n_186),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_512),
.B(n_264),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_617),
.B(n_264),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_659),
.B(n_231),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_659),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_616),
.B(n_15),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_655),
.B(n_556),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_591),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_564),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_591),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_591),
.B(n_15),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_522),
.B(n_16),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_522),
.B(n_16),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_637),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_631),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_563),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_622),
.B(n_18),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_598),
.B(n_610),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_650),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_598),
.B(n_62),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_648),
.B(n_60),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_543),
.B(n_19),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_69),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_621),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_650),
.B(n_19),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_642),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_618),
.B(n_77),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_648),
.B(n_59),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_557),
.A2(n_78),
.B1(n_161),
.B2(n_150),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_618),
.B(n_57),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_562),
.B(n_58),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_557),
.A2(n_55),
.B1(n_145),
.B2(n_138),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_645),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_627),
.B(n_646),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_565),
.B(n_20),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_648),
.B(n_164),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_532),
.B(n_24),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_641),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_627),
.B(n_136),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_563),
.B(n_28),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_589),
.B(n_29),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_589),
.Y(n_810)
);

AND2x6_ASAP7_75t_SL g811 ( 
.A(n_568),
.B(n_31),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_592),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_597),
.B(n_41),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_646),
.B(n_81),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_596),
.B(n_601),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_614),
.B(n_86),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_630),
.B(n_119),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_656),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_620),
.B(n_115),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_648),
.B(n_639),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_786),
.A2(n_585),
.B(n_529),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_786),
.A2(n_585),
.B(n_529),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_677),
.A2(n_585),
.B(n_529),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_718),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_688),
.A2(n_647),
.B(n_630),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_815),
.A2(n_529),
.B(n_585),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_679),
.A2(n_638),
.B(n_654),
.C(n_653),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_713),
.A2(n_647),
.B(n_652),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_679),
.A2(n_651),
.B(n_635),
.C(n_632),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_684),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_684),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_785),
.B(n_640),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_709),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_761),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_722),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_678),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_713),
.A2(n_628),
.B(n_612),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_801),
.A2(n_594),
.B(n_576),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_686),
.A2(n_594),
.B(n_576),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_772),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_776),
.B(n_812),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_663),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_810),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_671),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_689),
.A2(n_600),
.B(n_629),
.C(n_562),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_700),
.A2(n_612),
.B(n_628),
.Y(n_846)
);

AO21x1_ASAP7_75t_L g847 ( 
.A1(n_787),
.A2(n_562),
.B(n_587),
.Y(n_847)
);

INVx3_ASAP7_75t_SL g848 ( 
.A(n_783),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_704),
.B(n_99),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_667),
.B(n_629),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_727),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_707),
.B(n_41),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_671),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_667),
.B(n_628),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_778),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_699),
.B(n_612),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_707),
.A2(n_658),
.B(n_633),
.C(n_516),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_716),
.B(n_45),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_817),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_716),
.B(n_45),
.Y(n_860)
);

O2A1O1Ixp5_ASAP7_75t_L g861 ( 
.A1(n_691),
.A2(n_587),
.B(n_527),
.C(n_658),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_700),
.A2(n_633),
.B(n_516),
.Y(n_862)
);

AOI21x1_ASAP7_75t_L g863 ( 
.A1(n_820),
.A2(n_527),
.B(n_658),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_817),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_664),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_700),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_791),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_775),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_701),
.A2(n_658),
.B(n_633),
.C(n_516),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_669),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_699),
.B(n_633),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_781),
.A2(n_516),
.B(n_102),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_740),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_704),
.B(n_47),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_695),
.B(n_49),
.Y(n_875)
);

NAND2x1_ASAP7_75t_L g876 ( 
.A(n_818),
.B(n_100),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_774),
.A2(n_52),
.B(n_53),
.Y(n_877)
);

AO22x1_ASAP7_75t_L g878 ( 
.A1(n_789),
.A2(n_54),
.B1(n_813),
.B2(n_748),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_683),
.B(n_54),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_793),
.A2(n_800),
.B(n_697),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_702),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_774),
.A2(n_681),
.B(n_680),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_759),
.A2(n_703),
.B(n_794),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_660),
.B(n_740),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_673),
.B(n_693),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_759),
.A2(n_703),
.B(n_790),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_797),
.A2(n_806),
.B(n_814),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_775),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_789),
.B(n_756),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_728),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_816),
.A2(n_697),
.B(n_705),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_775),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_746),
.B(n_777),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_708),
.A2(n_672),
.B(n_733),
.Y(n_894)
);

NAND2xp33_ASAP7_75t_L g895 ( 
.A(n_690),
.B(n_674),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_706),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_729),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_743),
.B(n_745),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_726),
.A2(n_730),
.B(n_731),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_749),
.B(n_661),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_662),
.B(n_665),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_676),
.B(n_696),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_675),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_701),
.B(n_725),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_692),
.B(n_762),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_698),
.A2(n_803),
.B(n_795),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_788),
.A2(n_803),
.B(n_795),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_692),
.A2(n_747),
.B1(n_732),
.B2(n_751),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_782),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_685),
.B(n_668),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_725),
.B(n_732),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_741),
.B(n_751),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_788),
.B(n_796),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_741),
.B(n_747),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_802),
.A2(n_691),
.B1(n_792),
.B2(n_768),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_762),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_819),
.A2(n_682),
.B(n_753),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_715),
.A2(n_802),
.B(n_792),
.C(n_724),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_754),
.B(n_757),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_755),
.B(n_758),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_694),
.B(n_768),
.C(n_687),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_738),
.A2(n_773),
.B(n_737),
.C(n_742),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_764),
.B(n_720),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_763),
.B(n_769),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_750),
.B(n_760),
.C(n_739),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_805),
.A2(n_808),
.B(n_798),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_712),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_714),
.B(n_723),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_SL g929 ( 
.A1(n_738),
.A2(n_752),
.B(n_784),
.C(n_780),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_719),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_721),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_765),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_807),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_770),
.B(n_771),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_804),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_744),
.A2(n_767),
.B(n_666),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_676),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_717),
.A2(n_779),
.B(n_766),
.C(n_763),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_717),
.A2(n_779),
.B(n_769),
.C(n_676),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_696),
.B(n_736),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_804),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_734),
.A2(n_735),
.B(n_799),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_739),
.A2(n_804),
.B(n_809),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_809),
.A2(n_710),
.B(n_811),
.Y(n_944)
);

AOI21x1_ASAP7_75t_L g945 ( 
.A1(n_809),
.A2(n_820),
.B(n_774),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_688),
.A2(n_713),
.B(n_677),
.Y(n_946)
);

CKINVDCx10_ASAP7_75t_R g947 ( 
.A(n_809),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_671),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_695),
.A2(n_699),
.B1(n_679),
.B2(n_776),
.Y(n_949)
);

O2A1O1Ixp5_ASAP7_75t_L g950 ( 
.A1(n_691),
.A2(n_681),
.B(n_680),
.C(n_670),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_722),
.B(n_525),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_785),
.B(n_776),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_718),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_722),
.B(n_484),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_713),
.B(n_699),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_684),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_688),
.A2(n_689),
.B(n_672),
.C(n_670),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_785),
.B(n_776),
.Y(n_961)
);

CKINVDCx10_ASAP7_75t_R g962 ( 
.A(n_809),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_722),
.B(n_347),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_785),
.B(n_776),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_691),
.A2(n_681),
.B(n_680),
.C(n_670),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_820),
.A2(n_774),
.B(n_787),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_691),
.A2(n_681),
.B(n_680),
.C(n_670),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_789),
.A2(n_813),
.B1(n_707),
.B2(n_716),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_671),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_718),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_775),
.B(n_783),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_785),
.B(n_776),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_688),
.A2(n_689),
.B(n_672),
.C(n_670),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_713),
.A2(n_740),
.B1(n_785),
.B2(n_697),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_684),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_785),
.B(n_776),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_678),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_688),
.A2(n_713),
.B(n_677),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_785),
.B(n_776),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_783),
.B(n_574),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_785),
.B(n_776),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_785),
.B(n_776),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_722),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_786),
.A2(n_544),
.B(n_677),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_785),
.B(n_776),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_713),
.B(n_699),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_785),
.B(n_776),
.Y(n_992)
);

AOI211xp5_ASAP7_75t_L g993 ( 
.A1(n_717),
.A2(n_524),
.B(n_716),
.C(n_707),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_785),
.B(n_776),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_785),
.B(n_776),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_678),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_785),
.B(n_776),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_897),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_853),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_990),
.B(n_992),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_995),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_SL g1004 ( 
.A1(n_945),
.A2(n_880),
.B(n_877),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_951),
.B(n_835),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_908),
.B(n_949),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_SL g1007 ( 
.A1(n_880),
.A2(n_872),
.B(n_873),
.Y(n_1007)
);

AOI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_904),
.A2(n_914),
.B(n_912),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_997),
.B(n_952),
.Y(n_1009)
);

AO31x2_ASAP7_75t_L g1010 ( 
.A1(n_977),
.A2(n_875),
.A3(n_858),
.B(n_860),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_856),
.A2(n_871),
.B(n_882),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_967),
.A2(n_926),
.B(n_917),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_907),
.A2(n_826),
.B(n_821),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_952),
.B(n_961),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_980),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_822),
.A2(n_906),
.B(n_846),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_859),
.B(n_864),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_853),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_966),
.A2(n_975),
.B(n_969),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_961),
.B(n_964),
.Y(n_1020)
);

O2A1O1Ixp5_ASAP7_75t_L g1021 ( 
.A1(n_911),
.A2(n_970),
.B(n_887),
.C(n_874),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_982),
.A2(n_989),
.B(n_985),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_946),
.A2(n_981),
.B(n_955),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_946),
.A2(n_981),
.B(n_993),
.C(n_977),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_883),
.A2(n_886),
.B(n_854),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_958),
.A2(n_976),
.B(n_884),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_964),
.B(n_974),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_974),
.B(n_979),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_SL g1029 ( 
.A1(n_872),
.A2(n_873),
.B(n_922),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_828),
.A2(n_825),
.B(n_936),
.Y(n_1030)
);

BUFx2_ASAP7_75t_SL g1031 ( 
.A(n_996),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_836),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_867),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_979),
.B(n_983),
.Y(n_1034)
);

OAI21xp33_ASAP7_75t_SL g1035 ( 
.A1(n_991),
.A2(n_983),
.B(n_987),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_L g1036 ( 
.A1(n_889),
.A2(n_938),
.B(n_924),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_825),
.A2(n_891),
.B(n_838),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_954),
.B(n_835),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_894),
.A2(n_895),
.B(n_987),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_838),
.A2(n_861),
.B(n_899),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_862),
.A2(n_839),
.B(n_913),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_988),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_839),
.A2(n_913),
.B(n_942),
.Y(n_1043)
);

OAI22x1_ASAP7_75t_L g1044 ( 
.A1(n_921),
.A2(n_896),
.B1(n_940),
.B2(n_925),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_918),
.A2(n_852),
.B(n_915),
.C(n_910),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_988),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_986),
.A2(n_864),
.B1(n_859),
.B2(n_841),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_950),
.A2(n_968),
.B(n_965),
.C(n_847),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_834),
.A2(n_840),
.B(n_876),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_986),
.A2(n_841),
.B(n_827),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_905),
.B(n_932),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_859),
.B(n_864),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_SL g1053 ( 
.A1(n_943),
.A2(n_878),
.B1(n_963),
.B2(n_944),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_829),
.A2(n_919),
.B(n_832),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_927),
.B(n_931),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_928),
.A2(n_920),
.B(n_850),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_930),
.B(n_923),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_853),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_832),
.A2(n_934),
.B(n_866),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_889),
.B(n_916),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_898),
.B(n_890),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_939),
.B(n_943),
.C(n_879),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_831),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_845),
.A2(n_849),
.B(n_842),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_956),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_890),
.B(n_844),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_903),
.B(n_851),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_844),
.B(n_900),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_900),
.A2(n_833),
.B(n_830),
.C(n_978),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_901),
.B(n_881),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_866),
.A2(n_869),
.B(n_929),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_881),
.B(n_971),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_857),
.A2(n_885),
.B(n_937),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_865),
.B(n_824),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_881),
.A2(n_902),
.B(n_984),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_902),
.A2(n_973),
.B(n_972),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_948),
.B(n_971),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_868),
.B(n_892),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_843),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_948),
.A2(n_971),
.B(n_953),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_948),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_888),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_868),
.A2(n_892),
.A3(n_893),
.B(n_941),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_941),
.A2(n_933),
.B(n_973),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_973),
.A2(n_888),
.B(n_870),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_888),
.A2(n_870),
.B(n_935),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_870),
.A2(n_848),
.B(n_947),
.Y(n_1087)
);

OA22x2_ASAP7_75t_L g1088 ( 
.A1(n_962),
.A2(n_943),
.B1(n_908),
.B2(n_873),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_855),
.A2(n_959),
.B(n_957),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_859),
.B(n_864),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_909),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_831),
.Y(n_1094)
);

AO22x2_ASAP7_75t_L g1095 ( 
.A1(n_873),
.A2(n_977),
.B1(n_921),
.B2(n_943),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_908),
.A2(n_904),
.B(n_914),
.C(n_912),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_954),
.B(n_722),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_908),
.A2(n_904),
.B1(n_914),
.B2(n_912),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_990),
.B(n_992),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_L g1103 ( 
.A(n_859),
.B(n_864),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_990),
.B(n_992),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_908),
.A2(n_904),
.B(n_914),
.C(n_912),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_908),
.A2(n_904),
.B1(n_914),
.B2(n_912),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1109)
);

AOI22x1_ASAP7_75t_L g1110 ( 
.A1(n_894),
.A2(n_882),
.B1(n_913),
.B2(n_899),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_977),
.A2(n_875),
.A3(n_858),
.B(n_860),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_883),
.A2(n_886),
.B(n_958),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_883),
.A2(n_886),
.B(n_958),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_873),
.A2(n_955),
.B1(n_991),
.B2(n_904),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_980),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_867),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_980),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_990),
.B(n_992),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_980),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_897),
.Y(n_1124)
);

NAND2x1_ASAP7_75t_L g1125 ( 
.A(n_866),
.B(n_786),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_897),
.Y(n_1126)
);

OAI22x1_ASAP7_75t_L g1127 ( 
.A1(n_908),
.A2(n_789),
.B1(n_924),
.B2(n_736),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_954),
.B(n_722),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_837),
.A2(n_863),
.B(n_823),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_990),
.B(n_992),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_990),
.B(n_992),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_908),
.B(n_949),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_908),
.B(n_949),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_883),
.A2(n_886),
.B(n_958),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_856),
.A2(n_871),
.B(n_882),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_954),
.B(n_722),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_990),
.B(n_992),
.Y(n_1140)
);

OAI21xp33_ASAP7_75t_SL g1141 ( 
.A1(n_955),
.A2(n_713),
.B(n_991),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_912),
.A2(n_914),
.B(n_904),
.C(n_911),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_960),
.B(n_959),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_977),
.A2(n_875),
.A3(n_858),
.B(n_860),
.Y(n_1144)
);

OAI21xp33_ASAP7_75t_SL g1145 ( 
.A1(n_955),
.A2(n_713),
.B(n_991),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_908),
.A2(n_946),
.B(n_981),
.C(n_993),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1039),
.A2(n_1114),
.B(n_1112),
.Y(n_1147)
);

NAND2x1p5_ASAP7_75t_L g1148 ( 
.A(n_1078),
.B(n_999),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1123),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_1118),
.B(n_1119),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1127),
.A2(n_1133),
.B1(n_1006),
.B2(n_1134),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1135),
.A2(n_1029),
.B(n_1026),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1005),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_1036),
.A2(n_1054),
.B(n_1064),
.C(n_1089),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1088),
.A2(n_1133),
.B1(n_1006),
.B2(n_1134),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1098),
.B(n_1129),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1001),
.A2(n_1097),
.B(n_1090),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1039),
.A2(n_1056),
.B(n_1096),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1146),
.A2(n_1024),
.B(n_1045),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_998),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1161)
);

INVx3_ASAP7_75t_SL g1162 ( 
.A(n_1079),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1056),
.A2(n_1106),
.B(n_1100),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1110),
.A2(n_1019),
.B(n_1002),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1107),
.B(n_1146),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_SL g1166 ( 
.A1(n_1053),
.A2(n_1088),
.B1(n_1060),
.B2(n_1095),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1027),
.B(n_1028),
.Y(n_1167)
);

CKINVDCx11_ASAP7_75t_R g1168 ( 
.A(n_1117),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1034),
.A2(n_1009),
.B1(n_1000),
.B2(n_1140),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1015),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1032),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1057),
.B(n_1003),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1042),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1031),
.B(n_1075),
.Y(n_1175)
);

AOI222xp33_ASAP7_75t_L g1176 ( 
.A1(n_1044),
.A2(n_1104),
.B1(n_1132),
.B2(n_1121),
.C1(n_1102),
.C2(n_1131),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1060),
.A2(n_1137),
.B1(n_1062),
.B2(n_1033),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1124),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1078),
.B(n_1081),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1008),
.B(n_1115),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1038),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1051),
.B(n_1055),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1115),
.B(n_1035),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1061),
.A2(n_1047),
.B1(n_1067),
.B2(n_1095),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_1082),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1082),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_1023),
.A2(n_1050),
.B(n_1071),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1126),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_1046),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1070),
.B(n_1066),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1068),
.B(n_1093),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1018),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1019),
.A2(n_1022),
.B(n_1113),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1095),
.B(n_1077),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1082),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1075),
.B(n_1092),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_1018),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1022),
.A2(n_1113),
.B(n_1143),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1018),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1018),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1072),
.B(n_1010),
.Y(n_1201)
);

AND2x2_ASAP7_75t_SL g1202 ( 
.A(n_1103),
.B(n_1058),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1084),
.B(n_1076),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1074),
.A2(n_1052),
.B1(n_1017),
.B2(n_1145),
.Y(n_1204)
);

BUFx2_ASAP7_75t_SL g1205 ( 
.A(n_1058),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1023),
.B(n_1024),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1092),
.B(n_1089),
.Y(n_1207)
);

BUFx2_ASAP7_75t_SL g1208 ( 
.A(n_1058),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1091),
.A2(n_1138),
.B(n_1128),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1058),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1141),
.B(n_1144),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1086),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1085),
.B(n_1080),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1142),
.B(n_1144),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1073),
.A2(n_1069),
.B1(n_1007),
.B2(n_1059),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1063),
.B(n_1065),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1142),
.B(n_1010),
.Y(n_1217)
);

INVxp67_ASAP7_75t_SL g1218 ( 
.A(n_1063),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1083),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1091),
.A2(n_1139),
.B(n_1138),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1083),
.Y(n_1222)
);

INVx3_ASAP7_75t_SL g1223 ( 
.A(n_1065),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1087),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1010),
.B(n_1111),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1099),
.A2(n_1109),
.B(n_1108),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1059),
.A2(n_1094),
.B1(n_1071),
.B2(n_1144),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1010),
.B(n_1111),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1111),
.B(n_1144),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1004),
.B(n_1021),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1111),
.B(n_1021),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1043),
.B(n_1030),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_SL g1233 ( 
.A(n_1048),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1105),
.A2(n_1122),
.B(n_1139),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1105),
.A2(n_1122),
.B(n_1012),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1049),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_SL g1237 ( 
.A1(n_1048),
.A2(n_1025),
.B(n_1136),
.C(n_1011),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1037),
.A2(n_1013),
.B(n_1040),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1041),
.B(n_1101),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_R g1240 ( 
.A(n_1125),
.B(n_1116),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1016),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1120),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1130),
.B(n_1098),
.Y(n_1243)
);

BUFx2_ASAP7_75t_SL g1244 ( 
.A(n_1123),
.Y(n_1244)
);

NOR3xp33_ASAP7_75t_L g1245 ( 
.A(n_1036),
.B(n_924),
.C(n_970),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1014),
.A2(n_1027),
.B1(n_1028),
.B2(n_1020),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1098),
.B(n_1129),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1005),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1039),
.A2(n_713),
.B(n_700),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1112),
.A2(n_1135),
.B(n_1114),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1060),
.B(n_347),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1098),
.B(n_1129),
.Y(n_1255)
);

INVx3_ASAP7_75t_SL g1256 ( 
.A(n_1118),
.Y(n_1256)
);

OR2x6_ASAP7_75t_SL g1257 ( 
.A(n_1118),
.B(n_810),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1098),
.B(n_1129),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1078),
.B(n_868),
.Y(n_1259)
);

INVx5_ASAP7_75t_L g1260 ( 
.A(n_1082),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1039),
.A2(n_1114),
.B(n_1112),
.Y(n_1261)
);

INVx3_ASAP7_75t_SL g1262 ( 
.A(n_1118),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1005),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1078),
.B(n_868),
.Y(n_1268)
);

INVx2_ASAP7_75t_SL g1269 ( 
.A(n_1123),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1098),
.B(n_1129),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1031),
.B(n_1075),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_999),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1005),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1082),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1078),
.B(n_999),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1031),
.B(n_1075),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1079),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1015),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1014),
.B(n_1020),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_1078),
.B(n_859),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1036),
.A2(n_993),
.B(n_904),
.C(n_889),
.Y(n_1285)
);

INVx3_ASAP7_75t_SL g1286 ( 
.A(n_1118),
.Y(n_1286)
);

INVx6_ASAP7_75t_L g1287 ( 
.A(n_1260),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1168),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1285),
.A2(n_1151),
.B(n_1245),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1173),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1188),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1165),
.A2(n_1155),
.B1(n_1166),
.B2(n_1176),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1260),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1256),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1260),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1161),
.A2(n_1263),
.B1(n_1283),
.B2(n_1264),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1182),
.B(n_1172),
.Y(n_1297)
);

OR2x6_ASAP7_75t_L g1298 ( 
.A(n_1207),
.B(n_1159),
.Y(n_1298)
);

AOI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1251),
.A2(n_1238),
.B(n_1235),
.Y(n_1299)
);

OA21x2_ASAP7_75t_L g1300 ( 
.A1(n_1164),
.A2(n_1235),
.B(n_1193),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1282),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_SL g1302 ( 
.A(n_1149),
.Y(n_1302)
);

CKINVDCx11_ASAP7_75t_R g1303 ( 
.A(n_1257),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1284),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1153),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1165),
.A2(n_1177),
.B1(n_1264),
.B2(n_1266),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1178),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1169),
.B(n_1161),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1254),
.A2(n_1159),
.B1(n_1169),
.B2(n_1180),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1262),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1167),
.B(n_1249),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1189),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1156),
.B(n_1247),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1157),
.A2(n_1226),
.B(n_1234),
.Y(n_1314)
);

AO21x1_ASAP7_75t_L g1315 ( 
.A1(n_1246),
.A2(n_1183),
.B(n_1163),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1167),
.B(n_1249),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1171),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1281),
.Y(n_1318)
);

CKINVDCx6p67_ASAP7_75t_R g1319 ( 
.A(n_1286),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1152),
.A2(n_1253),
.B1(n_1183),
.B2(n_1246),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1230),
.A2(n_1215),
.B1(n_1283),
.B2(n_1252),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1250),
.A2(n_1252),
.B1(n_1267),
.B2(n_1279),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1153),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1250),
.A2(n_1267),
.B1(n_1263),
.B2(n_1279),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1191),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1170),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1266),
.B(n_1273),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1221),
.A2(n_1238),
.B(n_1147),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1190),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1147),
.A2(n_1261),
.B(n_1209),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1162),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1181),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1194),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1179),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1248),
.Y(n_1335)
);

BUFx2_ASAP7_75t_R g1336 ( 
.A(n_1244),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1185),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1198),
.A2(n_1158),
.B(n_1236),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1273),
.A2(n_1274),
.B1(n_1277),
.B2(n_1206),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1255),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1274),
.A2(n_1277),
.B1(n_1206),
.B2(n_1187),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1248),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1192),
.Y(n_1343)
);

INVx4_ASAP7_75t_SL g1344 ( 
.A(n_1284),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1265),
.A2(n_1275),
.B1(n_1229),
.B2(n_1225),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1184),
.A2(n_1204),
.B1(n_1265),
.B2(n_1275),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1201),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1197),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1269),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1210),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1224),
.A2(n_1280),
.B1(n_1271),
.B2(n_1175),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1230),
.A2(n_1215),
.B1(n_1258),
.B2(n_1270),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1243),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1228),
.A2(n_1261),
.B1(n_1211),
.B2(n_1231),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1218),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1223),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1211),
.A2(n_1232),
.B(n_1214),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1203),
.A2(n_1217),
.B1(n_1280),
.B2(n_1271),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1232),
.A2(n_1227),
.B(n_1239),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1185),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1242),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1233),
.A2(n_1202),
.B1(n_1280),
.B2(n_1175),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1268),
.B(n_1203),
.Y(n_1363)
);

BUFx2_ASAP7_75t_R g1364 ( 
.A(n_1205),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1199),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1213),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1175),
.A2(n_1271),
.B1(n_1207),
.B2(n_1196),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1216),
.B(n_1219),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1208),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1213),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1195),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1200),
.Y(n_1372)
);

BUFx2_ASAP7_75t_R g1373 ( 
.A(n_1212),
.Y(n_1373)
);

NAND2x1p5_ASAP7_75t_L g1374 ( 
.A(n_1174),
.B(n_1150),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1272),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1272),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1241),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1196),
.A2(n_1207),
.B1(n_1148),
.B2(n_1278),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1196),
.A2(n_1222),
.B1(n_1220),
.B2(n_1284),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1186),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1148),
.B(n_1278),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1186),
.Y(n_1382)
);

AOI222xp33_ASAP7_75t_L g1383 ( 
.A1(n_1154),
.A2(n_1237),
.B1(n_1174),
.B2(n_1186),
.C1(n_1276),
.C2(n_1241),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1240),
.A2(n_1241),
.B(n_1276),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1276),
.A2(n_889),
.B1(n_904),
.B2(n_756),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1153),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1196),
.B(n_1259),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_889),
.B1(n_924),
.B2(n_963),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1260),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1282),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_SL g1391 ( 
.A(n_1149),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1182),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1161),
.A2(n_908),
.B1(n_1249),
.B2(n_1167),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1157),
.A2(n_1226),
.B(n_1235),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1156),
.B(n_1247),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1160),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1260),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1254),
.A2(n_889),
.B1(n_924),
.B2(n_963),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1165),
.A2(n_889),
.B1(n_1053),
.B2(n_1088),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1333),
.B(n_1347),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1313),
.Y(n_1401)
);

BUFx2_ASAP7_75t_SL g1402 ( 
.A(n_1356),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1353),
.B(n_1354),
.Y(n_1403)
);

BUFx2_ASAP7_75t_SL g1404 ( 
.A(n_1356),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1335),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1342),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1388),
.A2(n_1398),
.B(n_1309),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1298),
.B(n_1289),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1394),
.A2(n_1314),
.B(n_1299),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1357),
.B(n_1320),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1297),
.A2(n_1298),
.B1(n_1311),
.B2(n_1316),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1298),
.B(n_1368),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1290),
.Y(n_1413)
);

INVx3_ASAP7_75t_L g1414 ( 
.A(n_1384),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1357),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1315),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1394),
.A2(n_1314),
.B(n_1338),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1305),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1312),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1384),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1327),
.B(n_1322),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1385),
.A2(n_1392),
.B1(n_1346),
.B2(n_1362),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_1340),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1359),
.A2(n_1320),
.B(n_1341),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1350),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1350),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1350),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1287),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1308),
.A2(n_1378),
.B(n_1300),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1322),
.B(n_1324),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1328),
.A2(n_1330),
.B(n_1351),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1330),
.A2(n_1306),
.B(n_1361),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1345),
.B(n_1341),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1345),
.B(n_1358),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1392),
.B(n_1317),
.Y(n_1436)
);

CKINVDCx8_ASAP7_75t_R g1437 ( 
.A(n_1344),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1344),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1307),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1323),
.Y(n_1440)
);

BUFx2_ASAP7_75t_SL g1441 ( 
.A(n_1392),
.Y(n_1441)
);

AO21x2_ASAP7_75t_L g1442 ( 
.A1(n_1361),
.A2(n_1377),
.B(n_1393),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_SL g1443 ( 
.A(n_1304),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1321),
.B(n_1358),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1339),
.B(n_1329),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1291),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1339),
.B(n_1352),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1386),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1396),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1387),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1301),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1367),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1363),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1363),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1390),
.B(n_1334),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1325),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1355),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1387),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1296),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1383),
.Y(n_1460)
);

INVx2_ASAP7_75t_SL g1461 ( 
.A(n_1287),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1381),
.B(n_1379),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1292),
.A2(n_1379),
.B(n_1324),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1415),
.Y(n_1464)
);

INVx4_ASAP7_75t_L g1465 ( 
.A(n_1443),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1410),
.B(n_1332),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1292),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1407),
.A2(n_1399),
.B1(n_1431),
.B2(n_1411),
.C(n_1447),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1459),
.B(n_1348),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1424),
.B(n_1343),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1415),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1426),
.B(n_1381),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1403),
.B(n_1375),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1403),
.B(n_1372),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1410),
.B(n_1376),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1447),
.A2(n_1303),
.B1(n_1288),
.B2(n_1334),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1421),
.B(n_1373),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1420),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1422),
.B(n_1344),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1420),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1432),
.B(n_1380),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1409),
.A2(n_1374),
.B(n_1382),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1406),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1408),
.B(n_1365),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1408),
.B(n_1371),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1452),
.B(n_1371),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1452),
.B(n_1389),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1442),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1414),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1414),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1445),
.B(n_1369),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1441),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1460),
.C(n_1416),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1466),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1405),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1483),
.B(n_1491),
.Y(n_1497)
);

AND4x1_ASAP7_75t_L g1498 ( 
.A(n_1468),
.B(n_1436),
.C(n_1460),
.D(n_1444),
.Y(n_1498)
);

OAI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1476),
.A2(n_1451),
.B1(n_1419),
.B2(n_1441),
.C(n_1401),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1477),
.B(n_1450),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1491),
.B(n_1413),
.Y(n_1501)
);

OAI221xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1476),
.A2(n_1444),
.B1(n_1477),
.B2(n_1434),
.C(n_1467),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1478),
.B(n_1414),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1484),
.B(n_1412),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1479),
.A2(n_1443),
.B(n_1438),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1484),
.B(n_1432),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1479),
.A2(n_1463),
.B1(n_1435),
.B2(n_1462),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1469),
.B(n_1416),
.C(n_1463),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1485),
.B(n_1462),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1402),
.Y(n_1510)
);

NAND4xp25_ASAP7_75t_L g1511 ( 
.A(n_1469),
.B(n_1423),
.C(n_1445),
.D(n_1456),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1485),
.B(n_1462),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1481),
.B(n_1463),
.C(n_1418),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1493),
.A2(n_1374),
.B1(n_1455),
.B2(n_1404),
.C(n_1402),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1485),
.B(n_1462),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_L g1517 ( 
.A1(n_1467),
.A2(n_1434),
.B(n_1435),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1470),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1486),
.B(n_1440),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1464),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1467),
.A2(n_1463),
.B1(n_1404),
.B2(n_1438),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1492),
.A2(n_1409),
.B(n_1417),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1482),
.A2(n_1453),
.B(n_1454),
.Y(n_1525)
);

OAI211xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1481),
.A2(n_1303),
.B(n_1456),
.C(n_1439),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1481),
.B(n_1446),
.C(n_1449),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1473),
.B(n_1400),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1473),
.B(n_1400),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1474),
.B(n_1458),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1466),
.A2(n_1437),
.B1(n_1336),
.B2(n_1364),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1465),
.B(n_1450),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1475),
.B(n_1458),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1474),
.B(n_1487),
.Y(n_1534)
);

NOR3xp33_ASAP7_75t_L g1535 ( 
.A(n_1465),
.B(n_1438),
.C(n_1429),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1474),
.B(n_1458),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1433),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1492),
.B(n_1446),
.C(n_1449),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1465),
.B(n_1438),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1521),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1521),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1519),
.B(n_1480),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1495),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1537),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1527),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1506),
.B(n_1480),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1503),
.B(n_1490),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1506),
.B(n_1480),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1524),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1503),
.B(n_1490),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1524),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1524),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1527),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1538),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1503),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1538),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1503),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_SL g1561 ( 
.A(n_1539),
.B(n_1465),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1513),
.B(n_1466),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1533),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1525),
.B(n_1490),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1517),
.B(n_1497),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1515),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1518),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1532),
.B(n_1490),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1534),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1504),
.B(n_1490),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1530),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1517),
.B(n_1464),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1520),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1556),
.B(n_1508),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1540),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1556),
.A2(n_1494),
.B1(n_1502),
.B2(n_1513),
.C(n_1508),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1566),
.B(n_1572),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1543),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1542),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1543),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1569),
.B(n_1535),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1572),
.B(n_1501),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1541),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1571),
.B(n_1510),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1556),
.B(n_1496),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1561),
.A2(n_1494),
.B1(n_1498),
.B2(n_1531),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1523),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1564),
.B(n_1505),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1572),
.B(n_1522),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1569),
.B(n_1490),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1541),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.B(n_1536),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1557),
.B(n_1294),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1563),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1528),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1563),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1529),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1472),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1571),
.B(n_1472),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1542),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1559),
.B(n_1545),
.Y(n_1605)
);

OAI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1559),
.A2(n_1507),
.B(n_1511),
.C(n_1499),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1545),
.B(n_1471),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1545),
.B(n_1554),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1487),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_L g1610 ( 
.A(n_1554),
.B(n_1505),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1487),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1563),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1576),
.Y(n_1614)
);

OR2x6_ASAP7_75t_SL g1615 ( 
.A(n_1575),
.B(n_1562),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1577),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1580),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1608),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1557),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1578),
.A2(n_1554),
.B(n_1562),
.C(n_1573),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1606),
.B(n_1570),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1498),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1582),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1573),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1581),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1583),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1587),
.B(n_1590),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1589),
.A2(n_1561),
.B1(n_1514),
.B2(n_1562),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1590),
.A2(n_1526),
.B1(n_1569),
.B2(n_1564),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1608),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1579),
.B(n_1568),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1582),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1610),
.B(n_1569),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1612),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1612),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1591),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1605),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1602),
.B(n_1557),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1585),
.B(n_1555),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1465),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1584),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1593),
.B(n_1555),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1596),
.B(n_1555),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1596),
.B(n_1586),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1598),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1602),
.B(n_1553),
.Y(n_1652)
);

INVxp67_ASAP7_75t_L g1653 ( 
.A(n_1575),
.Y(n_1653)
);

AND2x2_ASAP7_75t_SL g1654 ( 
.A(n_1584),
.B(n_1465),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1600),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1629),
.B(n_1584),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1654),
.B(n_1592),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1631),
.A2(n_1592),
.B1(n_1564),
.B2(n_1569),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1631),
.A2(n_1595),
.B1(n_1500),
.B2(n_1599),
.C(n_1601),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1654),
.B(n_1603),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1661)
);

AND3x1_ASAP7_75t_L g1662 ( 
.A(n_1624),
.B(n_1632),
.C(n_1622),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1624),
.A2(n_1564),
.B1(n_1604),
.B2(n_1488),
.Y(n_1663)
);

OR2x6_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_1288),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1642),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1646),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1614),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1637),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1647),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1653),
.A2(n_1564),
.B(n_1607),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1615),
.B(n_1310),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1615),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1613),
.B(n_1609),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1647),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1627),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1551),
.B(n_1549),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1626),
.B(n_1611),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1650),
.B(n_1544),
.Y(n_1681)
);

AND2x4_ASAP7_75t_SL g1682 ( 
.A(n_1634),
.B(n_1645),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1603),
.Y(n_1683)
);

AO22x1_ASAP7_75t_L g1684 ( 
.A1(n_1620),
.A2(n_1594),
.B1(n_1569),
.B2(n_1564),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1634),
.Y(n_1685)
);

OAI22x1_ASAP7_75t_L g1686 ( 
.A1(n_1620),
.A2(n_1594),
.B1(n_1558),
.B2(n_1560),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1630),
.B(n_1628),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1634),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1651),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1645),
.B(n_1594),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1655),
.B(n_1310),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1674),
.B(n_1621),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1662),
.A2(n_1633),
.B1(n_1635),
.B2(n_1639),
.C(n_1625),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1673),
.A2(n_1633),
.B1(n_1641),
.B2(n_1639),
.C(n_1636),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1691),
.B(n_1294),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1672),
.Y(n_1696)
);

OAI321xp33_ASAP7_75t_L g1697 ( 
.A1(n_1659),
.A2(n_1641),
.A3(n_1636),
.B1(n_1649),
.B2(n_1618),
.C(n_1619),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1661),
.B(n_1644),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1677),
.B(n_1643),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1656),
.B(n_1652),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1656),
.B(n_1648),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_1560),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1546),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1667),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1658),
.A2(n_1560),
.B1(n_1558),
.B2(n_1544),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1546),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1689),
.Y(n_1708)
);

OAI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1673),
.A2(n_1617),
.B1(n_1616),
.B2(n_1607),
.C(n_1558),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1678),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1665),
.B(n_1546),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1685),
.A2(n_1550),
.B1(n_1547),
.B2(n_1560),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1666),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1669),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1657),
.A2(n_1550),
.B(n_1547),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1669),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1688),
.B(n_1548),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1714),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1716),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1692),
.B(n_1687),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1701),
.B(n_1660),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1697),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1702),
.B(n_1668),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1701),
.B(n_1682),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1713),
.B(n_1668),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1694),
.B(n_1668),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1703),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1695),
.Y(n_1729)
);

NAND2x1p5_ASAP7_75t_L g1730 ( 
.A(n_1705),
.B(n_1657),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1700),
.B(n_1675),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.Y(n_1732)
);

AND3x1_ASAP7_75t_L g1733 ( 
.A(n_1693),
.B(n_1710),
.C(n_1708),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1709),
.A2(n_1664),
.B(n_1682),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1696),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1698),
.B(n_1699),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1704),
.B(n_1683),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1723),
.A2(n_1664),
.B1(n_1715),
.B2(n_1706),
.C(n_1663),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1723),
.A2(n_1664),
.B1(n_1690),
.B2(n_1717),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1729),
.A2(n_1707),
.B(n_1711),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1721),
.B(n_1683),
.Y(n_1741)
);

OAI21xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1727),
.A2(n_1663),
.B(n_1712),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1734),
.A2(n_1671),
.B(n_1690),
.C(n_1681),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1730),
.A2(n_1427),
.B(n_1425),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1725),
.B(n_1686),
.Y(n_1745)
);

OAI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1726),
.A2(n_1680),
.B(n_1664),
.C(n_1427),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1725),
.A2(n_1428),
.B(n_1326),
.C(n_1331),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_L g1748 ( 
.A1(n_1736),
.A2(n_1724),
.B(n_1728),
.C(n_1732),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1730),
.A2(n_1331),
.B(n_1428),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1733),
.A2(n_1686),
.B1(n_1684),
.B2(n_1679),
.C(n_1549),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_L g1751 ( 
.A(n_1748),
.B(n_1718),
.Y(n_1751)
);

OA22x2_ASAP7_75t_L g1752 ( 
.A1(n_1744),
.A2(n_1728),
.B1(n_1732),
.B2(n_1721),
.Y(n_1752)
);

NAND4xp25_ASAP7_75t_L g1753 ( 
.A(n_1739),
.B(n_1720),
.C(n_1722),
.D(n_1731),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1745),
.B(n_1719),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1741),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1749),
.B(n_1735),
.C(n_1737),
.Y(n_1756)
);

AOI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1742),
.A2(n_1326),
.B(n_1319),
.C(n_1349),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1750),
.A2(n_1565),
.B(n_1552),
.C(n_1549),
.Y(n_1758)
);

NOR2xp67_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1318),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1747),
.B(n_1318),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1740),
.B(n_1319),
.Y(n_1761)
);

NOR3x1_ASAP7_75t_L g1762 ( 
.A(n_1753),
.B(n_1738),
.C(n_1743),
.Y(n_1762)
);

NOR4xp25_ASAP7_75t_L g1763 ( 
.A(n_1755),
.B(n_1679),
.C(n_1551),
.D(n_1549),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1754),
.B(n_1548),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1751),
.B(n_1548),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1544),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1759),
.B(n_1349),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1767),
.B(n_1752),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1764),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1765),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1766),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1762),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1763),
.B(n_1757),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1764),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1768),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1768),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1769),
.Y(n_1777)
);

NOR2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1772),
.B(n_1761),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1770),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1777),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1777),
.B(n_1778),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1779),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1780),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1775),
.B1(n_1772),
.B2(n_1776),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1781),
.B1(n_1780),
.B2(n_1774),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1784),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1786),
.A2(n_1781),
.B(n_1782),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1785),
.B(n_1781),
.C(n_1782),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1771),
.B1(n_1782),
.B2(n_1773),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1787),
.A2(n_1760),
.B1(n_1758),
.B2(n_1391),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1789),
.A2(n_1302),
.B1(n_1558),
.B2(n_1565),
.Y(n_1791)
);

OAI221xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1791),
.A2(n_1790),
.B1(n_1337),
.B2(n_1360),
.C(n_1295),
.Y(n_1792)
);

AOI221xp5_ASAP7_75t_L g1793 ( 
.A1(n_1792),
.A2(n_1337),
.B1(n_1360),
.B2(n_1551),
.C(n_1565),
.Y(n_1793)
);

AOI211xp5_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1293),
.B(n_1397),
.C(n_1461),
.Y(n_1794)
);


endmodule