module real_jpeg_8790_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_328, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_328;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_10),
.B1(n_38),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_2),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_105),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_105),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_5),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_5),
.B(n_21),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_5),
.A2(n_9),
.B(n_27),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_42),
.B(n_55),
.C(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_42),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_6),
.A2(n_9),
.B(n_42),
.C(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_10),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_48),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_21),
.B1(n_22),
.B2(n_48),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_9),
.A2(n_38),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_9),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_54),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_11),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_39),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_11),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_81),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_79),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_73),
.Y(n_14)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.C(n_66),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_16),
.A2(n_17),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_51),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_18),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_18),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_18),
.A2(n_107),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_18),
.A2(n_51),
.B1(n_52),
.B2(n_107),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_19),
.A2(n_98),
.B(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_20),
.B(n_171),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_20),
.B(n_99),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_21),
.A2(n_34),
.B(n_56),
.Y(n_202)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_22),
.A2(n_29),
.B(n_34),
.C(n_167),
.Y(n_166)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_26),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_26),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_26),
.B(n_33),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_27),
.B(n_92),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_30),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_31),
.B(n_34),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_31),
.A2(n_207),
.B(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_34),
.B(n_92),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_35),
.A2(n_36),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_45),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_40),
.B(n_41),
.C(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_40),
.A2(n_49),
.B(n_77),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_42),
.B(n_44),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_43),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_46),
.B(n_103),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_49),
.B(n_77),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_50),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_55),
.B(n_63),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_55),
.A2(n_58),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_57),
.B(n_59),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_59),
.A2(n_145),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_60),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_64),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_64),
.A2(n_66),
.B1(n_250),
.B2(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_66),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_70),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_75),
.B(n_116),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_78),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_319),
.B(n_325),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_295),
.A3(n_314),
.B1(n_317),
.B2(n_318),
.C(n_328),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_273),
.B(n_294),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_254),
.B(n_272),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_153),
.B(n_236),
.C(n_253),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_136),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_87),
.B(n_136),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_112),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_101),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_89),
.B(n_101),
.C(n_112),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_90),
.B(n_97),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B(n_95),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_91),
.A2(n_92),
.B(n_151),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_94),
.B(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_93),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_93),
.B(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_176),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_98),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_106),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_107),
.B(n_299),
.C(n_304),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_110),
.B(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_123),
.B1(n_124),
.B2(n_135),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_122),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_114),
.B(n_122),
.C(n_123),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_127),
.B(n_193),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_142),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_137),
.A2(n_138),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_144),
.B(n_219),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_145),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_235),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_229),
.B(n_234),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_214),
.B(n_228),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_195),
.B(n_213),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_183),
.B(n_194),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_172),
.B(n_182),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_164),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_168),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_177),
.B(n_181),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_185),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_204),
.B1(n_205),
.B2(n_212),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_199),
.A2(n_200),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_199),
.A2(n_200),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_199),
.A2(n_287),
.B(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_200),
.B(n_269),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_201),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_224),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_223),
.C(n_227),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_232),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_237),
.B(n_238),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_251),
.B2(n_252),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_245),
.C(n_252),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_243),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_267),
.B2(n_268),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_268),
.C(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_264),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_275),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_292),
.B2(n_293),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_283),
.B1(n_290),
.B2(n_291),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_291),
.C(n_293),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B(n_282),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_297),
.C(n_306),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_282),
.B(n_297),
.CI(n_306),
.CON(n_316),
.SN(n_316)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_288),
.B2(n_289),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_284),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_285),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_307),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_307),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_299),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_309),
.C(n_313),
.Y(n_320)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_315),
.B(n_316),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_316),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_322),
.Y(n_324)
);


endmodule