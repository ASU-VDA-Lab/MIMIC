module real_jpeg_11663_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_3),
.A2(n_43),
.B1(n_49),
.B2(n_53),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_43),
.B1(n_68),
.B2(n_69),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_5),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_49),
.B1(n_53),
.B2(n_90),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_90),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_90),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_29),
.B(n_35),
.C(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_8),
.B(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_30),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_8),
.A2(n_30),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_64),
.C(n_69),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_8),
.A2(n_40),
.B1(n_49),
.B2(n_53),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_8),
.A2(n_84),
.B1(n_85),
.B2(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_112),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_49),
.B1(n_53),
.B2(n_58),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_10),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_68),
.B1(n_69),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_11),
.A2(n_49),
.B1(n_53),
.B2(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_88),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_88),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_13),
.A2(n_49),
.B1(n_53),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_13),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_13),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_76),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_49),
.B1(n_53),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_251)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_319),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_312),
.B(n_318),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_278),
.B(n_309),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_256),
.B(n_277),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_229),
.B(n_255),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_124),
.B(n_205),
.C(n_228),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_103),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_23),
.B(n_103),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_79),
.C(n_94),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_24),
.B(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_45),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_59),
.C(n_78),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_26),
.B(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_27),
.A2(n_28),
.B1(n_42),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_27),
.A2(n_28),
.B1(n_107),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_27),
.A2(n_222),
.B(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_27),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_27),
.A2(n_28),
.B1(n_290),
.B2(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_27),
.A2(n_273),
.B(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_28),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_29),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_30),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_30),
.A2(n_33),
.B(n_40),
.Y(n_93)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_SL g142 ( 
.A(n_31),
.B(n_51),
.C(n_53),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_40),
.B(n_85),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_40),
.B(n_67),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_44),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_44),
.B(n_274),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_59),
.B1(n_60),
.B2(n_78),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_47),
.A2(n_57),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_48),
.B1(n_102),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_111),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_47),
.A2(n_224),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g53 ( 
.A(n_49),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_49),
.A2(n_52),
.B(n_140),
.C(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_49),
.B(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_71),
.B(n_74),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_61),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_61),
.A2(n_67),
.B(n_71),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_62),
.A2(n_77),
.B1(n_135),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_77),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_62),
.A2(n_77),
.B1(n_158),
.B2(n_168),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_62),
.A2(n_77),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_62),
.A2(n_215),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_68),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_77),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_74),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_80),
.B1(n_94),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_91),
.B2(n_92),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_91),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_122),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_83),
.A2(n_86),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_84),
.A2(n_85),
.B1(n_171),
.B2(n_179),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_84),
.A2(n_173),
.B(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_84),
.A2(n_85),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_98),
.Y(n_122)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_87),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_86),
.B(n_145),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_97),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_104),
.B(n_115),
.C(n_123),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_113),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_106),
.B(n_108),
.C(n_113),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_109),
.B(n_247),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_110),
.A2(n_112),
.B(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_112),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_112),
.A2(n_248),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_116),
.B(n_119),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_118),
.B(n_136),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_203),
.B(n_204),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_146),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_127),
.B(n_130),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_137),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_137),
.B1(n_138),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_143),
.B1(n_144),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_145),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_159),
.B(n_202),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_151),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_157),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_196),
.B(n_201),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_185),
.B(n_195),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_174),
.B(n_184),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_169),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_166),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_183),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_191),
.C(n_194),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_200),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_227),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_227),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.C(n_217),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_216),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_220),
.C(n_226),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_226),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_254),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_240),
.B1(n_252),
.B2(n_253),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_253),
.C(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_235),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_237),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_235),
.A2(n_268),
.B(n_270),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_245),
.C(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_250),
.B(n_291),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_276),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_276),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_275),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_261),
.C(n_267),
.Y(n_307)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_267),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_265),
.B(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_281),
.C(n_293),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_266),
.B(n_281),
.CI(n_293),
.CON(n_308),
.SN(n_308)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_306),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_294),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_294),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_288),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_301),
.C(n_303),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_289),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_292),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_295),
.C(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_308),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_308),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_321),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.CI(n_317),
.CON(n_314),
.SN(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);


endmodule