module fake_jpeg_19452_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx4_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_17),
.Y(n_20)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_6),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_13),
.B1(n_8),
.B2(n_12),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_16),
.B1(n_8),
.B2(n_19),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_20),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_22),
.B1(n_19),
.B2(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_30),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_26),
.C(n_9),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_9),
.C(n_7),
.Y(n_39)
);

AOI21x1_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_41),
.B(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_33),
.C(n_9),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_43)
);

AND2x4_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_14),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_7),
.C(n_14),
.Y(n_46)
);

NOR4xp25_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_21),
.C(n_3),
.D(n_5),
.Y(n_47)
);


endmodule