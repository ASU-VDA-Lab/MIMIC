module real_jpeg_29752_n_12 (n_279, n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_279;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_203;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_273;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_0),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_40),
.B1(n_42),
.B2(n_94),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_0),
.A2(n_9),
.B1(n_33),
.B2(n_94),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_4),
.A2(n_9),
.B1(n_27),
.B2(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_4),
.A2(n_27),
.B1(n_40),
.B2(n_42),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_6),
.A2(n_9),
.B1(n_33),
.B2(n_181),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_181),
.Y(n_274)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_77),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_9),
.B1(n_33),
.B2(n_35),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_9),
.B(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_8),
.B(n_32),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_10),
.B(n_40),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_57),
.B(n_76),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_8),
.B(n_39),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_10),
.B1(n_33),
.B2(n_41),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_9),
.A2(n_35),
.B(n_117),
.C(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_11),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_270),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_261),
.B(n_269),
.Y(n_13)
);

OAI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_230),
.A3(n_254),
.B1(n_259),
.B2(n_260),
.C(n_279),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_211),
.B(n_229),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_192),
.B(n_210),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_110),
.B(n_173),
.C(n_191),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_98),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_19),
.B(n_98),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_64),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_20),
.B(n_65),
.C(n_83),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_50),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_21)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_22),
.B(n_49),
.C(n_50),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_22),
.A2(n_48),
.B1(n_67),
.B2(n_101),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_22),
.B(n_101),
.C(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_22),
.A2(n_48),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_22),
.B(n_240),
.C(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_24),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_26),
.A2(n_30),
.B(n_35),
.C(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_28),
.B(n_32),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_28),
.A2(n_32),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_35),
.A2(n_40),
.B(n_77),
.C(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_35),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_35),
.B(n_78),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_36),
.B(n_107),
.C(n_108),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_36),
.A2(n_49),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_36),
.A2(n_217),
.B(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_36),
.B(n_217),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_38),
.B(n_39),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_38),
.A2(n_39),
.B1(n_237),
.B2(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_39),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_42),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_47),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_45),
.B(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_54),
.A2(n_105),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_54),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_54),
.B(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_54),
.B(n_132),
.C(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_63),
.B(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_56),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_60),
.Y(n_59)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_59),
.B(n_60),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_59),
.A2(n_63),
.B1(n_93),
.B2(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_82),
.B2(n_83),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.C(n_79),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_69),
.B1(n_70),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_84),
.B1(n_85),
.B2(n_101),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_68),
.Y(n_238)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_74),
.B1(n_78),
.B2(n_87),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_74),
.A2(n_78),
.B1(n_203),
.B2(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_78),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_79),
.A2(n_102),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_79),
.A2(n_102),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_79),
.A2(n_102),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_79),
.B(n_236),
.C(n_239),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_79),
.B(n_246),
.C(n_253),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_80),
.A2(n_81),
.B(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_84),
.A2(n_85),
.B1(n_139),
.B2(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_84),
.B(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_101),
.C(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_85),
.B(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B(n_89),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_95),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_106),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_102),
.B(n_184),
.C(n_186),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_106),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_107),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_172),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_167),
.B(n_171),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_135),
.B(n_166),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_123),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_114),
.B(n_123),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_122),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_132),
.C(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_134),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_134),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_179),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_161),
.B(n_165),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_146),
.B(n_160),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_141),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_142),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_143),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B(n_159),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_156),
.B(n_158),
.Y(n_150)
);

INVx5_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_174),
.B(n_175),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_189),
.B2(n_190),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_183),
.C(n_190),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_189),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_209),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_201),
.C(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_205),
.B1(n_206),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_205),
.A2(n_206),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_221),
.B(n_223),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_212),
.B(n_213),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_227),
.B2(n_228),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_220),
.C(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_232),
.C(n_242),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_232),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_227),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_244),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_239),
.A2(n_240),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_243),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_266),
.CI(n_268),
.CON(n_263),
.SN(n_263)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_265),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);


endmodule