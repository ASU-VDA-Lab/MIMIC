module fake_jpeg_6586_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_2),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_25),
.Y(n_45)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_SL g28 ( 
.A1(n_21),
.A2(n_0),
.B(n_1),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_16),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_15),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_19),
.C(n_12),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_14),
.B1(n_24),
.B2(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_23),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_14),
.B1(n_12),
.B2(n_19),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

OAI21x1_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_51),
.B(n_57),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_22),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_11),
.C(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_22),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_35),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_23),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_59),
.B(n_13),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_45),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_51),
.C(n_47),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_77),
.C(n_64),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_51),
.C(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_76),
.B(n_73),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_78),
.A2(n_57),
.B(n_66),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_65),
.B(n_87),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_69),
.B1(n_71),
.B2(n_62),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_67),
.B1(n_62),
.B2(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.C(n_43),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_58),
.B(n_39),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_43),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_58),
.B1(n_85),
.B2(n_75),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_56),
.B1(n_61),
.B2(n_39),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.C(n_59),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_96),
.B(n_10),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_9),
.B(n_10),
.C(n_4),
.D(n_7),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_2),
.B1(n_3),
.B2(n_48),
.C(n_46),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_101),
.C(n_3),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_3),
.B(n_48),
.Y(n_104)
);


endmodule