module fake_netlist_6_1428_n_2090 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2090);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2090;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g207 ( 
.A(n_55),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_89),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_60),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_71),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_74),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_129),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_140),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_79),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_36),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_43),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_142),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_86),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_76),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_62),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_116),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_119),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_126),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_88),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_73),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_124),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_80),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_118),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_71),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_17),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_174),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_69),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_77),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_95),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_97),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_106),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_196),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_82),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_12),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_23),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_91),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_11),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_103),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_123),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_68),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_46),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_146),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_26),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_206),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_14),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_117),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_139),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_110),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_168),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_178),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_39),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_145),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_164),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_94),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_44),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_131),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_17),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_74),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_22),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_62),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_104),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_202),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_84),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_166),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_150),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_182),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_40),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_120),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_96),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_205),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_115),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_20),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_32),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_93),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_31),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_98),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_56),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_67),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_11),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_36),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_180),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_183),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_133),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_13),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_161),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_12),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_23),
.Y(n_338)
);

BUFx8_ASAP7_75t_SL g339 ( 
.A(n_64),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_125),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_16),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_132),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_107),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_203),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_30),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_48),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_68),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_155),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_160),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_26),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_111),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_5),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_187),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_130),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_152),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_41),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_78),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_81),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_56),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_184),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_45),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_57),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_112),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_16),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_39),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_34),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_43),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_144),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_35),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_46),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_201),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_35),
.Y(n_374)
);

BUFx5_ASAP7_75t_L g375 ( 
.A(n_29),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_108),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_65),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_37),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_189),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_200),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_27),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_34),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_137),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_113),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_22),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_122),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_92),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_172),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_85),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_55),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_52),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_75),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_52),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_13),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_66),
.Y(n_395)
);

BUFx8_ASAP7_75t_SL g396 ( 
.A(n_199),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_102),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_198),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_38),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_67),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_65),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_148),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_10),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_18),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_33),
.Y(n_405)
);

INVxp33_ASAP7_75t_R g406 ( 
.A(n_5),
.Y(n_406)
);

BUFx2_ASAP7_75t_SL g407 ( 
.A(n_177),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_0),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_128),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_149),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_44),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_73),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_53),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_90),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_101),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_75),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_375),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_380),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_225),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_218),
.B(n_1),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_335),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_339),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_262),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_297),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_267),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_218),
.B(n_2),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_208),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_259),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_263),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_313),
.B(n_2),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_208),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_218),
.B(n_3),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_235),
.B(n_3),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_269),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_270),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_367),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_208),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_271),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_283),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_235),
.B(n_4),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_208),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_208),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_235),
.B(n_4),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_345),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_345),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_345),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_345),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_209),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_408),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_266),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_314),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_316),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_295),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_343),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_286),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_316),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_389),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_232),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_266),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_288),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_292),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_359),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_302),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_210),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_340),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_304),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_308),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_359),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_310),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_317),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_207),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_224),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_257),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_261),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_265),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_268),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_319),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_287),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_293),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_210),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_320),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_325),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_324),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_359),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_334),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_344),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_258),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_254),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_330),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_337),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_348),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_275),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_276),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_279),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_351),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_359),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_284),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_354),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_213),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_363),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_371),
.B(n_6),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_385),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_211),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_213),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_285),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_290),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_301),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_211),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_212),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_214),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_413),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_429),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_501),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_435),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_R g532 ( 
.A(n_461),
.B(n_214),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_436),
.A2(n_305),
.B1(n_300),
.B2(n_274),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_432),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_441),
.B(n_220),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_435),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_448),
.B(n_220),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_442),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_478),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_443),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_446),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_447),
.Y(n_545)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_426),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_465),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_474),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_475),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_238),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_473),
.B(n_238),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_437),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_L g555 ( 
.A(n_417),
.B(n_418),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_417),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_418),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_463),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_445),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_445),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_451),
.B(n_223),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_449),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_419),
.B(n_223),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_477),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_449),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_471),
.B(n_378),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_464),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_480),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_481),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_420),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_483),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_525),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_476),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_420),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_458),
.B(n_236),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_468),
.A2(n_248),
.B1(n_346),
.B2(n_222),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_453),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_425),
.B(n_280),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_421),
.B(n_215),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_454),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_467),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_491),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_495),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_506),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_431),
.A2(n_401),
.B1(n_403),
.B2(n_374),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_471),
.B(n_378),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_479),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_424),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_499),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_456),
.B(n_230),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_484),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_424),
.A2(n_430),
.B(n_428),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_428),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_440),
.B(n_229),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_430),
.Y(n_602)
);

BUFx8_ASAP7_75t_L g603 ( 
.A(n_524),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_500),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_433),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_497),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_513),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_433),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_520),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_526),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_511),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_611),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_536),
.A2(n_422),
.B1(n_515),
.B2(n_459),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_611),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_580),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_515),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_580),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_581),
.B(n_521),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_472),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_532),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_609),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_601),
.B(n_434),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_581),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_536),
.B(n_494),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_534),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_599),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_573),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_615),
.Y(n_634)
);

INVx6_ASAP7_75t_L g635 ( 
.A(n_581),
.Y(n_635)
);

INVxp67_ASAP7_75t_SL g636 ( 
.A(n_573),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_540),
.B(n_522),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_573),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_601),
.B(n_229),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_581),
.B(n_523),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_600),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_603),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_540),
.B(n_438),
.Y(n_645)
);

CKINVDCx16_ASAP7_75t_R g646 ( 
.A(n_546),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_600),
.Y(n_648)
);

AND3x1_ASAP7_75t_L g649 ( 
.A(n_579),
.B(n_455),
.C(n_472),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_530),
.B(n_524),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_610),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_568),
.B(n_280),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_608),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_561),
.B(n_291),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_561),
.B(n_291),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_597),
.B(n_240),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_534),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_608),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_589),
.B(n_407),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_528),
.B(n_502),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_608),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_534),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_539),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_601),
.A2(n_329),
.B1(n_341),
.B2(n_306),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_556),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_603),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_551),
.B(n_233),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_576),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_552),
.A2(n_273),
.B1(n_282),
.B2(n_260),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_555),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_590),
.B(n_416),
.C(n_226),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_552),
.B(n_260),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_576),
.B(n_237),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_576),
.B(n_383),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_530),
.B(n_423),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_578),
.A2(n_543),
.B1(n_545),
.B2(n_544),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_597),
.B(n_273),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_539),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_556),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_560),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_603),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_556),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_542),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_557),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_548),
.B(n_549),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_539),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_557),
.B(n_240),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_577),
.B(n_282),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_542),
.A2(n_353),
.B1(n_331),
.B2(n_327),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_546),
.B(n_427),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_568),
.B(n_462),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_577),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_560),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_577),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_SL g700 ( 
.A(n_547),
.B(n_212),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_599),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_599),
.A2(n_593),
.B1(n_595),
.B2(n_592),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_592),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_560),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_240),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_550),
.B(n_289),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_599),
.B(n_289),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_595),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_555),
.B(n_311),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_595),
.B(n_240),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_602),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_602),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_602),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_531),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_564),
.B(n_230),
.Y(n_715)
);

INVx6_ASAP7_75t_L g716 ( 
.A(n_560),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_L g717 ( 
.A(n_590),
.B(n_307),
.C(n_303),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_547),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_531),
.Y(n_719)
);

INVx4_ASAP7_75t_SL g720 ( 
.A(n_560),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_593),
.B(n_462),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_570),
.B(n_311),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_613),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_537),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_582),
.B(n_333),
.Y(n_726)
);

INVx4_ASAP7_75t_SL g727 ( 
.A(n_560),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_575),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_575),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_571),
.B(n_333),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_591),
.Y(n_733)
);

BUFx4f_ASAP7_75t_L g734 ( 
.A(n_583),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_466),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_537),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_582),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_606),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_606),
.B(n_485),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_538),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_538),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_554),
.B(n_350),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_529),
.B(n_486),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_583),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_583),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_554),
.Y(n_746)
);

BUFx10_ASAP7_75t_L g747 ( 
.A(n_574),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_559),
.Y(n_748)
);

INVx4_ASAP7_75t_SL g749 ( 
.A(n_583),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_612),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_559),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_562),
.Y(n_752)
);

AOI21x1_ASAP7_75t_L g753 ( 
.A1(n_562),
.A2(n_482),
.B(n_476),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_565),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_585),
.B(n_231),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_588),
.B(n_350),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_565),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_596),
.B(n_231),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_553),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_566),
.B(n_356),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_607),
.B(n_321),
.C(n_309),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_566),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_567),
.B(n_356),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_567),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_583),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_572),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_572),
.B(n_384),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_587),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_587),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_735),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_637),
.B(n_604),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_645),
.B(n_604),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_702),
.B(n_240),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_629),
.B(n_579),
.C(n_323),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_640),
.B(n_605),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_739),
.B(n_338),
.C(n_322),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_640),
.B(n_605),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_L g779 ( 
.A(n_680),
.B(n_234),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_640),
.B(n_583),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_687),
.B(n_598),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_639),
.A2(n_384),
.B(n_486),
.C(n_487),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_671),
.B(n_586),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_671),
.B(n_586),
.Y(n_784)
);

OAI21xp33_ASAP7_75t_L g785 ( 
.A1(n_623),
.A2(n_488),
.B(n_487),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_739),
.B(n_234),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_671),
.B(n_586),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_627),
.B(n_586),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_627),
.B(n_586),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_628),
.B(n_245),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_628),
.B(n_586),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_635),
.A2(n_243),
.B1(n_249),
.B2(n_253),
.Y(n_792)
);

O2A1O1Ixp5_ASAP7_75t_L g793 ( 
.A1(n_639),
.A2(n_272),
.B(n_397),
.C(n_387),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_701),
.B(n_245),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_701),
.A2(n_707),
.B(n_623),
.C(n_681),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_624),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_630),
.Y(n_797)
);

BUFx6f_ASAP7_75t_SL g798 ( 
.A(n_634),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_658),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_616),
.B(n_216),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_735),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_635),
.A2(n_243),
.B1(n_249),
.B2(n_253),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_635),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_743),
.B(n_255),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_670),
.A2(n_622),
.B1(n_642),
.B2(n_677),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_SL g807 ( 
.A(n_689),
.B(n_533),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_632),
.B(n_245),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_769),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_769),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_621),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_743),
.B(n_255),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_687),
.B(n_254),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_678),
.A2(n_256),
.B1(n_298),
.B2(n_299),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_732),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_761),
.B(n_256),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

NOR3x1_ASAP7_75t_L g818 ( 
.A(n_718),
.B(n_406),
.C(n_488),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_617),
.B(n_298),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_618),
.B(n_219),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_746),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_706),
.B(n_299),
.Y(n_822)
);

AOI221xp5_ASAP7_75t_L g823 ( 
.A1(n_675),
.A2(n_533),
.B1(n_251),
.B2(n_217),
.C(n_227),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_655),
.B(n_221),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_706),
.B(n_312),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_656),
.B(n_244),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_748),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_632),
.A2(n_342),
.B1(n_245),
.B2(n_359),
.Y(n_828)
);

AND2x6_ASAP7_75t_SL g829 ( 
.A(n_662),
.B(n_715),
.Y(n_829)
);

INVx8_ASAP7_75t_L g830 ( 
.A(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_673),
.B(n_246),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_624),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_757),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_636),
.B(n_247),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_624),
.Y(n_835)
);

AND2x6_ASAP7_75t_SL g836 ( 
.A(n_755),
.B(n_489),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_624),
.Y(n_837)
);

NOR2xp67_ASAP7_75t_L g838 ( 
.A(n_758),
.B(n_679),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_676),
.A2(n_489),
.B(n_527),
.C(n_518),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_737),
.B(n_264),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_762),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_714),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_696),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_764),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_696),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_632),
.A2(n_342),
.B1(n_245),
.B2(n_359),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_634),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_714),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_768),
.B(n_277),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_723),
.B(n_312),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_719),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_719),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_718),
.B(n_254),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_650),
.B(n_490),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_278),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_725),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_723),
.A2(n_360),
.B1(n_362),
.B2(n_414),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_717),
.B(n_358),
.C(n_347),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_725),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_665),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_633),
.B(n_638),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_641),
.B(n_281),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_643),
.B(n_342),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_647),
.B(n_294),
.Y(n_864)
);

O2A1O1Ixp5_ASAP7_75t_L g865 ( 
.A1(n_676),
.A2(n_379),
.B(n_355),
.C(n_357),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_736),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_654),
.B(n_342),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_659),
.B(n_342),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_730),
.B(n_360),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_736),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_660),
.B(n_664),
.Y(n_871)
);

INVxp33_ASAP7_75t_L g872 ( 
.A(n_650),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_730),
.B(n_362),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_693),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_672),
.B(n_296),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_756),
.B(n_667),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_721),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_731),
.Y(n_878)
);

OAI22xp33_ASAP7_75t_L g879 ( 
.A1(n_728),
.A2(n_242),
.B1(n_239),
.B2(n_241),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_721),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_648),
.B(n_740),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_679),
.B(n_370),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_740),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_756),
.B(n_370),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_728),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_652),
.B(n_315),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_644),
.B(n_490),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_751),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_652),
.B(n_318),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_751),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_729),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_693),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_752),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_652),
.A2(n_376),
.B1(n_414),
.B2(n_410),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_752),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_754),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_754),
.B(n_326),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_766),
.Y(n_898)
);

OAI22xp33_ASAP7_75t_L g899 ( 
.A1(n_729),
.A2(n_661),
.B1(n_620),
.B2(n_731),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_733),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_648),
.B(n_359),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_626),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_738),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_733),
.B(n_492),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_626),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_620),
.B(n_492),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_766),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_648),
.B(n_359),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_767),
.A2(n_328),
.B1(n_332),
.B2(n_336),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_666),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_666),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_682),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_668),
.B(n_349),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_683),
.B(n_352),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_686),
.B(n_365),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_648),
.B(n_398),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_620),
.B(n_376),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_763),
.A2(n_402),
.B(n_415),
.C(n_409),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_682),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_688),
.B(n_386),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_648),
.B(n_386),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_691),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_690),
.B(n_388),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_620),
.B(n_661),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_691),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_703),
.B(n_388),
.Y(n_926)
);

INVx8_ASAP7_75t_L g927 ( 
.A(n_661),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_625),
.A2(n_410),
.B1(n_217),
.B2(n_395),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_697),
.B(n_482),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_694),
.B(n_227),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_767),
.B(n_693),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_699),
.B(n_498),
.Y(n_932)
);

BUFx5_ASAP7_75t_L g933 ( 
.A(n_767),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_722),
.B(n_493),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_712),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_649),
.A2(n_594),
.B1(n_373),
.B2(n_236),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_700),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_713),
.B(n_498),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_773),
.A2(n_734),
.B(n_709),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_771),
.B(n_708),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_803),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_876),
.A2(n_726),
.B1(n_669),
.B2(n_685),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_843),
.B(n_653),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_773),
.A2(n_734),
.B(n_657),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_876),
.A2(n_822),
.B(n_850),
.C(n_825),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_794),
.A2(n_734),
.B(n_657),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_794),
.A2(n_808),
.B(n_795),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_838),
.B(n_634),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_822),
.A2(n_700),
.B(n_760),
.C(n_742),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_772),
.B(n_805),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_845),
.B(n_711),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_809),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_808),
.A2(n_765),
.B(n_745),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_937),
.A2(n_646),
.B1(n_767),
.B2(n_695),
.Y(n_954)
);

AO22x1_ASAP7_75t_L g955 ( 
.A1(n_930),
.A2(n_242),
.B1(n_228),
.B2(n_239),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_788),
.A2(n_745),
.B(n_765),
.Y(n_956)
);

NOR2x1p5_ASAP7_75t_SL g957 ( 
.A(n_933),
.B(n_753),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_789),
.A2(n_684),
.B(n_704),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_881),
.A2(n_510),
.B(n_469),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_872),
.B(n_651),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_891),
.B(n_724),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_780),
.A2(n_765),
.B(n_745),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_874),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_877),
.B(n_684),
.Y(n_964)
);

OAI321xp33_ASAP7_75t_L g965 ( 
.A1(n_930),
.A2(n_493),
.A3(n_527),
.B1(n_518),
.B2(n_517),
.C(n_516),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_783),
.A2(n_744),
.B(n_698),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_809),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_880),
.B(n_684),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_810),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_828),
.A2(n_704),
.B(n_767),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_784),
.A2(n_698),
.B(n_744),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_770),
.B(n_704),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_854),
.B(n_750),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_828),
.A2(n_767),
.B(n_693),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_787),
.A2(n_698),
.B(n_744),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_775),
.A2(n_698),
.B(n_744),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_825),
.A2(n_510),
.B(n_496),
.C(n_503),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_934),
.B(n_904),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_801),
.B(n_716),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_846),
.A2(n_693),
.B(n_692),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_810),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_777),
.A2(n_791),
.B(n_861),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_846),
.B(n_716),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_885),
.B(n_663),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_861),
.A2(n_692),
.B(n_710),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_871),
.A2(n_705),
.B(n_710),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_842),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_903),
.B(n_558),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_842),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_796),
.A2(n_727),
.B(n_749),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_786),
.B(n_569),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_878),
.Y(n_992)
);

CKINVDCx8_ASAP7_75t_R g993 ( 
.A(n_902),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_782),
.A2(n_693),
.B(n_516),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_803),
.A2(n_584),
.B1(n_716),
.B2(n_759),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_815),
.B(n_720),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_782),
.A2(n_505),
.B(n_512),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_796),
.A2(n_720),
.B(n_749),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_790),
.A2(n_826),
.B(n_824),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_790),
.A2(n_834),
.B(n_886),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_817),
.B(n_720),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_848),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_786),
.B(n_663),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_SL g1004 ( 
.A(n_823),
.B(n_759),
.C(n_394),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_821),
.B(n_720),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_906),
.Y(n_1006)
);

AOI21x1_ASAP7_75t_L g1007 ( 
.A1(n_855),
.A2(n_470),
.B(n_466),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_830),
.B(n_663),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_878),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_827),
.B(n_674),
.Y(n_1010)
);

AND2x6_ASAP7_75t_SL g1011 ( 
.A(n_781),
.B(n_496),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_889),
.A2(n_503),
.B(n_517),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_831),
.A2(n_504),
.B(n_514),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_840),
.A2(n_931),
.B(n_929),
.Y(n_1014)
);

AOI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_850),
.A2(n_391),
.B(n_241),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_833),
.B(n_674),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_926),
.A2(n_514),
.B(n_512),
.C(n_509),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_848),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_835),
.A2(n_504),
.B(n_509),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_774),
.B(n_674),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_804),
.B(n_747),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_932),
.A2(n_505),
.B(n_228),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_852),
.A2(n_377),
.B(n_412),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_852),
.A2(n_890),
.B(n_888),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_900),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_841),
.B(n_747),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_844),
.B(n_747),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_874),
.B(n_83),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_888),
.A2(n_377),
.B(n_411),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_869),
.A2(n_412),
.B1(n_411),
.B2(n_404),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_869),
.A2(n_404),
.B1(n_395),
.B2(n_394),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_793),
.A2(n_368),
.B(n_392),
.Y(n_1032)
);

NAND2x1_ASAP7_75t_L g1033 ( 
.A(n_835),
.B(n_87),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_804),
.B(n_812),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_890),
.A2(n_393),
.B(n_392),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_935),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_873),
.A2(n_393),
.B1(n_391),
.B2(n_381),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_812),
.B(n_250),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_806),
.B(n_250),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_811),
.B(n_251),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_935),
.A2(n_366),
.B(n_252),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_926),
.A2(n_236),
.B(n_373),
.C(n_381),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_920),
.A2(n_366),
.B(n_372),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_873),
.A2(n_372),
.B1(n_369),
.B2(n_368),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_923),
.A2(n_369),
.B(n_364),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_862),
.A2(n_364),
.B(n_361),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_361),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_851),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_884),
.A2(n_252),
.B1(n_373),
.B2(n_194),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_900),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_813),
.B(n_853),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_874),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_864),
.A2(n_193),
.B(n_190),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_856),
.B(n_859),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_807),
.B(n_7),
.C(n_8),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_835),
.A2(n_837),
.B(n_832),
.Y(n_1056)
);

OR2x6_ASAP7_75t_SL g1057 ( 
.A(n_905),
.B(n_8),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_866),
.B(n_9),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_835),
.A2(n_176),
.B(n_175),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_870),
.B(n_9),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_875),
.A2(n_173),
.B1(n_170),
.B2(n_169),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_819),
.A2(n_10),
.B(n_15),
.C(n_18),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_832),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_883),
.B(n_15),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_893),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_819),
.A2(n_19),
.B(n_24),
.C(n_27),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_897),
.A2(n_159),
.B(n_158),
.Y(n_1067)
);

INVx11_ASAP7_75t_L g1068 ( 
.A(n_847),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_SL g1069 ( 
.A(n_874),
.B(n_19),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_899),
.B(n_882),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_895),
.A2(n_157),
.B(n_154),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_896),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_892),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_830),
.B(n_927),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_898),
.A2(n_907),
.B(n_911),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_800),
.B(n_24),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_798),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_829),
.B(n_28),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_776),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_909),
.A2(n_147),
.B1(n_143),
.B2(n_141),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_910),
.A2(n_127),
.B(n_121),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_917),
.B(n_899),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_887),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_778),
.A2(n_799),
.B(n_797),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_820),
.B(n_33),
.Y(n_1086)
);

AND2x6_ASAP7_75t_L g1087 ( 
.A(n_892),
.B(n_100),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_901),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_860),
.A2(n_47),
.B(n_48),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_849),
.B(n_47),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_909),
.A2(n_72),
.B1(n_51),
.B2(n_54),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_779),
.B(n_49),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_922),
.B(n_49),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_816),
.B(n_51),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_917),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_892),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_912),
.A2(n_925),
.B(n_919),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_938),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_858),
.B(n_58),
.C(n_59),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_814),
.B(n_58),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_921),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_1101)
);

AOI33xp33_ASAP7_75t_L g1102 ( 
.A1(n_879),
.A2(n_63),
.A3(n_64),
.B1(n_66),
.B2(n_69),
.B3(n_70),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_785),
.B(n_70),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_887),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_938),
.A2(n_72),
.B(n_913),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_914),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_887),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_894),
.A2(n_792),
.B(n_802),
.C(n_865),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_L g1109 ( 
.A(n_933),
.B(n_927),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_857),
.B(n_928),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_915),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_830),
.A2(n_927),
.B1(n_921),
.B2(n_936),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_933),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_916),
.A2(n_908),
.B(n_901),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_879),
.B(n_933),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_933),
.B(n_839),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_916),
.A2(n_908),
.B(n_868),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_918),
.A2(n_867),
.B(n_868),
.C(n_863),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_863),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_867),
.A2(n_933),
.B1(n_798),
.B2(n_836),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_924),
.A2(n_795),
.B(n_808),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_818),
.B(n_771),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_809),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_1121),
.A2(n_1071),
.B(n_947),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1024),
.A2(n_971),
.B(n_966),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_975),
.A2(n_956),
.B(n_953),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1034),
.B(n_950),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_952),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_956),
.A2(n_953),
.B(n_976),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_967),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_1009),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_939),
.A2(n_944),
.B(n_982),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1006),
.B(n_1074),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1014),
.A2(n_1056),
.B(n_939),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_978),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_963),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_1014),
.A2(n_959),
.B(n_958),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_1087),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_945),
.B(n_1051),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1003),
.B(n_1106),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1083),
.A2(n_947),
.B(n_1110),
.C(n_1015),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_944),
.A2(n_946),
.B(n_1000),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_993),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_980),
.A2(n_1102),
.B(n_965),
.C(n_1100),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1068),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1021),
.B(n_973),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_1115),
.B(n_949),
.Y(n_1148)
);

BUFx12f_ASAP7_75t_L g1149 ( 
.A(n_1011),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_977),
.A2(n_946),
.A3(n_1118),
.B(n_1066),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1095),
.B(n_991),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_963),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_963),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_SL g1154 ( 
.A1(n_1105),
.A2(n_1082),
.B(n_970),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1000),
.A2(n_974),
.B(n_1116),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_1047),
.B(n_960),
.C(n_961),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1122),
.B(n_1120),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_940),
.B(n_1038),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1114),
.A2(n_1113),
.B(n_1097),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_943),
.B(n_1050),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_992),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1036),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1020),
.A2(n_1070),
.B1(n_1004),
.B2(n_942),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1117),
.A2(n_1085),
.B(n_1098),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1117),
.A2(n_998),
.B(n_990),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_1052),
.B(n_1081),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1111),
.B(n_951),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_969),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1074),
.B(n_1008),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1119),
.A2(n_972),
.B(n_1108),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_986),
.A2(n_985),
.B(n_987),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_995),
.B(n_988),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1039),
.B(n_1040),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1084),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_981),
.A2(n_989),
.B(n_1002),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1054),
.B(n_964),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1052),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_999),
.A2(n_1001),
.B(n_1005),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1052),
.B(n_1081),
.Y(n_1180)
);

AND3x1_ASAP7_75t_SL g1181 ( 
.A(n_1057),
.B(n_1078),
.C(n_955),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1099),
.B(n_1092),
.C(n_1030),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1081),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1063),
.A2(n_1123),
.B(n_1018),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_943),
.B(n_1035),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_941),
.B(n_1072),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1010),
.B(n_1016),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_968),
.A2(n_979),
.B(n_996),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_941),
.A2(n_1027),
.B1(n_1026),
.B2(n_1073),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1076),
.A2(n_1086),
.B(n_1090),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1063),
.A2(n_1048),
.B(n_1065),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1041),
.B(n_1022),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1007),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1073),
.A2(n_1033),
.B(n_1028),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_1042),
.A2(n_1044),
.B(n_1037),
.Y(n_1195)
);

AO21x1_ASAP7_75t_L g1196 ( 
.A1(n_1049),
.A2(n_1105),
.B(n_1053),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1058),
.A2(n_1060),
.B(n_1064),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_994),
.A2(n_1112),
.B(n_1080),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1023),
.B(n_1029),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1093),
.A2(n_1053),
.B(n_1103),
.C(n_1069),
.Y(n_1201)
);

CKINVDCx8_ASAP7_75t_R g1202 ( 
.A(n_1008),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1096),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1023),
.B(n_1025),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_948),
.A2(n_1094),
.B(n_1061),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_954),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1096),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_984),
.A2(n_1012),
.B(n_1013),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1043),
.A2(n_1045),
.B(n_1046),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1104),
.B(n_1107),
.Y(n_1210)
);

NAND2x1_ASAP7_75t_L g1211 ( 
.A(n_1096),
.B(n_1087),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1031),
.B(n_1046),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1059),
.A2(n_1019),
.B(n_997),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1013),
.B(n_1012),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1079),
.A2(n_1101),
.B(n_1062),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1091),
.A2(n_1032),
.B(n_1089),
.Y(n_1216)
);

AOI33xp33_ASAP7_75t_L g1217 ( 
.A1(n_1017),
.A2(n_1088),
.A3(n_1055),
.B1(n_1008),
.B2(n_1074),
.B3(n_1087),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1067),
.A2(n_957),
.B(n_1087),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1067),
.B(n_1087),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1034),
.B(n_950),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_945),
.B(n_950),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_978),
.B(n_1051),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1034),
.B(n_950),
.Y(n_1223)
);

CKINVDCx8_ASAP7_75t_R g1224 ( 
.A(n_1011),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_973),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1034),
.B(n_950),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1034),
.B(n_950),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_945),
.A2(n_974),
.B(n_970),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_945),
.A2(n_947),
.B(n_795),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1075),
.A2(n_808),
.B(n_939),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1006),
.B(n_1074),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_952),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_978),
.B(n_1051),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1074),
.B(n_830),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1036),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_978),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_945),
.B(n_950),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1087),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1034),
.B(n_950),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1034),
.B(n_950),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1034),
.B(n_950),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_945),
.A2(n_1034),
.B1(n_1083),
.B2(n_629),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_945),
.A2(n_876),
.B(n_1034),
.C(n_1083),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1250)
);

BUFx5_ASAP7_75t_L g1251 ( 
.A(n_1087),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_978),
.B(n_1051),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1036),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_952),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_945),
.A2(n_947),
.B(n_795),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1034),
.B(n_950),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_993),
.Y(n_1258)
);

CKINVDCx8_ASAP7_75t_R g1259 ( 
.A(n_1011),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_945),
.A2(n_876),
.B(n_1034),
.C(n_1083),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1095),
.B(n_902),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_978),
.B(n_1051),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1034),
.B(n_950),
.Y(n_1265)
);

OA22x2_ASAP7_75t_L g1266 ( 
.A1(n_1034),
.A2(n_579),
.B1(n_533),
.B2(n_936),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_SL g1267 ( 
.A1(n_945),
.A2(n_974),
.B(n_970),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_963),
.B(n_1052),
.Y(n_1268)
);

OAI21xp33_ASAP7_75t_L g1269 ( 
.A1(n_1034),
.A2(n_1015),
.B(n_629),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1034),
.B(n_950),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1036),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_945),
.A2(n_947),
.B(n_795),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_952),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1024),
.A2(n_962),
.B(n_1075),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_945),
.B(n_950),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1009),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1009),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1006),
.B(n_1074),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1034),
.B(n_950),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_SL g1282 ( 
.A1(n_1121),
.A2(n_1071),
.B(n_947),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_963),
.B(n_1052),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_947),
.A2(n_950),
.B(n_944),
.Y(n_1284)
);

OR2x2_ASAP7_75t_SL g1285 ( 
.A(n_1172),
.B(n_1156),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1248),
.A2(n_1141),
.B1(n_1260),
.B2(n_1249),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1128),
.B(n_1220),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1269),
.A2(n_1151),
.B1(n_1157),
.B2(n_1147),
.Y(n_1289)
);

INVx6_ASAP7_75t_L g1290 ( 
.A(n_1237),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1222),
.B(n_1236),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1152),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1146),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1225),
.B(n_1173),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1216),
.A2(n_1209),
.B(n_1256),
.C(n_1274),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1252),
.B(n_1264),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1253),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1185),
.B(n_1136),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1136),
.B(n_1239),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1228),
.B(n_1244),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1238),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1258),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1152),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1152),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1249),
.A2(n_1260),
.B1(n_1281),
.B2(n_1271),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1257),
.B(n_1265),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1215),
.A2(n_1182),
.B1(n_1195),
.B2(n_1266),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1132),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1158),
.B(n_1167),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1142),
.A2(n_1187),
.B(n_1277),
.C(n_1140),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1125),
.A2(n_1282),
.B(n_1232),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1258),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1239),
.B(n_1187),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1152),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1278),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1142),
.B(n_1163),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1206),
.A2(n_1148),
.B(n_1171),
.C(n_1190),
.Y(n_1321)
);

INVxp67_ASAP7_75t_SL g1322 ( 
.A(n_1166),
.Y(n_1322)
);

NOR2xp67_ASAP7_75t_SL g1323 ( 
.A(n_1139),
.B(n_1242),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1277),
.B(n_1212),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1279),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1129),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1160),
.B(n_1210),
.Y(n_1327)
);

AOI222xp33_ASAP7_75t_L g1328 ( 
.A1(n_1149),
.A2(n_1157),
.B1(n_1192),
.B2(n_1145),
.C1(n_1263),
.C2(n_1266),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1139),
.A2(n_1242),
.B1(n_1251),
.B2(n_1144),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1134),
.A2(n_1280),
.B1(n_1234),
.B2(n_1189),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1145),
.A2(n_1284),
.B(n_1262),
.C(n_1261),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1161),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1273),
.Y(n_1334)
);

OAI21xp33_ASAP7_75t_L g1335 ( 
.A1(n_1204),
.A2(n_1200),
.B(n_1198),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1174),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1177),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1190),
.B(n_1186),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1229),
.A2(n_1267),
.B1(n_1139),
.B2(n_1242),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1144),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1134),
.B(n_1234),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1280),
.B(n_1170),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1231),
.A2(n_1247),
.B(n_1262),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1131),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1169),
.B(n_1139),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1168),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1177),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1178),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1235),
.B(n_1255),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1275),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1205),
.A2(n_1201),
.B(n_1197),
.C(n_1196),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1231),
.A2(n_1261),
.B(n_1241),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1155),
.A2(n_1205),
.B(n_1217),
.C(n_1201),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1242),
.A2(n_1155),
.B1(n_1175),
.B2(n_1176),
.Y(n_1354)
);

OR2x2_ASAP7_75t_SL g1355 ( 
.A(n_1181),
.B(n_1259),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1183),
.B(n_1203),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1217),
.B(n_1251),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1251),
.A2(n_1181),
.B1(n_1154),
.B2(n_1224),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1202),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1177),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1208),
.A2(n_1218),
.B(n_1214),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1251),
.B(n_1203),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1137),
.B(n_1153),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1137),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1251),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1251),
.B(n_1183),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1180),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1180),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1208),
.A2(n_1143),
.B1(n_1193),
.B2(n_1164),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1191),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1268),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1153),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1143),
.A2(n_1218),
.B(n_1176),
.C(n_1188),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1184),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1219),
.A2(n_1283),
.B(n_1268),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1219),
.A2(n_1283),
.B(n_1194),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1207),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1213),
.A2(n_1135),
.B(n_1159),
.C(n_1138),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1207),
.B(n_1150),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1150),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1165),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1150),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1150),
.B(n_1219),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1133),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1233),
.B(n_1124),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1126),
.B(n_1243),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1226),
.B(n_1250),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1179),
.B(n_1130),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1127),
.B(n_1270),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1230),
.A2(n_1254),
.B1(n_1272),
.B2(n_1276),
.Y(n_1390)
);

NAND2x1_ASAP7_75t_L g1391 ( 
.A(n_1183),
.B(n_1063),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1225),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1269),
.B(n_1034),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1166),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1147),
.B(n_978),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1211),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1269),
.B(n_1034),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1162),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1211),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1156),
.B(n_905),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1258),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1161),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1129),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1129),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1161),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1248),
.A2(n_945),
.B(n_1260),
.C(n_1249),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1269),
.B(n_1034),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1225),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1128),
.B(n_1220),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1196),
.A2(n_945),
.B(n_1199),
.C(n_1034),
.Y(n_1413)
);

AOI21xp33_ASAP7_75t_L g1414 ( 
.A1(n_1269),
.A2(n_1034),
.B(n_945),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1147),
.B(n_978),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1132),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1269),
.A2(n_807),
.B1(n_991),
.B2(n_988),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1418)
);

NOR2x1_ASAP7_75t_L g1419 ( 
.A(n_1258),
.B(n_1144),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1129),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_SL g1421 ( 
.A(n_1269),
.B(n_1034),
.C(n_945),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1128),
.B(n_1220),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1269),
.A2(n_1248),
.B1(n_876),
.B2(n_1034),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1248),
.A2(n_945),
.B1(n_1141),
.B2(n_1034),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_SL g1425 ( 
.A(n_1258),
.B(n_902),
.Y(n_1425)
);

BUFx4f_ASAP7_75t_L g1426 ( 
.A(n_1178),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1147),
.B(n_978),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1428)
);

HAxp5_ASAP7_75t_L g1429 ( 
.A(n_1181),
.B(n_406),
.CON(n_1429),
.SN(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1152),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1129),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1199),
.A2(n_1240),
.B(n_1221),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1196),
.A2(n_945),
.B(n_1199),
.C(n_1034),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1129),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1225),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1128),
.B(n_1220),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1136),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1237),
.B(n_1169),
.Y(n_1438)
);

OR2x6_ASAP7_75t_SL g1439 ( 
.A(n_1146),
.B(n_902),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1129),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1392),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1323),
.B(n_1380),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1291),
.B(n_1297),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1319),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1311),
.B(n_1299),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1349),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1345),
.Y(n_1448)
);

AO21x1_ASAP7_75t_SL g1449 ( 
.A1(n_1311),
.A2(n_1357),
.B(n_1382),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1417),
.A2(n_1355),
.B1(n_1285),
.B2(n_1358),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1324),
.B(n_1320),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1350),
.Y(n_1452)
);

AO21x1_ASAP7_75t_SL g1453 ( 
.A1(n_1414),
.A2(n_1379),
.B(n_1338),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1326),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1430),
.Y(n_1455)
);

OA21x2_ASAP7_75t_L g1456 ( 
.A1(n_1343),
.A2(n_1352),
.B(n_1353),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1345),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1423),
.B(n_1320),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1393),
.A2(n_1409),
.B1(n_1397),
.B2(n_1424),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1344),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1313),
.A2(n_1309),
.B1(n_1287),
.B2(n_1411),
.Y(n_1461)
);

AO21x1_ASAP7_75t_L g1462 ( 
.A1(n_1286),
.A2(n_1310),
.B(n_1304),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1319),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1423),
.B(n_1393),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1303),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1325),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1390),
.A2(n_1361),
.B(n_1385),
.Y(n_1467)
);

AOI222xp33_ASAP7_75t_L g1468 ( 
.A1(n_1421),
.A2(n_1409),
.B1(n_1397),
.B2(n_1415),
.C1(n_1427),
.C2(n_1395),
.Y(n_1468)
);

NOR2x1_ASAP7_75t_SL g1469 ( 
.A(n_1339),
.B(n_1293),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1425),
.A2(n_1290),
.B1(n_1308),
.B2(n_1412),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1421),
.A2(n_1328),
.B1(n_1358),
.B2(n_1342),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1353),
.A2(n_1413),
.B(n_1433),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1325),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1389),
.A2(n_1378),
.B(n_1388),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1346),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1388),
.A2(n_1389),
.B(n_1408),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1410),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1430),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1392),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1288),
.B(n_1301),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1396),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1306),
.A2(n_1422),
.B1(n_1436),
.B2(n_1289),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1401),
.A2(n_1317),
.B1(n_1315),
.B2(n_1295),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1329),
.B(n_1398),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1331),
.A2(n_1293),
.B1(n_1435),
.B2(n_1359),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1413),
.A2(n_1433),
.B(n_1332),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1396),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1381),
.A2(n_1432),
.B(n_1428),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1296),
.A2(n_1321),
.B1(n_1407),
.B2(n_1335),
.C(n_1341),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1317),
.A2(n_1315),
.B1(n_1438),
.B2(n_1412),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1400),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1333),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1407),
.A2(n_1312),
.B1(n_1290),
.B2(n_1365),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1381),
.A2(n_1418),
.B(n_1387),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1336),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1416),
.Y(n_1496)
);

BUFx12f_ASAP7_75t_L g1497 ( 
.A(n_1316),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1290),
.Y(n_1498)
);

AO21x1_ASAP7_75t_L g1499 ( 
.A1(n_1351),
.A2(n_1314),
.B(n_1354),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1327),
.B(n_1300),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1336),
.Y(n_1501)
);

HB1xp67_ASAP7_75t_L g1502 ( 
.A(n_1312),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1437),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1403),
.Y(n_1504)
);

CKINVDCx11_ASAP7_75t_R g1505 ( 
.A(n_1439),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1437),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1400),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1293),
.A2(n_1330),
.B1(n_1359),
.B2(n_1398),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1360),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1404),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1405),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1406),
.A2(n_1340),
.B1(n_1402),
.B2(n_1366),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1330),
.A2(n_1438),
.B1(n_1329),
.B2(n_1394),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1292),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1429),
.A2(n_1426),
.B1(n_1383),
.B2(n_1322),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1420),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1292),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1292),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1322),
.A2(n_1394),
.B1(n_1434),
.B2(n_1431),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1429),
.A2(n_1426),
.B1(n_1348),
.B2(n_1296),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1419),
.A2(n_1334),
.B1(n_1302),
.B2(n_1440),
.Y(n_1521)
);

BUFx2_ASAP7_75t_R g1522 ( 
.A(n_1348),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1292),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_SL g1524 ( 
.A1(n_1367),
.A2(n_1377),
.B1(n_1294),
.B2(n_1368),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1356),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1370),
.B(n_1384),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1386),
.A2(n_1369),
.B(n_1374),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1356),
.Y(n_1528)
);

BUFx4f_ASAP7_75t_SL g1529 ( 
.A(n_1318),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1298),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1369),
.A2(n_1376),
.B(n_1375),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1363),
.Y(n_1532)
);

BUFx8_ASAP7_75t_L g1533 ( 
.A(n_1318),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1399),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1378),
.A2(n_1373),
.B(n_1332),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1362),
.B(n_1371),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1318),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1367),
.A2(n_1372),
.B1(n_1364),
.B2(n_1371),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1391),
.A2(n_1373),
.B(n_1305),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1307),
.A2(n_1318),
.B1(n_1337),
.B2(n_1347),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1337),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1337),
.B(n_1347),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1337),
.Y(n_1543)
);

BUFx8_ASAP7_75t_L g1544 ( 
.A(n_1347),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1321),
.B(n_1347),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1313),
.B(n_1287),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1349),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1349),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1417),
.A2(n_945),
.B1(n_1248),
.B2(n_1141),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1313),
.B(n_1287),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1349),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1430),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1392),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1320),
.A2(n_1083),
.B1(n_1269),
.B2(n_1004),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1349),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1324),
.B(n_1320),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1349),
.Y(n_1557)
);

BUFx2_ASAP7_75t_R g1558 ( 
.A(n_1439),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1320),
.A2(n_807),
.B1(n_1003),
.B2(n_991),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1349),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1417),
.A2(n_807),
.B1(n_991),
.B2(n_598),
.Y(n_1561)
);

INVx5_ASAP7_75t_SL g1562 ( 
.A(n_1293),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1303),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1410),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1349),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1303),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1320),
.A2(n_807),
.B1(n_1003),
.B2(n_991),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1303),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1349),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1349),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1349),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1417),
.A2(n_945),
.B1(n_1248),
.B2(n_1141),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1423),
.A2(n_945),
.B(n_1034),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1392),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1349),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1430),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1349),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1417),
.A2(n_945),
.B1(n_1248),
.B2(n_1141),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1430),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1349),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1319),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1320),
.A2(n_1083),
.B1(n_1269),
.B2(n_1004),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1410),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1423),
.A2(n_945),
.B(n_1034),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1349),
.Y(n_1585)
);

BUFx12f_ASAP7_75t_L g1586 ( 
.A(n_1303),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1320),
.A2(n_1083),
.B1(n_1269),
.B2(n_1004),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1458),
.B(n_1464),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1480),
.B(n_1461),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1526),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1545),
.Y(n_1591)
);

BUFx4f_ASAP7_75t_SL g1592 ( 
.A(n_1497),
.Y(n_1592)
);

INVxp67_ASAP7_75t_R g1593 ( 
.A(n_1531),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1480),
.B(n_1546),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1526),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1533),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1526),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1466),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1473),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1550),
.B(n_1482),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1451),
.B(n_1556),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1476),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1458),
.B(n_1464),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1446),
.B(n_1449),
.Y(n_1604)
);

BUFx5_ASAP7_75t_L g1605 ( 
.A(n_1452),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1527),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1451),
.B(n_1556),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1527),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1559),
.A2(n_1567),
.B1(n_1450),
.B2(n_1561),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1499),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1499),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1477),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1573),
.A2(n_1584),
.B(n_1459),
.Y(n_1613)
);

AO31x2_ASAP7_75t_L g1614 ( 
.A1(n_1462),
.A2(n_1578),
.A3(n_1549),
.B(n_1572),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1446),
.B(n_1449),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1456),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1472),
.Y(n_1617)
);

INVx2_ASAP7_75t_SL g1618 ( 
.A(n_1473),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1531),
.B(n_1462),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1581),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1486),
.B(n_1483),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1536),
.B(n_1453),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1533),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1535),
.B(n_1489),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1535),
.B(n_1490),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1536),
.B(n_1453),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1468),
.B(n_1447),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1495),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1506),
.B(n_1562),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1501),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1445),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1547),
.B(n_1548),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1551),
.B(n_1555),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1557),
.B(n_1560),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1554),
.A2(n_1587),
.B1(n_1582),
.B2(n_1470),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1539),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1562),
.B(n_1500),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1469),
.B(n_1448),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1463),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1565),
.B(n_1569),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1454),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1467),
.A2(n_1488),
.B(n_1494),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1532),
.B(n_1441),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1460),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1475),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1443),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1478),
.A2(n_1579),
.B(n_1552),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1539),
.A2(n_1471),
.B(n_1511),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1474),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1519),
.A2(n_1493),
.B(n_1510),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1479),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1516),
.A2(n_1530),
.B(n_1534),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1575),
.B(n_1577),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1442),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1553),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1574),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1580),
.B(n_1585),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1533),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1502),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1444),
.B(n_1564),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1538),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1481),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1544),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1484),
.B(n_1562),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1583),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1513),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1487),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1485),
.A2(n_1508),
.B(n_1540),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1628),
.B(n_1562),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1640),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1657),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1496),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1588),
.B(n_1515),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1643),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1640),
.B(n_1498),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1625),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1588),
.B(n_1520),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1603),
.B(n_1541),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1643),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1626),
.B(n_1484),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1647),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1625),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1649),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1618),
.Y(n_1691)
);

OAI33xp33_ASAP7_75t_L g1692 ( 
.A1(n_1609),
.A2(n_1512),
.A3(n_1543),
.B1(n_1465),
.B2(n_1566),
.B3(n_1521),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1603),
.B(n_1518),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1637),
.B(n_1524),
.C(n_1505),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1604),
.B(n_1518),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1609),
.A2(n_1505),
.B1(n_1586),
.B2(n_1497),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1604),
.B(n_1518),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1615),
.B(n_1542),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1618),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1594),
.B(n_1492),
.Y(n_1700)
);

INVx5_ASAP7_75t_L g1701 ( 
.A(n_1638),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1640),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1612),
.B(n_1465),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1617),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1620),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1591),
.B(n_1509),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1615),
.B(n_1542),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1566),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1670),
.B(n_1568),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1591),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1638),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1613),
.A2(n_1586),
.B1(n_1504),
.B2(n_1563),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1600),
.B(n_1568),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1607),
.B(n_1504),
.Y(n_1714)
);

BUFx12f_ASAP7_75t_L g1715 ( 
.A(n_1650),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1622),
.B(n_1523),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1627),
.B(n_1523),
.Y(n_1717)
);

INVx6_ASAP7_75t_L g1718 ( 
.A(n_1646),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1621),
.B(n_1525),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1659),
.B(n_1590),
.Y(n_1720)
);

INVxp67_ASAP7_75t_SL g1721 ( 
.A(n_1630),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1620),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1645),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1627),
.B(n_1523),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1656),
.Y(n_1725)
);

OAI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1589),
.A2(n_1525),
.B1(n_1528),
.B2(n_1491),
.C(n_1507),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1629),
.A2(n_1563),
.B1(n_1528),
.B2(n_1507),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1601),
.B(n_1517),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1621),
.B(n_1491),
.Y(n_1729)
);

NAND4xp25_ASAP7_75t_L g1730 ( 
.A(n_1629),
.B(n_1537),
.C(n_1558),
.D(n_1579),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1660),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1661),
.B(n_1664),
.Y(n_1732)
);

NOR4xp25_ASAP7_75t_SL g1733 ( 
.A(n_1671),
.B(n_1522),
.C(n_1443),
.D(n_1544),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1624),
.B(n_1517),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1590),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1624),
.B(n_1514),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_SL g1737 ( 
.A(n_1692),
.B(n_1666),
.C(n_1611),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1611),
.C(n_1610),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1694),
.A2(n_1671),
.B1(n_1619),
.B2(n_1610),
.C(n_1639),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1694),
.B(n_1632),
.C(n_1633),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1725),
.A2(n_1641),
.B1(n_1634),
.B2(n_1648),
.C(n_1635),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_L g1743 ( 
.A(n_1712),
.B(n_1639),
.C(n_1599),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1723),
.B(n_1598),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1727),
.A2(n_1596),
.B1(n_1668),
.B2(n_1663),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_SL g1746 ( 
.A1(n_1727),
.A2(n_1683),
.B1(n_1726),
.B2(n_1619),
.C(n_1679),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1734),
.B(n_1619),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1683),
.A2(n_1619),
.B1(n_1631),
.B2(n_1614),
.C(n_1635),
.Y(n_1748)
);

NOR2xp67_ASAP7_75t_L g1749 ( 
.A(n_1701),
.B(n_1602),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1713),
.A2(n_1623),
.B1(n_1663),
.B2(n_1668),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1731),
.B(n_1619),
.C(n_1653),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1734),
.B(n_1593),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1736),
.B(n_1593),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1732),
.B(n_1614),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1680),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1706),
.B(n_1646),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1673),
.B1(n_1646),
.B2(n_1651),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1676),
.B(n_1606),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1614),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1678),
.B(n_1614),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1676),
.B(n_1702),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1676),
.B(n_1608),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1679),
.A2(n_1714),
.B(n_1700),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1678),
.B(n_1614),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1685),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1728),
.B(n_1614),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1695),
.B(n_1697),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1706),
.B(n_1646),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1733),
.A2(n_1623),
.B1(n_1663),
.B2(n_1596),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1682),
.B(n_1655),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1689),
.A2(n_1634),
.B1(n_1636),
.B2(n_1658),
.C(n_1648),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_L g1772 ( 
.A(n_1708),
.B(n_1653),
.C(n_1658),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1697),
.B(n_1720),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1720),
.B(n_1616),
.Y(n_1774)
);

NAND3xp33_ASAP7_75t_L g1775 ( 
.A(n_1703),
.B(n_1653),
.C(n_1662),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1693),
.B(n_1655),
.Y(n_1776)
);

NOR3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1709),
.B(n_1595),
.C(n_1597),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1693),
.B(n_1636),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1718),
.B(n_1592),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1720),
.B(n_1716),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1691),
.B(n_1653),
.C(n_1699),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1686),
.A2(n_1673),
.B1(n_1651),
.B2(n_1669),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_L g1783 ( 
.A(n_1705),
.B(n_1642),
.C(n_1662),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1720),
.B(n_1602),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1717),
.B(n_1724),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1722),
.B(n_1642),
.C(n_1672),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1686),
.A2(n_1673),
.B1(n_1651),
.B2(n_1669),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1724),
.B(n_1595),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1684),
.B(n_1605),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1684),
.B(n_1605),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1719),
.A2(n_1623),
.B1(n_1596),
.B2(n_1668),
.Y(n_1791)
);

OA21x2_ASAP7_75t_L g1792 ( 
.A1(n_1677),
.A2(n_1644),
.B(n_1654),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1710),
.B(n_1597),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1719),
.B(n_1672),
.C(n_1667),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1718),
.B(n_1651),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_SL g1796 ( 
.A1(n_1740),
.A2(n_1715),
.B1(n_1718),
.B2(n_1707),
.Y(n_1796)
);

AND2x4_ASAP7_75t_SL g1797 ( 
.A(n_1777),
.B(n_1681),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1741),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1741),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1754),
.B(n_1685),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1760),
.B(n_1687),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1773),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1755),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1767),
.B(n_1675),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.B(n_1675),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1755),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1764),
.B(n_1687),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1744),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1765),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1740),
.B(n_1681),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1765),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1774),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1774),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1815)
);

INVxp67_ASAP7_75t_SL g1816 ( 
.A(n_1786),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1793),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1776),
.B(n_1729),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1766),
.B(n_1674),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1785),
.B(n_1698),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1749),
.B(n_1701),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1770),
.B(n_1688),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1759),
.B(n_1704),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1792),
.Y(n_1824)
);

NOR2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1738),
.B(n_1715),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1793),
.Y(n_1826)
);

BUFx3_ASAP7_75t_L g1827 ( 
.A(n_1779),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1758),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1749),
.B(n_1701),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1775),
.B(n_1704),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1752),
.B(n_1707),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1763),
.B(n_1690),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1752),
.B(n_1735),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1811),
.B(n_1761),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1808),
.B(n_1763),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1816),
.B(n_1775),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1830),
.B(n_1772),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1830),
.B(n_1772),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1799),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1799),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1825),
.A2(n_1738),
.B1(n_1745),
.B2(n_1743),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1815),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1761),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1799),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1818),
.B(n_1783),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1806),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1806),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1806),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1824),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1821),
.B(n_1783),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1810),
.A2(n_1743),
.B(n_1739),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1796),
.B(n_1750),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1821),
.B(n_1786),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1798),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1832),
.B(n_1778),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1796),
.A2(n_1746),
.B(n_1751),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1818),
.B(n_1748),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1832),
.B(n_1742),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1819),
.B(n_1789),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1797),
.A2(n_1751),
.B(n_1756),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1798),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1803),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1804),
.B(n_1753),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1819),
.B(n_1790),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1804),
.B(n_1753),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1794),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1805),
.B(n_1784),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1827),
.B(n_1768),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1821),
.B(n_1762),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1802),
.B(n_1788),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1802),
.B(n_1788),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1803),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1821),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1809),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1809),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1801),
.B(n_1771),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1812),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1824),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1869),
.B(n_1813),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1866),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1869),
.B(n_1813),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1850),
.B(n_1829),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1869),
.B(n_1814),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1854),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1847),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1800),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1854),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1837),
.B(n_1800),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1861),
.Y(n_1889)
);

NAND2xp33_ASAP7_75t_L g1890 ( 
.A(n_1851),
.B(n_1825),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1861),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1850),
.B(n_1829),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1873),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1835),
.Y(n_1894)
);

NOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1836),
.B(n_1827),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1876),
.B(n_1820),
.Y(n_1896)
);

NAND2x1_ASAP7_75t_SL g1897 ( 
.A(n_1841),
.B(n_1829),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1866),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1862),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1869),
.B(n_1814),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1847),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1850),
.B(n_1827),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1862),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1872),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1849),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1873),
.B(n_1833),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1872),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1856),
.B(n_1797),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1874),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1874),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1837),
.B(n_1801),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1853),
.B(n_1817),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1875),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1868),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1855),
.B(n_1836),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1849),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1875),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1853),
.B(n_1829),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1877),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1877),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1852),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1857),
.B(n_1831),
.Y(n_1923)
);

AOI21xp33_ASAP7_75t_L g1924 ( 
.A1(n_1838),
.A2(n_1757),
.B(n_1791),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1857),
.B(n_1831),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1860),
.B(n_1797),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1840),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1840),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1902),
.B(n_1853),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1905),
.Y(n_1930)
);

OAI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1922),
.A2(n_1838),
.B1(n_1782),
.B2(n_1787),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1902),
.B(n_1842),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1893),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1919),
.B(n_1842),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1895),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1910),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1888),
.B(n_1845),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1884),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1919),
.B(n_1834),
.Y(n_1939)
);

OAI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1895),
.A2(n_1845),
.B1(n_1864),
.B2(n_1859),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1915),
.B(n_1859),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1882),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1884),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1901),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1894),
.B(n_1870),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1919),
.B(n_1834),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1919),
.B(n_1843),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1887),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1897),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1888),
.B(n_1864),
.Y(n_1950)
);

AO22x1_ASAP7_75t_L g1951 ( 
.A1(n_1880),
.A2(n_1769),
.B1(n_1878),
.B2(n_1863),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1897),
.B(n_1652),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1912),
.B(n_1807),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1882),
.B(n_1839),
.Y(n_1954)
);

INVx1_ASAP7_75t_SL g1955 ( 
.A(n_1909),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1886),
.B(n_1870),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1887),
.Y(n_1957)
);

BUFx2_ASAP7_75t_L g1958 ( 
.A(n_1882),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1912),
.B(n_1807),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1923),
.B(n_1871),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1901),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1898),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1890),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1901),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1906),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1926),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1889),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1882),
.B(n_1843),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1889),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1958),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1938),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1949),
.A2(n_1925),
.B1(n_1896),
.B2(n_1916),
.Y(n_1972)
);

OAI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1935),
.A2(n_1924),
.B1(n_1893),
.B2(n_1781),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1963),
.A2(n_1737),
.B1(n_1781),
.B2(n_1913),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1958),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1938),
.Y(n_1976)
);

OAI222xp33_ASAP7_75t_L g1977 ( 
.A1(n_1955),
.A2(n_1913),
.B1(n_1892),
.B2(n_1907),
.C1(n_1904),
.C2(n_1883),
.Y(n_1977)
);

A2O1A1Ixp33_ASAP7_75t_L g1978 ( 
.A1(n_1966),
.A2(n_1892),
.B(n_1907),
.C(n_1904),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1962),
.B(n_1879),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1943),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1941),
.B(n_1892),
.Y(n_1981)
);

NAND4xp25_ASAP7_75t_L g1982 ( 
.A(n_1937),
.B(n_1892),
.C(n_1881),
.D(n_1883),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1960),
.B(n_1879),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1933),
.Y(n_1984)
);

OAI31xp33_ASAP7_75t_L g1985 ( 
.A1(n_1940),
.A2(n_1900),
.A3(n_1881),
.B(n_1885),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1933),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1942),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1929),
.B(n_1900),
.Y(n_1988)
);

O2A1O1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1931),
.A2(n_1885),
.B(n_1899),
.C(n_1891),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1943),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1932),
.B(n_1871),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1948),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1932),
.B(n_1867),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1945),
.B(n_1937),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1930),
.A2(n_1899),
.B1(n_1891),
.B2(n_1921),
.C(n_1920),
.Y(n_1995)
);

AND3x2_ASAP7_75t_L g1996 ( 
.A(n_1930),
.B(n_1908),
.C(n_1903),
.Y(n_1996)
);

AOI21xp33_ASAP7_75t_SL g1997 ( 
.A1(n_1951),
.A2(n_1952),
.B(n_1942),
.Y(n_1997)
);

OR2x6_ASAP7_75t_L g1998 ( 
.A(n_1952),
.B(n_1652),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1951),
.A2(n_1908),
.B(n_1903),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1984),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1970),
.B(n_1984),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1975),
.B(n_1936),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1988),
.B(n_1929),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1996),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1971),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1986),
.B(n_1936),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1976),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1987),
.B(n_1939),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1980),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1994),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1990),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1978),
.B(n_1939),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1983),
.B(n_1946),
.Y(n_2013)
);

NOR2x1_ASAP7_75t_L g2014 ( 
.A(n_1973),
.B(n_1933),
.Y(n_2014)
);

INVxp33_ASAP7_75t_L g2015 ( 
.A(n_1981),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_1979),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1992),
.B(n_1946),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1993),
.B(n_1947),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1991),
.B(n_1947),
.Y(n_2019)
);

INVxp67_ASAP7_75t_L g2020 ( 
.A(n_1972),
.Y(n_2020)
);

AOI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_1985),
.A2(n_1952),
.B1(n_1968),
.B2(n_1934),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1982),
.B(n_1968),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1974),
.A2(n_1952),
.B1(n_1934),
.B2(n_1950),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1989),
.B(n_1956),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_2014),
.A2(n_1974),
.B(n_1999),
.Y(n_2025)
);

AOI21xp33_ASAP7_75t_L g2026 ( 
.A1(n_2014),
.A2(n_1997),
.B(n_1952),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_2020),
.A2(n_1998),
.B1(n_1995),
.B2(n_1950),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2000),
.B(n_1954),
.Y(n_2028)
);

OAI222xp33_ASAP7_75t_L g2029 ( 
.A1(n_2023),
.A2(n_1998),
.B1(n_1954),
.B2(n_1977),
.C1(n_1953),
.C2(n_1959),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2004),
.A2(n_1998),
.B1(n_1954),
.B2(n_1961),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2004),
.B(n_1954),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2024),
.A2(n_1961),
.B(n_1944),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2001),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_2010),
.B(n_1953),
.Y(n_2034)
);

NOR3x1_ASAP7_75t_L g2035 ( 
.A(n_2006),
.B(n_1957),
.C(n_1948),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2015),
.A2(n_1964),
.B(n_1944),
.Y(n_2036)
);

AOI211xp5_ASAP7_75t_L g2037 ( 
.A1(n_2012),
.A2(n_1964),
.B(n_1967),
.C(n_1957),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_2021),
.A2(n_1969),
.B(n_1967),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2012),
.A2(n_1969),
.B(n_1965),
.C(n_1959),
.Y(n_2039)
);

OAI21xp33_ASAP7_75t_L g2040 ( 
.A1(n_2022),
.A2(n_1965),
.B(n_1914),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2028),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2031),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2033),
.B(n_2010),
.Y(n_2043)
);

NOR3x1_ASAP7_75t_L g2044 ( 
.A(n_2034),
.B(n_2002),
.C(n_2008),
.Y(n_2044)
);

NOR3xp33_ASAP7_75t_SL g2045 ( 
.A(n_2029),
.B(n_2013),
.C(n_2007),
.Y(n_2045)
);

NOR3xp33_ASAP7_75t_L g2046 ( 
.A(n_2025),
.B(n_2016),
.C(n_2007),
.Y(n_2046)
);

AOI21xp33_ASAP7_75t_L g2047 ( 
.A1(n_2027),
.A2(n_2017),
.B(n_2011),
.Y(n_2047)
);

NOR2x1_ASAP7_75t_L g2048 ( 
.A(n_2036),
.B(n_2011),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_2026),
.A2(n_2017),
.B(n_2003),
.Y(n_2049)
);

NOR2xp67_ASAP7_75t_L g2050 ( 
.A(n_2032),
.B(n_2017),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2040),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_L g2052 ( 
.A(n_2038),
.B(n_2005),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2039),
.B(n_2018),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2045),
.A2(n_2030),
.B1(n_2037),
.B2(n_2019),
.C(n_2009),
.Y(n_2054)
);

NOR2xp67_ASAP7_75t_L g2055 ( 
.A(n_2050),
.B(n_2003),
.Y(n_2055)
);

NAND3xp33_ASAP7_75t_SL g2056 ( 
.A(n_2046),
.B(n_2009),
.C(n_2005),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_2042),
.Y(n_2057)
);

AOI211xp5_ASAP7_75t_L g2058 ( 
.A1(n_2047),
.A2(n_2019),
.B(n_2018),
.C(n_2035),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2049),
.B(n_2018),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_2051),
.B(n_2018),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2055),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_2058),
.B(n_2041),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_2059),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2060),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_2054),
.A2(n_2052),
.B1(n_2053),
.B2(n_2056),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2057),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_2057),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2055),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_2063),
.Y(n_2069)
);

OR5x1_ASAP7_75t_L g2070 ( 
.A(n_2065),
.B(n_2044),
.C(n_2048),
.D(n_2043),
.E(n_1906),
.Y(n_2070)
);

OAI31xp33_ASAP7_75t_L g2071 ( 
.A1(n_2061),
.A2(n_1906),
.A3(n_1917),
.B(n_1914),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2068),
.B(n_2064),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_2062),
.B(n_1917),
.C(n_1911),
.Y(n_2073)
);

NAND4xp75_ASAP7_75t_L g2074 ( 
.A(n_2066),
.B(n_1917),
.C(n_1911),
.D(n_1921),
.Y(n_2074)
);

XOR2x2_ASAP7_75t_L g2075 ( 
.A(n_2072),
.B(n_2067),
.Y(n_2075)
);

NOR2x1p5_ASAP7_75t_L g2076 ( 
.A(n_2074),
.B(n_2067),
.Y(n_2076)
);

AND2x4_ASAP7_75t_L g2077 ( 
.A(n_2069),
.B(n_1918),
.Y(n_2077)
);

OAI221xp5_ASAP7_75t_L g2078 ( 
.A1(n_2071),
.A2(n_1920),
.B1(n_1918),
.B2(n_1928),
.C(n_1927),
.Y(n_2078)
);

OAI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_2076),
.A2(n_2073),
.B1(n_1928),
.B2(n_1927),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2075),
.Y(n_2080)
);

NAND5xp2_ASAP7_75t_L g2081 ( 
.A(n_2080),
.B(n_2070),
.C(n_2078),
.D(n_2077),
.E(n_1795),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2081),
.Y(n_2082)
);

OAI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_2081),
.A2(n_2079),
.B1(n_1878),
.B2(n_1839),
.Y(n_2083)
);

AOI22xp5_ASAP7_75t_L g2084 ( 
.A1(n_2082),
.A2(n_1844),
.B1(n_1848),
.B2(n_1846),
.Y(n_2084)
);

AOI21xp33_ASAP7_75t_L g2085 ( 
.A1(n_2083),
.A2(n_1848),
.B(n_1846),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_2084),
.B(n_1844),
.Y(n_2086)
);

AOI21xp33_ASAP7_75t_L g2087 ( 
.A1(n_2086),
.A2(n_2085),
.B(n_1822),
.Y(n_2087)
);

AOI322xp5_ASAP7_75t_L g2088 ( 
.A1(n_2087),
.A2(n_1817),
.A3(n_1826),
.B1(n_1863),
.B2(n_1865),
.C1(n_1824),
.C2(n_1828),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_2088),
.A2(n_1529),
.B1(n_1715),
.B2(n_1824),
.Y(n_2089)
);

AOI211xp5_ASAP7_75t_L g2090 ( 
.A1(n_2089),
.A2(n_1552),
.B(n_1455),
.C(n_1576),
.Y(n_2090)
);


endmodule