module fake_jpeg_810_n_362 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_362);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_362;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_53),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_57),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_30),
.B(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_70),
.Y(n_120)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_67),
.Y(n_127)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_6),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_93),
.Y(n_133)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_9),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_25),
.B(n_9),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_99),
.Y(n_126)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_42),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_27),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_22),
.B(n_10),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_16),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_29),
.B1(n_45),
.B2(n_27),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_103),
.A2(n_104),
.B1(n_112),
.B2(n_122),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_45),
.B1(n_27),
.B2(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_37),
.B1(n_45),
.B2(n_42),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_81),
.B1(n_54),
.B2(n_82),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_40),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_43),
.B1(n_34),
.B2(n_22),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_51),
.A2(n_43),
.B1(n_34),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_36),
.B1(n_33),
.B2(n_21),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_139),
.B1(n_147),
.B2(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_129),
.B(n_144),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_33),
.B1(n_21),
.B2(n_3),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_148),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_50),
.A2(n_21),
.B1(n_33),
.B2(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_11),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_72),
.A2(n_33),
.B1(n_1),
.B2(n_4),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g148 ( 
.A(n_94),
.B(n_2),
.CON(n_148),
.SN(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_66),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_56),
.B(n_5),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_58),
.A2(n_14),
.B1(n_16),
.B2(n_63),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_149),
.B1(n_147),
.B2(n_104),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_16),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_102),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_68),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_166),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_179),
.B1(n_181),
.B2(n_186),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_60),
.B1(n_91),
.B2(n_75),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_178),
.Y(n_208)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_173),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_96),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_174),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_96),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_177),
.C(n_200),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_110),
.A2(n_64),
.B(n_92),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_78),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_103),
.A2(n_86),
.B1(n_90),
.B2(n_77),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_185),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_106),
.A2(n_150),
.B1(n_123),
.B2(n_135),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_184),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_141),
.B1(n_101),
.B2(n_125),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_126),
.A2(n_154),
.B1(n_134),
.B2(n_139),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_153),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_111),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_192),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_137),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_195),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_107),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_140),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_146),
.B1(n_156),
.B2(n_157),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_132),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_107),
.A2(n_108),
.B1(n_101),
.B2(n_142),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_136),
.B1(n_148),
.B2(n_117),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_205),
.A2(n_231),
.B1(n_200),
.B2(n_193),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_159),
.B(n_122),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_209),
.C(n_222),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_140),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_166),
.A2(n_198),
.B1(n_162),
.B2(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_226),
.B1(n_175),
.B2(n_163),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_152),
.C(n_136),
.Y(n_222)
);

BUFx24_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_157),
.B1(n_156),
.B2(n_140),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_229),
.A2(n_203),
.B1(n_218),
.B2(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_156),
.B1(n_157),
.B2(n_185),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_SL g232 ( 
.A(n_170),
.B(n_190),
.C(n_177),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_191),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_228),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_234),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_189),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_235),
.B(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

O2A1O1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_185),
.B(n_175),
.C(n_188),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_206),
.B(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_256),
.Y(n_275)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_171),
.B1(n_172),
.B2(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_248),
.B(n_231),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_227),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_250),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_203),
.A2(n_200),
.B(n_174),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_167),
.C(n_164),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_161),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_219),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_169),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_255),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_183),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_205),
.A2(n_168),
.B1(n_176),
.B2(n_184),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_184),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_265),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_225),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_252),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_271),
.B(n_273),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_237),
.A2(n_220),
.B(n_213),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_225),
.B(n_222),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_274),
.A2(n_240),
.B(n_255),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_241),
.A2(n_207),
.B(n_217),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_239),
.B(n_204),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_243),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_207),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_253),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_240),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_295),
.C(n_280),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_293),
.Y(n_310)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_244),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_256),
.B1(n_254),
.B2(n_238),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_298),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_260),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_303),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_274),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_311),
.C(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_282),
.B(n_270),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_312),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_258),
.C(n_260),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_258),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_306),
.A2(n_294),
.B1(n_287),
.B2(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_306),
.A2(n_287),
.B1(n_277),
.B2(n_265),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_283),
.C(n_264),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_325),
.C(n_308),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_283),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_313),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_263),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_326),
.Y(n_334)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_263),
.C(n_271),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_309),
.Y(n_326)
);

OAI321xp33_ASAP7_75t_L g341 ( 
.A1(n_328),
.A2(n_273),
.A3(n_278),
.B1(n_279),
.B2(n_288),
.C(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_321),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_319),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_337),
.B(n_331),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_319),
.A3(n_318),
.B1(n_317),
.B2(n_307),
.C(n_305),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_333),
.B(n_318),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_343),
.Y(n_347)
);

AOI31xp33_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_342),
.A3(n_327),
.B(n_314),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_334),
.A2(n_317),
.B(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_346),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_348),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_330),
.C(n_332),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_327),
.C(n_296),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_338),
.A2(n_293),
.B1(n_267),
.B2(n_259),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_349),
.B(n_275),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_347),
.B(n_210),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g357 ( 
.A1(n_350),
.A2(n_352),
.B(n_212),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_275),
.B(n_202),
.Y(n_352)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_254),
.B(n_210),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_356),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_217),
.C(n_254),
.Y(n_356)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_357),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_353),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_358),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_212),
.Y(n_362)
);


endmodule