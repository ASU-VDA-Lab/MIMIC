module fake_jpeg_14762_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_27),
.Y(n_111)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_34),
.CON(n_68),
.SN(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_25),
.B(n_26),
.C(n_43),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_24),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_91),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_50),
.A2(n_44),
.B1(n_30),
.B2(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_30),
.B1(n_44),
.B2(n_39),
.Y(n_101)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_28),
.Y(n_91)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_99),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_91),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_115),
.B1(n_119),
.B2(n_76),
.Y(n_157)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_30),
.B1(n_44),
.B2(n_24),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_105),
.B1(n_125),
.B2(n_76),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_39),
.B1(n_23),
.B2(n_25),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g141 ( 
.A(n_107),
.Y(n_141)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_111),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_117),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_68),
.B(n_58),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_123),
.B(n_57),
.C(n_47),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_56),
.B1(n_47),
.B2(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_62),
.Y(n_120)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g151 ( 
.A(n_121),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_39),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_55),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_32),
.B1(n_26),
.B2(n_43),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_27),
.B(n_37),
.C(n_38),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_41),
.Y(n_138)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_133),
.Y(n_164)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_135),
.B1(n_139),
.B2(n_156),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_146),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_69),
.B1(n_116),
.B2(n_127),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_97),
.B1(n_89),
.B2(n_127),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_157),
.B1(n_123),
.B2(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_92),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_150),
.Y(n_180)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_129),
.C(n_134),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_169),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_153),
.B1(n_133),
.B2(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_168),
.B1(n_175),
.B2(n_143),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_163),
.B1(n_111),
.B2(n_118),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_120),
.B1(n_103),
.B2(n_99),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_113),
.B1(n_103),
.B2(n_123),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_114),
.C(n_55),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_114),
.C(n_77),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_109),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_122),
.B1(n_111),
.B2(n_124),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_182),
.B(n_193),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_190),
.B1(n_191),
.B2(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_151),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_176),
.B(n_178),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_110),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_96),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_139),
.B1(n_131),
.B2(n_158),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_124),
.B1(n_143),
.B2(n_144),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_195),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_126),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_167),
.B1(n_142),
.B2(n_166),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_101),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_198),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_137),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_165),
.B(n_168),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_203),
.A2(n_217),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_181),
.B(n_162),
.CI(n_172),
.CON(n_205),
.SN(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_194),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_207),
.A2(n_215),
.B1(n_219),
.B2(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_209),
.C(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_176),
.C(n_137),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_184),
.B(n_191),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_178),
.C(n_57),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_29),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_183),
.Y(n_232)
);

AOI22x1_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_141),
.B1(n_167),
.B2(n_179),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_26),
.B(n_43),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_141),
.B(n_155),
.C(n_70),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_141),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_196),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_182),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_41),
.B1(n_38),
.B2(n_37),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_193),
.B1(n_35),
.B2(n_33),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_236),
.C(n_212),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_227),
.A2(n_230),
.B(n_241),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_229),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_187),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_234),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_240),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_215),
.B1(n_217),
.B2(n_205),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_249),
.B1(n_211),
.B2(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

XNOR2x2_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_192),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_205),
.A2(n_191),
.B1(n_190),
.B2(n_199),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_197),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_269),
.C(n_256),
.Y(n_281)
);

OA21x2_ASAP7_75t_L g253 ( 
.A1(n_231),
.A2(n_219),
.B(n_211),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_35),
.B(n_25),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_188),
.Y(n_258)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_260),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_218),
.Y(n_262)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_238),
.B(n_203),
.C(n_219),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_270),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_214),
.B1(n_219),
.B2(n_152),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_248),
.B1(n_230),
.B2(n_243),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_29),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_42),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_22),
.Y(n_269)
);

AOI32xp33_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_238),
.A3(n_245),
.B1(n_244),
.B2(n_231),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_242),
.B(n_249),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_277),
.B(n_283),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_276),
.B1(n_280),
.B2(n_288),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_258),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_275),
.B(n_254),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_236),
.B1(n_136),
.B2(n_82),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_35),
.B(n_33),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_136),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_279),
.B(n_282),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_257),
.B1(n_271),
.B2(n_261),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_251),
.C(n_252),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_33),
.B(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_257),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_82),
.B1(n_80),
.B2(n_73),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_289),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_299),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_303),
.C(n_305),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_265),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_262),
.B1(n_252),
.B2(n_267),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_288),
.B1(n_276),
.B2(n_274),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_264),
.C(n_253),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_1),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_264),
.C(n_254),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_80),
.C(n_73),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_291),
.C(n_48),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_308),
.B(n_313),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_291),
.B1(n_282),
.B2(n_283),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_310),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_279),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_321),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_296),
.C(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_48),
.C(n_42),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_8),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_293),
.A2(n_298),
.B1(n_306),
.B2(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_20),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_307),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_311),
.A2(n_307),
.B1(n_2),
.B2(n_5),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_324),
.B1(n_326),
.B2(n_310),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_324)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_328),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_8),
.B(n_9),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_29),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_22),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_316),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_315),
.C(n_313),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_337),
.C(n_40),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_40),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_336),
.B(n_340),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_317),
.C(n_22),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_328),
.B(n_10),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_338),
.B(n_11),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_11),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_11),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_326),
.B1(n_12),
.B2(n_13),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_345),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_344),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_347),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_12),
.Y(n_347)
);

AOI31xp33_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_334),
.A3(n_333),
.B(n_14),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_348),
.B(n_13),
.Y(n_353)
);

NAND4xp25_ASAP7_75t_SL g355 ( 
.A(n_353),
.B(n_354),
.C(n_18),
.D(n_13),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_349),
.A2(n_351),
.B(n_350),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_12),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_14),
.C(n_15),
.Y(n_357)
);

OA21x2_ASAP7_75t_SL g358 ( 
.A1(n_357),
.A2(n_15),
.B(n_16),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_18),
.C(n_16),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_359),
.A2(n_17),
.B(n_18),
.Y(n_360)
);


endmodule