module fake_netlist_1_11982_n_715 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_715);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_715;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_704;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_101), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_106), .Y(n_206) );
BUFx10_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_54), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_114), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_91), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_157), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_125), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_103), .B(n_78), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_105), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_113), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_22), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_176), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_141), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_17), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_42), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_143), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_129), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_75), .Y(n_223) );
INVxp33_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_65), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_145), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_118), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_138), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_73), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_89), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_123), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_100), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_79), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_18), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_120), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_13), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_10), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_43), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_117), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_55), .Y(n_241) );
INVxp67_ASAP7_75t_L g242 ( .A(n_202), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_188), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_45), .Y(n_244) );
INVxp33_ASAP7_75t_L g245 ( .A(n_119), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_3), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_165), .Y(n_247) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_111), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_23), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_131), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_160), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_68), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_63), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_164), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_135), .B(n_27), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_47), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_97), .Y(n_257) );
BUFx8_ASAP7_75t_SL g258 ( .A(n_72), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_191), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_64), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_88), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_163), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_3), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_21), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_71), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_27), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_124), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_130), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_77), .Y(n_269) );
INVxp67_ASAP7_75t_SL g270 ( .A(n_70), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_151), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_4), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_87), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_196), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_53), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_128), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_169), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_10), .B(n_74), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_99), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_146), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_24), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_148), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_67), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_98), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_8), .Y(n_286) );
INVxp67_ASAP7_75t_SL g287 ( .A(n_174), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_170), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_33), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_134), .Y(n_290) );
BUFx2_ASAP7_75t_SL g291 ( .A(n_121), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_51), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_76), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_24), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_127), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_20), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_197), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_153), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_108), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_38), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_58), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_102), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_175), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_40), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_22), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_90), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_56), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_21), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_0), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_203), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_66), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_122), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_13), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_11), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_240), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_308), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_240), .Y(n_317) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_248), .B(n_34), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_245), .B(n_0), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_273), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_210), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_241), .B(n_35), .Y(n_323) );
OA21x2_ASAP7_75t_L g324 ( .A1(n_206), .A2(n_37), .B(n_36), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_241), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_245), .B(n_1), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_210), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_275), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_275), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_208), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_277), .B(n_2), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_277), .B(n_4), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_295), .B(n_5), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_298), .B(n_6), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_298), .B(n_6), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_218), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_219), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_216), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_207), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_224), .B(n_7), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_259), .B(n_7), .Y(n_341) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_334), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_319), .Y(n_343) );
AND2x6_ASAP7_75t_L g344 ( .A(n_334), .B(n_209), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_317), .B(n_246), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_339), .Y(n_346) );
NOR2x1p5_ASAP7_75t_L g347 ( .A(n_339), .B(n_294), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_339), .B(n_225), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_341), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_320), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_325), .B(n_264), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_325), .B(n_235), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_334), .B(n_288), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_329), .B(n_266), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_329), .B(n_272), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_315), .B(n_309), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_331), .A2(n_237), .B1(n_249), .B2(n_238), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_326), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_320), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_328), .B(n_225), .Y(n_361) );
INVx3_ASAP7_75t_L g362 ( .A(n_322), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_332), .A2(n_263), .B1(n_286), .B2(n_282), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_348), .B(n_340), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_348), .B(n_340), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_343), .B(n_333), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_346), .B(n_338), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_349), .B(n_333), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_351), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_351), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_362), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_362), .Y(n_372) );
NOR2xp67_ASAP7_75t_L g373 ( .A(n_362), .B(n_322), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_359), .B(n_335), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_342), .Y(n_375) );
OR2x6_ASAP7_75t_L g376 ( .A(n_347), .B(n_335), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_360), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_350), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_342), .B(n_318), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_346), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_361), .B(n_341), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_345), .B(n_205), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_361), .B(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_355), .B(n_330), .Y(n_385) );
AND2x6_ASAP7_75t_SL g386 ( .A(n_356), .B(n_316), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_352), .B(n_336), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_323), .B(n_337), .C(n_336), .Y(n_390) );
BUFx12f_ASAP7_75t_L g391 ( .A(n_386), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_364), .B(n_357), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_388), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_365), .B(n_344), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
NOR2xp33_ASAP7_75t_SL g396 ( .A(n_379), .B(n_256), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_382), .B(n_344), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_387), .A2(n_354), .B1(n_285), .B2(n_300), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_387), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_363), .B(n_358), .C(n_354), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_369), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_375), .B(n_214), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_368), .B(n_374), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_316), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_380), .A2(n_304), .B1(n_313), .B2(n_270), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_367), .A2(n_296), .B(n_289), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_370), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_376), .B(n_305), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_375), .B(n_217), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_390), .A2(n_324), .B(n_270), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_324), .B(n_287), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_376), .B(n_314), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
OAI21x1_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_324), .B(n_299), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_373), .Y(n_419) );
AOI22x1_ASAP7_75t_L g420 ( .A1(n_389), .A2(n_287), .B1(n_223), .B2(n_321), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_376), .B(n_258), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_394), .A2(n_381), .B(n_383), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
AOI21x1_ASAP7_75t_L g424 ( .A1(n_414), .A2(n_324), .B(n_371), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_402), .Y(n_425) );
BUFx10_ASAP7_75t_L g426 ( .A(n_421), .Y(n_426) );
CKINVDCx9p33_ASAP7_75t_R g427 ( .A(n_401), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_406), .B(n_384), .Y(n_428) );
INVx4_ASAP7_75t_L g429 ( .A(n_399), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g430 ( .A1(n_391), .A2(n_244), .B1(n_301), .B2(n_242), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_397), .A2(n_405), .B(n_414), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
O2A1O1Ixp33_ASAP7_75t_SL g433 ( .A1(n_395), .A2(n_372), .B(n_378), .C(n_377), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_413), .A2(n_381), .B(n_244), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_404), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_396), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_212), .B(n_211), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_400), .A2(n_278), .B(n_255), .C(n_215), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_SL g440 ( .A1(n_419), .A2(n_220), .B(n_222), .C(n_221), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_415), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_409), .A2(n_417), .B(n_410), .C(n_407), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_403), .B(n_291), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_420), .B(n_213), .C(n_210), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_418), .A2(n_227), .B(n_226), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_407), .A2(n_229), .B(n_228), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_417), .A2(n_231), .B(n_232), .C(n_230), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_408), .B(n_9), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
AO31x2_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_236), .A3(n_239), .B(n_234), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_247), .B(n_251), .C(n_250), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_441), .A2(n_254), .B1(n_257), .B2(n_252), .Y(n_453) );
OAI21x1_ASAP7_75t_L g454 ( .A1(n_424), .A2(n_303), .B(n_293), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_431), .A2(n_262), .B(n_260), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_437), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_446), .A2(n_268), .B(n_267), .Y(n_457) );
OAI21x1_ASAP7_75t_L g458 ( .A1(n_434), .A2(n_271), .B(n_269), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_442), .B(n_9), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_425), .Y(n_460) );
BUFx6f_ASAP7_75t_SL g461 ( .A(n_426), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_428), .B(n_233), .Y(n_462) );
OR2x6_ASAP7_75t_L g463 ( .A(n_444), .B(n_276), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_433), .A2(n_280), .B(n_279), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_449), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_422), .A2(n_284), .B(n_283), .Y(n_466) );
BUFx8_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_436), .B(n_243), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_450), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_430), .A2(n_307), .B1(n_292), .B2(n_302), .C(n_311), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_438), .A2(n_213), .B(n_297), .C(n_312), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_451), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_443), .A2(n_253), .B(n_210), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_452), .A2(n_253), .B(n_281), .C(n_312), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_448), .A2(n_12), .B(n_14), .C(n_15), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_440), .A2(n_253), .B1(n_281), .B2(n_312), .C(n_310), .Y(n_476) );
OR2x6_ASAP7_75t_L g477 ( .A(n_447), .B(n_12), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_445), .A2(n_327), .B(n_321), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_429), .B(n_14), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_435), .A2(n_327), .B(n_321), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_451), .B(n_16), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_429), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_426), .A2(n_290), .B1(n_265), .B2(n_306), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_432), .B(n_16), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_432), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_444), .B(n_17), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_434), .A2(n_327), .B(n_321), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_423), .B(n_18), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_423), .B(n_19), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g491 ( .A1(n_423), .A2(n_274), .B1(n_261), .B2(n_327), .C1(n_25), .C2(n_26), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_423), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_439), .A2(n_20), .B(n_23), .Y(n_494) );
AOI211xp5_ASAP7_75t_L g495 ( .A1(n_470), .A2(n_25), .B(n_26), .C(n_28), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_465), .B(n_29), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_492), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_494), .A2(n_30), .B(n_31), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_469), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_490), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_482), .B(n_31), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_489), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_493), .Y(n_503) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_473), .A2(n_32), .B(n_33), .Y(n_504) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_488), .A2(n_454), .B(n_472), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_459), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_488), .A2(n_204), .B(n_39), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_481), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_477), .Y(n_510) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_464), .A2(n_41), .B(n_44), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_456), .B(n_46), .Y(n_512) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_478), .A2(n_48), .B(n_49), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_455), .A2(n_50), .B(n_52), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_479), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_467), .Y(n_517) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_458), .A2(n_57), .B(n_59), .Y(n_518) );
AO21x1_ASAP7_75t_SL g519 ( .A1(n_484), .A2(n_60), .B(n_61), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_463), .B(n_62), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_491), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_462), .B(n_69), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_476), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_453), .B(n_80), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_475), .Y(n_526) );
OAI33xp33_ASAP7_75t_L g527 ( .A1(n_468), .A2(n_81), .A3(n_82), .B1(n_83), .B2(n_84), .B3(n_85), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_461), .A2(n_86), .B1(n_92), .B2(n_93), .Y(n_528) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_474), .A2(n_94), .B(n_95), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_471), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_466), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_480), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_483), .B(n_96), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_487), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_477), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_487), .Y(n_537) );
INVx5_ASAP7_75t_L g538 ( .A(n_486), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_487), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_477), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_477), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_487), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_482), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_465), .B(n_104), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_467), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_465), .B(n_107), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_465), .A2(n_109), .B1(n_110), .B2(n_112), .C(n_115), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_499), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_503), .B(n_116), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_535), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_503), .B(n_126), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_537), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_508), .B(n_132), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_536), .A2(n_133), .B1(n_136), .B2(n_137), .Y(n_559) );
NAND2x1p5_ASAP7_75t_SL g560 ( .A(n_549), .B(n_139), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_509), .Y(n_561) );
INVx4_ASAP7_75t_L g562 ( .A(n_538), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_540), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
OR2x6_ASAP7_75t_L g565 ( .A(n_539), .B(n_140), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_544), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_546), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_520), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_547), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_510), .Y(n_571) );
OAI21xp33_ASAP7_75t_SL g572 ( .A1(n_541), .A2(n_142), .B(n_144), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_541), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_514), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_501), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_543), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_542), .B(n_149), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_539), .B(n_150), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_522), .A2(n_152), .B1(n_154), .B2(n_155), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_496), .B(n_156), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_496), .B(n_158), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_545), .B(n_159), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_517), .B(n_161), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_521), .B(n_162), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_545), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_502), .B(n_166), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_500), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_168), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_516), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_538), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_512), .B(n_171), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_522), .B(n_172), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_526), .B(n_173), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_534), .B(n_177), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_498), .B(n_178), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_548), .B(n_179), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_534), .B(n_180), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_495), .A2(n_181), .B(n_182), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_523), .B(n_183), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_534), .B(n_184), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_525), .B(n_185), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_519), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_532), .B(n_186), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_504), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_531), .B(n_189), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_524), .A2(n_190), .B1(n_192), .B2(n_193), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_597), .B(n_518), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_571), .B(n_530), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_555), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_576), .B(n_527), .Y(n_614) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_606), .B(n_528), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_568), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_575), .B(n_574), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_608), .B(n_568), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_554), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_557), .B(n_515), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_570), .B(n_524), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_597), .B(n_507), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_563), .B(n_511), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_566), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_567), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_569), .B(n_533), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_574), .B(n_513), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_552), .B(n_551), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_565), .B(n_529), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_589), .B(n_551), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_564), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_561), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_591), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_591), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_605), .B(n_195), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_577), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_600), .B(n_198), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_594), .B(n_199), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_607), .B(n_200), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_579), .B(n_201), .Y(n_641) );
BUFx2_ASAP7_75t_SL g642 ( .A(n_562), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_609), .B(n_578), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_573), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_580), .B(n_578), .Y(n_645) );
OR2x6_ASAP7_75t_L g646 ( .A(n_637), .B(n_606), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_618), .B(n_592), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_616), .B(n_596), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_618), .B(n_600), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_642), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_617), .B(n_603), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_613), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_632), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_621), .B(n_603), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_624), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_625), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_633), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_634), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_612), .B(n_565), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_614), .A2(n_572), .B(n_559), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_626), .B(n_558), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_626), .B(n_560), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_612), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_638), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_636), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_637), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_620), .B(n_595), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_644), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_643), .B(n_586), .Y(n_670) );
AND2x4_ASAP7_75t_L g671 ( .A(n_620), .B(n_585), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_614), .B(n_583), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_628), .B(n_582), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_648), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_670), .B(n_627), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_664), .B(n_623), .Y(n_676) );
INVx4_ASAP7_75t_L g677 ( .A(n_646), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_653), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_656), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_672), .B(n_645), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_658), .B(n_622), .Y(n_681) );
NAND4xp25_ASAP7_75t_L g682 ( .A(n_661), .B(n_629), .C(n_581), .D(n_622), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_669), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_659), .B(n_630), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_667), .A2(n_637), .B1(n_615), .B2(n_639), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_647), .B(n_631), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_654), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_657), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_678), .Y(n_689) );
NAND4xp25_ASAP7_75t_L g690 ( .A(n_682), .B(n_661), .C(n_651), .D(n_673), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_680), .A2(n_651), .B(n_663), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_684), .B(n_668), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_675), .B(n_671), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_677), .B(n_559), .C(n_601), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_674), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_681), .B(n_665), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_683), .A2(n_646), .B(n_660), .C(n_655), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_690), .B(n_688), .C(n_679), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_689), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_691), .A2(n_676), .B(n_685), .Y(n_700) );
INVx2_ASAP7_75t_SL g701 ( .A(n_693), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g702 ( .A1(n_694), .A2(n_649), .A3(n_650), .B1(n_686), .B2(n_652), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_692), .B1(n_696), .B2(n_697), .C(n_695), .Y(n_703) );
NOR3xp33_ASAP7_75t_L g704 ( .A(n_698), .B(n_610), .C(n_640), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g705 ( .A(n_704), .B(n_700), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_703), .B(n_699), .C(n_598), .Y(n_706) );
OAI211xp5_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_701), .B(n_641), .C(n_604), .Y(n_707) );
NAND5xp2_ASAP7_75t_L g708 ( .A(n_705), .B(n_611), .C(n_602), .D(n_593), .E(n_599), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_707), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_709), .B(n_708), .Y(n_710) );
AO22x2_ASAP7_75t_L g711 ( .A1(n_710), .A2(n_584), .B1(n_590), .B2(n_588), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_590), .B(n_588), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_712), .A2(n_687), .B1(n_666), .B2(n_662), .Y(n_713) );
OAI31xp33_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_553), .A3(n_556), .B(n_635), .Y(n_714) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_553), .B(n_556), .Y(n_715) );
endmodule