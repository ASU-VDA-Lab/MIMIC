module fake_jpeg_7285_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_33),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_30),
.B1(n_20),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_49),
.B1(n_59),
.B2(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_51),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g57 ( 
.A1(n_34),
.A2(n_25),
.B(n_26),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_20),
.B2(n_24),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_22),
.C(n_31),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_27),
.B(n_18),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_35),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_27),
.B1(n_18),
.B2(n_17),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_79),
.B1(n_87),
.B2(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_17),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_0),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_16),
.B1(n_29),
.B2(n_21),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_85),
.B1(n_89),
.B2(n_44),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_78),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_32),
.B1(n_26),
.B2(n_29),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_90),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_54),
.B1(n_66),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_26),
.B1(n_29),
.B2(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_25),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_93),
.B(n_109),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_69),
.B(n_16),
.C(n_21),
.Y(n_129)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_55),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_58),
.B1(n_51),
.B2(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_53),
.B1(n_62),
.B2(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_62),
.B1(n_44),
.B2(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_73),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_19),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_19),
.C(n_21),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_110),
.Y(n_116)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_84),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_120),
.B(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_123),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_88),
.B1(n_82),
.B2(n_89),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_76),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_74),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_129),
.B1(n_23),
.B2(n_48),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_69),
.B1(n_16),
.B2(n_29),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_101),
.B1(n_113),
.B2(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_114),
.B1(n_95),
.B2(n_91),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_23),
.B1(n_44),
.B2(n_3),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_138),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_103),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_19),
.C(n_23),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_112),
.C(n_107),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_144),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_147),
.C(n_156),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_135),
.B1(n_129),
.B2(n_137),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_109),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_96),
.C(n_25),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_0),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_139),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_23),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_130),
.C(n_136),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_141),
.C(n_147),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_23),
.B1(n_1),
.B2(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_2),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_168),
.B(n_177),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_155),
.B1(n_154),
.B2(n_156),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_133),
.B1(n_139),
.B2(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_185),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_140),
.B(n_144),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_138),
.C(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_116),
.B1(n_23),
.B2(n_4),
.Y(n_186)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_2),
.C(n_3),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_188),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_149),
.B1(n_146),
.B2(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_192),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_205),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_177),
.B1(n_186),
.B2(n_153),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_157),
.B(n_158),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_173),
.B(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_180),
.B1(n_178),
.B2(n_169),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_143),
.C(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_207),
.C(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_163),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_199),
.A2(n_175),
.B1(n_179),
.B2(n_185),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_220),
.B1(n_207),
.B2(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_219),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_224),
.B(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_170),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_182),
.B1(n_164),
.B2(n_183),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_204),
.C(n_193),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_167),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_210),
.B(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_224),
.B1(n_205),
.B2(n_218),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_202),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_234),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_187),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_196),
.B(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_200),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_238),
.B(n_159),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_231),
.B1(n_200),
.B2(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_245),
.B1(n_212),
.B2(n_221),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_246),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_214),
.C(n_224),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_230),
.CI(n_235),
.CON(n_248),
.SN(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_253),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_249),
.A2(n_251),
.A3(n_255),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_229),
.B1(n_182),
.B2(n_176),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_239),
.B1(n_214),
.B2(n_240),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_234),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_153),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_214),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_247),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_248),
.B1(n_254),
.B2(n_250),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_153),
.B1(n_4),
.B2(n_5),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_7),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_2),
.C(n_4),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_260),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_12),
.B(n_13),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_256),
.C(n_258),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_9),
.B(n_12),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_263),
.B(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_13),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_270),
.C(n_13),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_14),
.Y(n_274)
);


endmodule