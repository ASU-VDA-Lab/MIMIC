module fake_netlist_6_4645_n_1659 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1659);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1659;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx3_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_94),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_45),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_25),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_78),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_36),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_48),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_101),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_34),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_98),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_25),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_26),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_12),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_112),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_108),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_65),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_51),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_104),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_99),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_162),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_57),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_46),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_142),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_31),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_74),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_45),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_53),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_83),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_49),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_52),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_82),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_106),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_95),
.Y(n_240)
);

BUFx2_ASAP7_75t_SL g241 ( 
.A(n_69),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_123),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_20),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_87),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_40),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_26),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_39),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_39),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_169),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_5),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_72),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_42),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_167),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_44),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_75),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_97),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_144),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_103),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_124),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_165),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_132),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_54),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_56),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_48),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_35),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_88),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_85),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_161),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_159),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_44),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_121),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_17),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_150),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_13),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_68),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_130),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_62),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_59),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_126),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_76),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_89),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_84),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_146),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_114),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_16),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_4),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_129),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_110),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_149),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_28),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_22),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_58),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_32),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_100),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_29),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_81),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_19),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_16),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_51),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_1),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_40),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_154),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_29),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_18),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_140),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_30),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_32),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_7),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_66),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_160),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_0),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_42),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_151),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_90),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_122),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_158),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_14),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_11),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_221),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_227),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_242),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_240),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_222),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_213),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_180),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_247),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_260),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_180),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_180),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_0),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_177),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_223),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_180),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_178),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_208),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_180),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_224),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_180),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_226),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_229),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_180),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_238),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_243),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_272),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_246),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_172),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_L g378 ( 
.A(n_216),
.B(n_2),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_172),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_311),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_264),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_191),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_328),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_175),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_191),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_266),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_268),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_270),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_239),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_239),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_271),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_249),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_249),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_286),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_286),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_322),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_315),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_255),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_216),
.B(n_3),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_206),
.B(n_4),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_225),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_206),
.B(n_5),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_298),
.B(n_6),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_184),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_186),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_228),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_R g414 ( 
.A(n_173),
.B(n_109),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_204),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_218),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_298),
.B(n_7),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_236),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_173),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_196),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_174),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_174),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_251),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_265),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_230),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_276),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_231),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_196),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_382),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_215),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_215),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_343),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_348),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_358),
.B(n_176),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_347),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_363),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_365),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_366),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_351),
.A2(n_357),
.B1(n_382),
.B2(n_345),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

AND3x2_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_304),
.C(n_269),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_377),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_368),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_352),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_350),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_371),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_385),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_419),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_370),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_373),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_376),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_346),
.A2(n_263),
.B1(n_261),
.B2(n_253),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_350),
.B(n_219),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_384),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_421),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_383),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_R g468 ( 
.A(n_406),
.B(n_179),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_422),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_388),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_354),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_389),
.B(n_219),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_393),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_402),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_400),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_354),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_279),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_410),
.Y(n_483)
);

NAND2xp33_ASAP7_75t_SL g484 ( 
.A(n_360),
.B(n_186),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_416),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_361),
.B(n_269),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_410),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_425),
.B(n_427),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_386),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_361),
.B(n_304),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_355),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_405),
.B(n_309),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_407),
.B(n_309),
.Y(n_494)
);

BUFx8_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_355),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_359),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_378),
.B(n_404),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_359),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_362),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_349),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_464),
.B(n_279),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_428),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_480),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_464),
.B(n_362),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_464),
.B(n_364),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_488),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_409),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_468),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_353),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_279),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_481),
.A2(n_330),
.B1(n_290),
.B2(n_308),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_429),
.B(n_279),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_429),
.B(n_279),
.Y(n_524)
);

BUFx4f_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_432),
.B(n_367),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_432),
.B(n_181),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_436),
.B(n_486),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_447),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_491),
.A2(n_190),
.B1(n_281),
.B2(n_340),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_434),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_473),
.B(n_182),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_433),
.B(n_426),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_492),
.B(n_367),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_451),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_433),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_369),
.Y(n_539)
);

CKINVDCx14_ASAP7_75t_R g540 ( 
.A(n_435),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_411),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_463),
.B(n_443),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_209),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_451),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_440),
.B(n_195),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_500),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_471),
.B(n_443),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_498),
.B(n_444),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_369),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_481),
.B(n_185),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_443),
.B(n_189),
.Y(n_554)
);

BUFx8_ASAP7_75t_SL g555 ( 
.A(n_439),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_446),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_456),
.B(n_194),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_472),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_465),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_459),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_442),
.B(n_426),
.Y(n_564)
);

CKINVDCx6p67_ASAP7_75t_R g565 ( 
.A(n_430),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_448),
.B(n_415),
.Y(n_566)
);

BUFx10_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_497),
.B(n_183),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_461),
.B(n_462),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_465),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_485),
.B(n_415),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_467),
.B(n_198),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_459),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_465),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_499),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_482),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_445),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_424),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_445),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_431),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_485),
.B(n_438),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_484),
.B(n_273),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_485),
.B(n_241),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_450),
.B(n_200),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_478),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_482),
.B(n_418),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_437),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_437),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_490),
.A2(n_307),
.B1(n_319),
.B2(n_321),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_466),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_445),
.B(n_424),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_495),
.B(n_202),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_495),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_476),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_476),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

INVxp33_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_495),
.A2(n_179),
.B1(n_281),
.B2(n_340),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_455),
.B(n_285),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_477),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_477),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_479),
.B(n_212),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_479),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

CKINVDCx14_ASAP7_75t_R g610 ( 
.A(n_458),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_466),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_469),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_464),
.B(n_423),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_464),
.B(n_217),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_464),
.B(n_220),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_493),
.A2(n_317),
.B1(n_320),
.B2(n_325),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_493),
.A2(n_341),
.B1(n_423),
.B2(n_256),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_464),
.B(n_232),
.Y(n_620)
);

INVx4_ASAP7_75t_SL g621 ( 
.A(n_428),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_235),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_454),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_464),
.B(n_237),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_489),
.A2(n_293),
.B1(n_292),
.B2(n_291),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_493),
.B(n_245),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_454),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_428),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_428),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_444),
.A2(n_257),
.B1(n_342),
.B2(n_335),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_493),
.A2(n_334),
.B1(n_295),
.B2(n_299),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_433),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_234),
.C(n_326),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_464),
.B(n_248),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_428),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_449),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_459),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_454),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g640 ( 
.A(n_433),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_510),
.B(n_258),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_550),
.A2(n_293),
.B1(n_274),
.B2(n_259),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_277),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_525),
.B(n_262),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_526),
.B(n_267),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_525),
.B(n_414),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_632),
.B(n_327),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_547),
.B(n_278),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_555),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_622),
.A2(n_312),
.B1(n_282),
.B2(n_289),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_505),
.B(n_294),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_614),
.B(n_337),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_632),
.B(n_187),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_614),
.B(n_187),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_545),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_207),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_506),
.B(n_190),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_518),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_640),
.B(n_193),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_640),
.B(n_529),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_639),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_517),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_529),
.B(n_193),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_552),
.B(n_197),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_550),
.A2(n_300),
.B1(n_214),
.B2(n_211),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_552),
.B(n_197),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_583),
.B(n_188),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_566),
.B(n_207),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_519),
.A2(n_301),
.B1(n_214),
.B2(n_211),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_538),
.B(n_199),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_518),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_622),
.A2(n_205),
.B1(n_188),
.B2(n_192),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_507),
.B(n_199),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_531),
.B(n_201),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_511),
.B(n_201),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_535),
.B(n_203),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_622),
.B(n_259),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_622),
.B(n_522),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_542),
.A2(n_300),
.B1(n_339),
.B2(n_338),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_542),
.A2(n_306),
.B1(n_314),
.B2(n_305),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_622),
.B(n_274),
.Y(n_684)
);

AND2x4_ASAP7_75t_SL g685 ( 
.A(n_556),
.B(n_311),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_522),
.B(n_284),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_533),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_615),
.B(n_284),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_631),
.A2(n_333),
.B(n_287),
.C(n_291),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_631),
.A2(n_205),
.B1(n_336),
.B2(n_332),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_537),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_524),
.B(n_287),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_537),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_524),
.B(n_292),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_582),
.A2(n_314),
.B(n_297),
.Y(n_696)
);

BUFx2_ASAP7_75t_L g697 ( 
.A(n_609),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_527),
.A2(n_305),
.B1(n_339),
.B2(n_333),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_501),
.B(n_207),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_626),
.B(n_233),
.C(n_244),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_618),
.A2(n_192),
.B1(n_210),
.B2(n_275),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_568),
.B(n_297),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_544),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_513),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_623),
.B(n_301),
.Y(n_705)
);

AO221x1_ASAP7_75t_L g706 ( 
.A1(n_592),
.A2(n_311),
.B1(n_399),
.B2(n_397),
.C(n_396),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_593),
.B(n_210),
.Y(n_707)
);

AOI221xp5_ASAP7_75t_L g708 ( 
.A1(n_618),
.A2(n_332),
.B1(n_275),
.B2(n_280),
.C(n_283),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_508),
.B(n_306),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_543),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_516),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_634),
.B(n_338),
.Y(n_712)
);

INVx8_ASAP7_75t_L g713 ( 
.A(n_584),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_620),
.B(n_250),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_541),
.B(n_401),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_584),
.A2(n_252),
.B1(n_323),
.B2(n_283),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_516),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_609),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_555),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_586),
.B(n_401),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_521),
.B(n_399),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_625),
.B(n_280),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_573),
.B(n_288),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_624),
.B(n_288),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_586),
.B(n_397),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_521),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_635),
.B(n_302),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_627),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_551),
.B(n_536),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_581),
.B(n_396),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_539),
.B(n_553),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_573),
.B(n_302),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_512),
.B(n_303),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_619),
.A2(n_303),
.B1(n_313),
.B2(n_331),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_619),
.A2(n_313),
.B1(n_331),
.B2(n_336),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_595),
.B(n_575),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_534),
.B(n_8),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_616),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_549),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_594),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_572),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_534),
.B(n_8),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_571),
.B(n_395),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_577),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_569),
.B(n_67),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_527),
.B(n_9),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_577),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_503),
.A2(n_394),
.B(n_392),
.C(n_391),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_515),
.A2(n_392),
.B1(n_391),
.B2(n_387),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_557),
.B(n_617),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_633),
.Y(n_751)
);

BUFx8_ASAP7_75t_L g752 ( 
.A(n_608),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_554),
.B(n_9),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_560),
.B(n_387),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_561),
.B(n_55),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_554),
.B(n_10),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_626),
.A2(n_170),
.B1(n_157),
.B2(n_152),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_637),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_617),
.B(n_10),
.Y(n_759)
);

OAI22xp33_ASAP7_75t_L g760 ( 
.A1(n_584),
.A2(n_548),
.B1(n_603),
.B2(n_604),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_576),
.B(n_139),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_588),
.B(n_562),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_588),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_138),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_567),
.B(n_14),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_575),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_559),
.B(n_136),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_559),
.B(n_504),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_515),
.B(n_127),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_607),
.B(n_19),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_520),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_558),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_558),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_585),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_504),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_604),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_604),
.Y(n_777)
);

INVx8_ASAP7_75t_L g778 ( 
.A(n_595),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_509),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_548),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_607),
.A2(n_115),
.B1(n_113),
.B2(n_111),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_520),
.A2(n_107),
.B1(n_105),
.B2(n_96),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_630),
.A2(n_24),
.B1(n_27),
.B2(n_34),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_509),
.B(n_530),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_556),
.B(n_27),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_530),
.B(n_93),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_569),
.B(n_548),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_570),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_643),
.B(n_763),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_643),
.A2(n_606),
.B(n_605),
.C(n_540),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_762),
.A2(n_528),
.B(n_570),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_590),
.Y(n_793)
);

AO32x1_ASAP7_75t_L g794 ( 
.A1(n_783),
.A2(n_766),
.A3(n_772),
.B1(n_773),
.B2(n_751),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_681),
.A2(n_580),
.B(n_598),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_731),
.A2(n_599),
.B(n_580),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_720),
.B(n_595),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_725),
.B(n_595),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_740),
.B(n_595),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_645),
.A2(n_599),
.B(n_608),
.C(n_597),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_737),
.A2(n_613),
.B(n_612),
.C(n_638),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_662),
.B(n_629),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_658),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

AO21x2_ASAP7_75t_L g805 ( 
.A1(n_645),
.A2(n_621),
.B(n_629),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_731),
.A2(n_580),
.B(n_621),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_726),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_662),
.B(n_628),
.Y(n_808)
);

BUFx4f_ASAP7_75t_L g809 ( 
.A(n_718),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_715),
.B(n_628),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_744),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_697),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_785),
.A2(n_580),
.B(n_621),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_670),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_726),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_747),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_784),
.A2(n_532),
.B1(n_591),
.B2(n_602),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_665),
.A2(n_567),
.B1(n_565),
.B2(n_611),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_732),
.A2(n_737),
.B(n_742),
.C(n_770),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_665),
.B(n_636),
.Y(n_820)
);

OR2x6_ASAP7_75t_SL g821 ( 
.A(n_669),
.B(n_610),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_742),
.A2(n_610),
.B(n_602),
.C(n_574),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_778),
.B(n_546),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_657),
.B(n_589),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_726),
.Y(n_826)
);

AOI21x1_ASAP7_75t_L g827 ( 
.A1(n_646),
.A2(n_502),
.B(n_600),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_719),
.B(n_92),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_666),
.A2(n_502),
.B(n_563),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_654),
.A2(n_736),
.B(n_652),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_711),
.B(n_574),
.Y(n_831)
);

INVx11_ASAP7_75t_L g832 ( 
.A(n_752),
.Y(n_832)
);

INVx11_ASAP7_75t_L g833 ( 
.A(n_704),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_648),
.B(n_655),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_717),
.B(n_563),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_784),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_SL g837 ( 
.A1(n_769),
.A2(n_41),
.B(n_46),
.C(n_50),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_647),
.A2(n_676),
.B(n_767),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_770),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_699),
.B(n_54),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_63),
.B1(n_601),
.B2(n_750),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_655),
.B(n_601),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_661),
.B(n_743),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_651),
.B1(n_677),
.B2(n_756),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_788),
.A2(n_712),
.B1(n_668),
.B2(n_677),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_726),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_768),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_777),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_707),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_702),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_789),
.A2(n_781),
.B(n_787),
.Y(n_851)
);

OAI21xp33_ASAP7_75t_L g852 ( 
.A1(n_691),
.A2(n_735),
.B(n_734),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_746),
.A2(n_753),
.B(n_756),
.C(n_759),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_660),
.Y(n_854)
);

AND2x6_ASAP7_75t_L g855 ( 
.A(n_753),
.B(n_746),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_759),
.A2(n_712),
.B(n_642),
.C(n_667),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_675),
.B(n_682),
.C(n_683),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_775),
.A2(n_779),
.B(n_692),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_748),
.A2(n_690),
.B(n_741),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_679),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_674),
.A2(n_687),
.B(n_694),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_663),
.A2(n_728),
.B1(n_664),
.B2(n_688),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_721),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_738),
.B(n_760),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_686),
.A2(n_693),
.B(n_695),
.C(n_745),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_703),
.A2(n_758),
.B(n_739),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_650),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_659),
.B(n_649),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_656),
.B(n_738),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_776),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_684),
.A2(n_689),
.B1(n_714),
.B2(n_760),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_672),
.A2(n_764),
.B(n_768),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_755),
.A2(n_761),
.B(n_705),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_755),
.A2(n_761),
.B(n_778),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_754),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_738),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_714),
.B(n_733),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_L g878 ( 
.A1(n_691),
.A2(n_734),
.B(n_735),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_724),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_680),
.A2(n_651),
.B(n_724),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_727),
.A2(n_696),
.B(n_678),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_718),
.B(n_777),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_727),
.A2(n_713),
.B(n_709),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_771),
.A2(n_722),
.B(n_723),
.C(n_780),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_713),
.A2(n_782),
.B(n_749),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_780),
.A2(n_765),
.B(n_786),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_718),
.B(n_700),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_713),
.B(n_716),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_671),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_698),
.B(n_749),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_757),
.A2(n_706),
.B(n_685),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_708),
.A2(n_701),
.B(n_710),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_701),
.A2(n_729),
.B(n_681),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_662),
.B(n_525),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_729),
.A2(n_525),
.B(n_762),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_731),
.A2(n_729),
.B(n_526),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_643),
.B(n_699),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_774),
.B(n_643),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_641),
.B(n_595),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_643),
.A2(n_510),
.B(n_732),
.C(n_662),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_774),
.B(n_643),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_729),
.A2(n_525),
.B(n_762),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_731),
.A2(n_729),
.B(n_526),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_643),
.B(n_673),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_774),
.B(n_643),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_729),
.A2(n_525),
.B(n_762),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_643),
.B(n_732),
.C(n_677),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_774),
.B(n_643),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_774),
.B(n_643),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_643),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_729),
.A2(n_525),
.B(n_762),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_657),
.B(n_508),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_774),
.B(n_643),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_697),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_774),
.B(n_643),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_641),
.A2(n_770),
.B(n_756),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_774),
.B(n_643),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_744),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_L g919 ( 
.A(n_643),
.B(n_430),
.C(n_630),
.Y(n_919)
);

BUFx12f_ASAP7_75t_L g920 ( 
.A(n_752),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_643),
.B(n_673),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_752),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_711),
.B(n_717),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_774),
.B(n_643),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_770),
.A2(n_643),
.B1(n_677),
.B2(n_737),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_662),
.B(n_525),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_774),
.B(n_643),
.Y(n_927)
);

OAI321xp33_ASAP7_75t_L g928 ( 
.A1(n_784),
.A2(n_643),
.A3(n_770),
.B1(n_641),
.B2(n_780),
.C(n_510),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_643),
.B(n_673),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_662),
.A2(n_643),
.B1(n_774),
.B2(n_510),
.Y(n_930)
);

OAI22x1_ASAP7_75t_L g931 ( 
.A1(n_643),
.A2(n_543),
.B1(n_770),
.B2(n_591),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_643),
.B(n_732),
.C(n_677),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_643),
.A2(n_510),
.B(n_732),
.C(n_662),
.Y(n_933)
);

AOI21x1_ASAP7_75t_L g934 ( 
.A1(n_731),
.A2(n_729),
.B(n_526),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_643),
.A2(n_732),
.B(n_691),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_729),
.A2(n_681),
.B(n_641),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_653),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_650),
.Y(n_938)
);

A2O1A1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_643),
.A2(n_510),
.B(n_732),
.C(n_662),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_914),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_830),
.A2(n_823),
.B(n_895),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_897),
.B(n_904),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_812),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_853),
.A2(n_844),
.B(n_900),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_831),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_898),
.B(n_901),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_L g947 ( 
.A(n_855),
.B(n_856),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_851),
.A2(n_796),
.B(n_806),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_930),
.B(n_845),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_933),
.B(n_939),
.Y(n_950)
);

BUFx8_ASAP7_75t_SL g951 ( 
.A(n_938),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_804),
.B(n_920),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_905),
.B(n_908),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_909),
.B(n_910),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_813),
.A2(n_903),
.B(n_896),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_844),
.A2(n_878),
.B1(n_852),
.B2(n_857),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_825),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_934),
.A2(n_858),
.B(n_792),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_831),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_842),
.A2(n_926),
.B(n_894),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_884),
.A2(n_834),
.B(n_928),
.C(n_880),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_807),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_911),
.B(n_906),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_843),
.B(n_790),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_913),
.B(n_915),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_916),
.A2(n_795),
.B(n_936),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_928),
.A2(n_892),
.B(n_893),
.C(n_924),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_936),
.B(n_893),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_807),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_917),
.B(n_927),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_849),
.B(n_860),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_867),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_921),
.A2(n_929),
.B(n_850),
.Y(n_973)
);

OAI21x1_ASAP7_75t_SL g974 ( 
.A1(n_881),
.A2(n_886),
.B(n_885),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_807),
.Y(n_975)
);

AO31x2_ASAP7_75t_L g976 ( 
.A1(n_865),
.A2(n_802),
.A3(n_808),
.B(n_873),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_849),
.B(n_860),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_912),
.B(n_815),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_820),
.A2(n_827),
.B(n_872),
.Y(n_979)
);

AO31x2_ASAP7_75t_L g980 ( 
.A1(n_793),
.A2(n_838),
.A3(n_891),
.B(n_874),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_815),
.B(n_826),
.Y(n_981)
);

AOI221x1_ASAP7_75t_L g982 ( 
.A1(n_919),
.A2(n_829),
.B1(n_931),
.B2(n_836),
.C(n_791),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_855),
.B(n_875),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_800),
.A2(n_866),
.B(n_861),
.Y(n_984)
);

NAND2x1_ASAP7_75t_L g985 ( 
.A(n_826),
.B(n_811),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_855),
.B(n_868),
.Y(n_986)
);

OAI21x1_ASAP7_75t_SL g987 ( 
.A1(n_877),
.A2(n_883),
.B(n_836),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_859),
.A2(n_890),
.B(n_855),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_846),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_810),
.A2(n_869),
.B(n_899),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_846),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_889),
.B(n_879),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_876),
.B(n_847),
.Y(n_993)
);

NAND3xp33_ASAP7_75t_L g994 ( 
.A(n_803),
.B(n_814),
.C(n_801),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_816),
.B(n_918),
.Y(n_995)
);

OA21x2_ASAP7_75t_L g996 ( 
.A1(n_829),
.A2(n_871),
.B(n_864),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_841),
.A2(n_862),
.B1(n_839),
.B2(n_840),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_923),
.B(n_863),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_816),
.A2(n_847),
.B(n_805),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_937),
.B(n_846),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_923),
.B(n_817),
.Y(n_1001)
);

NAND2x1_ASAP7_75t_L g1002 ( 
.A(n_887),
.B(n_882),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_870),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_828),
.A2(n_888),
.B(n_794),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_848),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_882),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_835),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_812),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_824),
.B(n_818),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_SL g1010 ( 
.A1(n_822),
.A2(n_817),
.B(n_837),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_809),
.B(n_835),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_794),
.A2(n_833),
.B(n_821),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_832),
.B(n_922),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_907),
.B(n_932),
.Y(n_1014)
);

BUFx4_ASAP7_75t_SL g1015 ( 
.A(n_938),
.Y(n_1015)
);

AOI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_852),
.A2(n_878),
.B1(n_935),
.B2(n_643),
.C(n_932),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_900),
.B(n_939),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_830),
.A2(n_525),
.B(n_823),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_907),
.A2(n_932),
.B1(n_819),
.B2(n_853),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_916),
.A2(n_853),
.A3(n_819),
.B(n_844),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_898),
.B(n_901),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_930),
.B(n_898),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_812),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_907),
.A2(n_932),
.B(n_935),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_830),
.A2(n_525),
.B(n_823),
.Y(n_1025)
);

AO31x2_ASAP7_75t_L g1026 ( 
.A1(n_916),
.A2(n_853),
.A3(n_819),
.B(n_844),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_812),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_854),
.Y(n_1028)
);

AO32x2_ASAP7_75t_L g1029 ( 
.A1(n_844),
.A2(n_836),
.A3(n_839),
.B1(n_928),
.B2(n_916),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_897),
.B(n_904),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_900),
.B(n_939),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_812),
.Y(n_1032)
);

AOI21x1_ASAP7_75t_SL g1033 ( 
.A1(n_797),
.A2(n_798),
.B(n_799),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_854),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_901),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_900),
.B(n_939),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_923),
.B(n_711),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_925),
.A2(n_819),
.B(n_933),
.C(n_900),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_854),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_930),
.B(n_898),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_907),
.B(n_932),
.C(n_935),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_804),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_930),
.B(n_898),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_795),
.A2(n_936),
.B(n_893),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_SL g1049 ( 
.A1(n_907),
.A2(n_932),
.B1(n_643),
.B2(n_844),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_851),
.A2(n_796),
.B(n_806),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_938),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_854),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_851),
.A2(n_796),
.B(n_806),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_897),
.B(n_904),
.Y(n_1055)
);

O2A1O1Ixp5_ASAP7_75t_L g1056 ( 
.A1(n_925),
.A2(n_819),
.B(n_933),
.C(n_900),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_819),
.A2(n_853),
.B(n_844),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_907),
.A2(n_932),
.B1(n_819),
.B2(n_853),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_851),
.A2(n_796),
.B(n_806),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_812),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_SL g1061 ( 
.A(n_835),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1032),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_943),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_977),
.B(n_1023),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_953),
.B(n_964),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_962),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_971),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_964),
.B(n_970),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_957),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_969),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_1051),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1049),
.A2(n_949),
.B1(n_1044),
.B2(n_1052),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_941),
.A2(n_947),
.B(n_963),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_970),
.B(n_946),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_1008),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_1046),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1022),
.B(n_1042),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1047),
.B(n_954),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_965),
.B(n_1021),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_940),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_990),
.A2(n_961),
.B(n_988),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_951),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1036),
.B(n_942),
.Y(n_1083)
);

AND2x2_ASAP7_75t_SL g1084 ( 
.A(n_1016),
.B(n_996),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_1023),
.B(n_1027),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1030),
.B(n_1055),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1027),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1006),
.B(n_998),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1060),
.Y(n_1089)
);

AOI221x1_ASAP7_75t_L g1090 ( 
.A1(n_1035),
.A2(n_1045),
.B1(n_1041),
.B2(n_1057),
.C(n_1052),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_973),
.B(n_992),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1060),
.B(n_998),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1035),
.A2(n_1057),
.B1(n_1045),
.B2(n_1043),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1041),
.A2(n_1043),
.B1(n_944),
.B2(n_1058),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_944),
.A2(n_1039),
.B(n_1056),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1024),
.A2(n_967),
.B(n_1058),
.C(n_1019),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1005),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1038),
.B(n_1007),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_945),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_972),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1015),
.Y(n_1101)
);

INVxp67_ASAP7_75t_L g1102 ( 
.A(n_959),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_952),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_950),
.A2(n_1037),
.B(n_1031),
.Y(n_1104)
);

OR2x6_ASAP7_75t_SL g1105 ( 
.A(n_1019),
.B(n_997),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1014),
.B(n_1001),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_986),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_986),
.Y(n_1108)
);

AOI21xp33_ASAP7_75t_L g1109 ( 
.A1(n_956),
.A2(n_1017),
.B(n_997),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1002),
.B(n_1011),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_956),
.B(n_982),
.C(n_994),
.Y(n_1111)
);

AND2x4_ASAP7_75t_SL g1112 ( 
.A(n_1038),
.B(n_1013),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_1007),
.B(n_978),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_969),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1000),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_962),
.Y(n_1116)
);

INVx6_ASAP7_75t_SL g1117 ( 
.A(n_952),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_955),
.A2(n_958),
.B(n_974),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_983),
.B(n_1053),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_1000),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_983),
.B(n_1003),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1028),
.B(n_1034),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_996),
.B(n_1020),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1010),
.A2(n_987),
.B1(n_1040),
.B2(n_1061),
.Y(n_1124)
);

INVx5_ASAP7_75t_L g1125 ( 
.A(n_962),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_993),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_991),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1020),
.B(n_1026),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_991),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1013),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_1004),
.B(n_1061),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_989),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1029),
.A2(n_1048),
.B1(n_968),
.B2(n_969),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1012),
.B(n_1020),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_952),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1136)
);

INVx3_ASAP7_75t_SL g1137 ( 
.A(n_975),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_981),
.B(n_985),
.Y(n_1138)
);

CKINVDCx11_ASAP7_75t_R g1139 ( 
.A(n_1026),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_966),
.B(n_968),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_976),
.B(n_995),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_976),
.B(n_960),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_999),
.B(n_980),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_979),
.B(n_948),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_984),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1029),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1050),
.A2(n_1054),
.B(n_1059),
.C(n_1033),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_964),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_980),
.A2(n_1025),
.B(n_1018),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1049),
.A2(n_907),
.B1(n_932),
.B2(n_819),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1032),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1006),
.B(n_998),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1006),
.B(n_998),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1049),
.A2(n_907),
.B1(n_932),
.B2(n_819),
.Y(n_1154)
);

AOI221x1_ASAP7_75t_L g1155 ( 
.A1(n_1035),
.A2(n_1041),
.B1(n_1052),
.B2(n_1045),
.C(n_1043),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_SL g1156 ( 
.A1(n_1009),
.A2(n_932),
.B1(n_907),
.B2(n_786),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1006),
.B(n_998),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_943),
.B(n_907),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1006),
.B(n_998),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_953),
.B(n_964),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_971),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_943),
.B(n_907),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1023),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_1049),
.B(n_932),
.C(n_907),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1049),
.B(n_932),
.C(n_907),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_951),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_953),
.B(n_964),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_942),
.B(n_1030),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_SL g1169 ( 
.A1(n_944),
.A2(n_643),
.B(n_1057),
.C(n_1052),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1032),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_942),
.B(n_1030),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_1046),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1016),
.A2(n_907),
.B(n_932),
.C(n_935),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1049),
.A2(n_907),
.B1(n_932),
.B2(n_819),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_969),
.B(n_815),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_962),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_957),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_1051),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_943),
.B(n_907),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_943),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_SL g1181 ( 
.A1(n_961),
.A2(n_853),
.B(n_819),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_962),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_969),
.B(n_815),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_957),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_971),
.B(n_946),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1019),
.A2(n_1058),
.B(n_956),
.Y(n_1186)
);

CKINVDCx8_ASAP7_75t_R g1187 ( 
.A(n_972),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1149),
.A2(n_1073),
.B(n_1081),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1086),
.B(n_1168),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1164),
.A2(n_1165),
.B(n_1173),
.Y(n_1190)
);

BUFx4_ASAP7_75t_SL g1191 ( 
.A(n_1100),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1072),
.A2(n_1150),
.B1(n_1154),
.B2(n_1174),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1077),
.B(n_1078),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1119),
.Y(n_1194)
);

BUFx8_ASAP7_75t_L g1195 ( 
.A(n_1076),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1065),
.A2(n_1160),
.B1(n_1167),
.B2(n_1068),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_1082),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1110),
.B(n_1126),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1116),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1164),
.A2(n_1165),
.B1(n_1094),
.B2(n_1093),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1186),
.A2(n_1156),
.B1(n_1109),
.B2(n_1111),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1077),
.B(n_1083),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1107),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1107),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1177),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1184),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1110),
.B(n_1098),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1074),
.A2(n_1078),
.B1(n_1079),
.B2(n_1106),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1112),
.Y(n_1209)
);

CKINVDCx14_ASAP7_75t_R g1210 ( 
.A(n_1178),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1108),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1070),
.B(n_1114),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1122),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1147),
.A2(n_1169),
.B(n_1095),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1115),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1098),
.B(n_1088),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1109),
.A2(n_1111),
.B1(n_1095),
.B2(n_1091),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1120),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1079),
.B(n_1171),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1158),
.A2(n_1162),
.B1(n_1179),
.B2(n_1088),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1070),
.B(n_1114),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1118),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1090),
.A2(n_1155),
.B(n_1142),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_1157),
.B2(n_1159),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1105),
.A2(n_1185),
.B1(n_1161),
.B2(n_1067),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1145),
.A2(n_1141),
.B(n_1144),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1166),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1132),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1089),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1163),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1087),
.A2(n_1062),
.B1(n_1151),
.B2(n_1170),
.Y(n_1231)
);

CKINVDCx6p67_ASAP7_75t_R g1232 ( 
.A(n_1172),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1116),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1092),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1121),
.Y(n_1235)
);

AO21x1_ASAP7_75t_SL g1236 ( 
.A1(n_1148),
.A2(n_1128),
.B(n_1146),
.Y(n_1236)
);

BUFx12f_ASAP7_75t_L g1237 ( 
.A(n_1135),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1064),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1075),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1133),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1123),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1084),
.Y(n_1242)
);

NAND2x1p5_ASAP7_75t_L g1243 ( 
.A(n_1125),
.B(n_1113),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1085),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1071),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1096),
.A2(n_1140),
.B(n_1128),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1124),
.A2(n_1097),
.B1(n_1181),
.B2(n_1102),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1097),
.A2(n_1099),
.B1(n_1180),
.B2(n_1063),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1127),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1139),
.A2(n_1104),
.B1(n_1117),
.B2(n_1134),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1131),
.A2(n_1101),
.B1(n_1103),
.B2(n_1113),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1080),
.Y(n_1252)
);

CKINVDCx6p67_ASAP7_75t_R g1253 ( 
.A(n_1137),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1066),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1143),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1136),
.B(n_1129),
.Y(n_1256)
);

INVx11_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1176),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1125),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1176),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1175),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1187),
.B(n_1130),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1176),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1182),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1182),
.B(n_1125),
.Y(n_1265)
);

BUFx8_ASAP7_75t_SL g1266 ( 
.A(n_1138),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1138),
.A2(n_907),
.B1(n_932),
.B2(n_928),
.Y(n_1267)
);

CKINVDCx8_ASAP7_75t_R g1268 ( 
.A(n_1183),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1065),
.A2(n_932),
.B1(n_907),
.B2(n_845),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1150),
.A2(n_907),
.B1(n_932),
.B2(n_786),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1185),
.B(n_1161),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1116),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1072),
.A2(n_935),
.B1(n_932),
.B2(n_907),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1098),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1150),
.A2(n_907),
.B1(n_932),
.B2(n_786),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1069),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1069),
.Y(n_1277)
);

BUFx8_ASAP7_75t_L g1278 ( 
.A(n_1076),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1107),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1069),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1086),
.B(n_1168),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1156),
.A2(n_907),
.B1(n_932),
.B2(n_935),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1098),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1267),
.A2(n_1190),
.B(n_1282),
.C(n_1269),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1222),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1240),
.B(n_1223),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1241),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1241),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1223),
.B(n_1246),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1266),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1246),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1266),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1193),
.B(n_1196),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1223),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1203),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1242),
.B(n_1236),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1226),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1188),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1214),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1193),
.B(n_1217),
.Y(n_1300)
);

AO21x2_ASAP7_75t_L g1301 ( 
.A1(n_1267),
.A2(n_1256),
.B(n_1255),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1198),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1198),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1255),
.A2(n_1225),
.B(n_1247),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1208),
.A2(n_1206),
.A3(n_1205),
.B(n_1194),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1191),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1192),
.B(n_1217),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1204),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1192),
.B(n_1204),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1201),
.B(n_1200),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1201),
.B(n_1200),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1211),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1211),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1279),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1279),
.B(n_1250),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1250),
.A2(n_1280),
.B(n_1276),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1273),
.A2(n_1228),
.B(n_1235),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1270),
.A2(n_1275),
.B(n_1273),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1271),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1238),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1215),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1207),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1207),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1220),
.A2(n_1202),
.B(n_1244),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1218),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1191),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1243),
.B(n_1212),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1229),
.B(n_1219),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_1231),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1230),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_1231),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1213),
.B(n_1277),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1234),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1216),
.B(n_1283),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1189),
.B(n_1281),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1239),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1248),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1249),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1212),
.A2(n_1221),
.B(n_1261),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1286),
.B(n_1254),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1289),
.B(n_1260),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1289),
.B(n_1258),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1299),
.A2(n_1263),
.B(n_1264),
.Y(n_1344)
);

OAI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1319),
.A2(n_1251),
.B1(n_1224),
.B2(n_1209),
.C(n_1252),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1287),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1319),
.A2(n_1237),
.B1(n_1210),
.B2(n_1245),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1289),
.B(n_1216),
.Y(n_1348)
);

NOR4xp25_ASAP7_75t_SL g1349 ( 
.A(n_1284),
.B(n_1307),
.C(n_1327),
.D(n_1330),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1291),
.B(n_1216),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1291),
.B(n_1265),
.Y(n_1352)
);

INVx4_ASAP7_75t_R g1353 ( 
.A(n_1290),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1287),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_1314),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1285),
.B(n_1274),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1299),
.B(n_1262),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1297),
.B(n_1272),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1314),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1293),
.B(n_1210),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1284),
.A2(n_1245),
.B1(n_1237),
.B2(n_1232),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1295),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1311),
.A2(n_1253),
.B1(n_1195),
.B2(n_1278),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1286),
.B(n_1259),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1303),
.B(n_1272),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1294),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1286),
.B(n_1259),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1328),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1298),
.A2(n_1268),
.B(n_1233),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1305),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_L g1371 ( 
.A(n_1293),
.B(n_1199),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1301),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1300),
.B(n_1199),
.Y(n_1373)
);

AOI221xp5_ASAP7_75t_L g1374 ( 
.A1(n_1347),
.A2(n_1338),
.B1(n_1300),
.B2(n_1330),
.C(n_1332),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1348),
.B(n_1364),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_1345),
.B(n_1325),
.C(n_1311),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1361),
.B(n_1325),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1348),
.B(n_1296),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1347),
.A2(n_1338),
.B1(n_1332),
.B2(n_1312),
.C(n_1311),
.Y(n_1379)
);

OAI21xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1361),
.A2(n_1312),
.B(n_1308),
.Y(n_1380)
);

NAND4xp25_ASAP7_75t_L g1381 ( 
.A(n_1360),
.B(n_1312),
.C(n_1308),
.D(n_1320),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1363),
.B(n_1323),
.Y(n_1382)
);

OAI221xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1345),
.A2(n_1308),
.B1(n_1316),
.B2(n_1310),
.C(n_1329),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1357),
.B(n_1306),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1360),
.A2(n_1316),
.B1(n_1304),
.B2(n_1324),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1364),
.B(n_1296),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1363),
.B(n_1323),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1371),
.A2(n_1316),
.B(n_1310),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1372),
.A2(n_1292),
.B1(n_1290),
.B2(n_1339),
.Y(n_1389)
);

NAND4xp25_ASAP7_75t_L g1390 ( 
.A(n_1373),
.B(n_1329),
.C(n_1333),
.D(n_1339),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1366),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1357),
.A2(n_1304),
.B1(n_1324),
.B2(n_1323),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1373),
.A2(n_1329),
.B(n_1310),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1364),
.B(n_1367),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1357),
.A2(n_1304),
.B1(n_1324),
.B2(n_1323),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1342),
.B(n_1306),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1349),
.B(n_1318),
.C(n_1331),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1349),
.B(n_1318),
.C(n_1331),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1372),
.A2(n_1321),
.B1(n_1326),
.B2(n_1322),
.C(n_1334),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1367),
.B(n_1301),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1343),
.B(n_1322),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1367),
.B(n_1301),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1343),
.B(n_1301),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1343),
.B(n_1326),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1351),
.B(n_1288),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1346),
.B(n_1309),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1346),
.B(n_1309),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1372),
.B(n_1318),
.C(n_1321),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1358),
.A2(n_1317),
.B(n_1340),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1368),
.A2(n_1304),
.B1(n_1324),
.B2(n_1323),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_SL g1411 ( 
.A1(n_1365),
.A2(n_1336),
.B(n_1335),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1354),
.B(n_1313),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1359),
.B(n_1315),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1403),
.B(n_1341),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1391),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1391),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1376),
.A2(n_1324),
.B1(n_1323),
.B2(n_1302),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1375),
.B(n_1350),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1406),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1375),
.B(n_1350),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1403),
.B(n_1341),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1412),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1394),
.B(n_1350),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1412),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1394),
.B(n_1350),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1407),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1393),
.B(n_1356),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1414),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1396),
.B(n_1341),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1413),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1400),
.B(n_1362),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1408),
.B(n_1344),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1393),
.B(n_1355),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1390),
.B(n_1355),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1409),
.B(n_1350),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1384),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1390),
.B(n_1315),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1402),
.B(n_1350),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1405),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1405),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1402),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1378),
.B(n_1368),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1386),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1386),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1417),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1416),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1434),
.B(n_1389),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1417),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1416),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1434),
.B(n_1408),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1446),
.B(n_1440),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1441),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1436),
.A2(n_1377),
.B(n_1383),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1415),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.B(n_1410),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1443),
.B(n_1411),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1420),
.B(n_1399),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1439),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1411),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1433),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1441),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1421),
.B(n_1392),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1442),
.Y(n_1466)
);

INVxp67_ASAP7_75t_SL g1467 ( 
.A(n_1435),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1420),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1422),
.B(n_1370),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1421),
.B(n_1395),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1437),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1433),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1388),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1437),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1437),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1426),
.B(n_1388),
.Y(n_1476)
);

CKINVDCx16_ASAP7_75t_R g1477 ( 
.A(n_1444),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1455),
.B(n_1428),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1477),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1475),
.B(n_1437),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1474),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1467),
.B(n_1429),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1447),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1447),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1475),
.B(n_1444),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1477),
.B(n_1445),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1474),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1467),
.B(n_1427),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1450),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1461),
.B(n_1427),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1460),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1462),
.B(n_1445),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1450),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1454),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1428),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1449),
.A2(n_1380),
.B1(n_1389),
.B2(n_1381),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1448),
.Y(n_1497)
);

NAND2x1_ASAP7_75t_L g1498 ( 
.A(n_1452),
.B(n_1353),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1449),
.A2(n_1398),
.B(n_1397),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1460),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1438),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1423),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1462),
.B(n_1423),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1454),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1430),
.Y(n_1506)
);

AOI21xp33_ASAP7_75t_L g1507 ( 
.A1(n_1452),
.A2(n_1387),
.B(n_1382),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1464),
.Y(n_1508)
);

NAND2xp67_ASAP7_75t_L g1509 ( 
.A(n_1458),
.B(n_1337),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1448),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1468),
.B(n_1430),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1464),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1425),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1468),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1448),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1369),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1466),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1466),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1432),
.Y(n_1520)
);

CKINVDCx16_ASAP7_75t_R g1521 ( 
.A(n_1496),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.Y(n_1523)
);

CKINVDCx16_ASAP7_75t_R g1524 ( 
.A(n_1479),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1492),
.B(n_1476),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1498),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1487),
.Y(n_1527)
);

OR2x6_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1380),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1502),
.B(n_1476),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1499),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1483),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1484),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1499),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1493),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1494),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1499),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1478),
.Y(n_1538)
);

NAND2xp33_ASAP7_75t_L g1539 ( 
.A(n_1495),
.B(n_1227),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1505),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1508),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1488),
.B(n_1463),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1503),
.B(n_1476),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1518),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1490),
.B(n_1463),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1497),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1515),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1475),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1501),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1486),
.B(n_1475),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1531),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1530),
.A2(n_1500),
.B(n_1507),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1530),
.A2(n_1500),
.B(n_1379),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1506),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1534),
.B(n_1506),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1520),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1532),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1521),
.A2(n_1520),
.B1(n_1381),
.B2(n_1480),
.Y(n_1566)
);

NAND4xp25_ASAP7_75t_SL g1567 ( 
.A(n_1538),
.B(n_1374),
.C(n_1385),
.D(n_1482),
.Y(n_1567)
);

AOI322xp5_ASAP7_75t_L g1568 ( 
.A1(n_1521),
.A2(n_1472),
.A3(n_1459),
.B1(n_1470),
.B2(n_1465),
.C1(n_1512),
.C2(n_1456),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1525),
.B(n_1485),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1537),
.A2(n_1517),
.B(n_1398),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1525),
.B(n_1485),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1537),
.B(n_1397),
.C(n_1418),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1555),
.B(n_1504),
.Y(n_1573)
);

INVxp33_ASAP7_75t_L g1574 ( 
.A(n_1552),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1522),
.B(n_1480),
.Y(n_1575)
);

OAI21xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1537),
.A2(n_1475),
.B(n_1471),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1532),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1554),
.Y(n_1578)
);

OAI32xp33_ASAP7_75t_L g1579 ( 
.A1(n_1538),
.A2(n_1517),
.A3(n_1471),
.B1(n_1511),
.B2(n_1469),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1522),
.B(n_1480),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1522),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1549),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1555),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1582),
.B(n_1549),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1585)
);

AND2x2_ASAP7_75t_SL g1586 ( 
.A(n_1561),
.B(n_1539),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1574),
.B(n_1550),
.Y(n_1587)
);

OAI221xp5_ASAP7_75t_L g1588 ( 
.A1(n_1566),
.A2(n_1526),
.B1(n_1528),
.B2(n_1551),
.C(n_1547),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1578),
.B(n_1526),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1581),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1573),
.B(n_1547),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1560),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1575),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1523),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1569),
.B(n_1529),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1529),
.Y(n_1597)
);

NAND2x1_ASAP7_75t_L g1598 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1526),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1562),
.B(n_1542),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1580),
.B(n_1543),
.Y(n_1602)
);

NAND4xp25_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1568),
.C(n_1558),
.D(n_1564),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1599),
.A2(n_1583),
.B(n_1558),
.Y(n_1604)
);

AOI322xp5_ASAP7_75t_L g1605 ( 
.A1(n_1587),
.A2(n_1557),
.A3(n_1577),
.B1(n_1563),
.B2(n_1565),
.C1(n_1567),
.C2(n_1543),
.Y(n_1605)
);

AOI31xp33_ASAP7_75t_L g1606 ( 
.A1(n_1592),
.A2(n_1227),
.A3(n_1572),
.B(n_1570),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1588),
.A2(n_1579),
.B1(n_1584),
.B2(n_1589),
.C(n_1601),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1598),
.A2(n_1528),
.B1(n_1570),
.B2(n_1527),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1602),
.A2(n_1528),
.B1(n_1556),
.B2(n_1576),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1595),
.B(n_1523),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1584),
.B(n_1527),
.C(n_1528),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1595),
.B(n_1527),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1594),
.A2(n_1536),
.B1(n_1533),
.B2(n_1535),
.C(n_1546),
.Y(n_1613)
);

NOR4xp75_ASAP7_75t_SL g1614 ( 
.A(n_1585),
.B(n_1195),
.C(n_1278),
.D(n_1353),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1607),
.B(n_1593),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1610),
.B(n_1591),
.Y(n_1616)
);

NOR2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1612),
.B(n_1585),
.Y(n_1617)
);

NOR4xp25_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1594),
.C(n_1601),
.D(n_1590),
.Y(n_1618)
);

NOR4xp25_ASAP7_75t_L g1619 ( 
.A(n_1603),
.B(n_1600),
.C(n_1597),
.D(n_1596),
.Y(n_1619)
);

AOI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1608),
.A2(n_1556),
.B(n_1540),
.C(n_1533),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1613),
.Y(n_1621)
);

AOI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1611),
.A2(n_1540),
.B(n_1535),
.C(n_1536),
.Y(n_1622)
);

NOR2x1_ASAP7_75t_L g1623 ( 
.A(n_1606),
.B(n_1541),
.Y(n_1623)
);

NOR4xp75_ASAP7_75t_L g1624 ( 
.A(n_1614),
.B(n_1553),
.C(n_1586),
.D(n_1471),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1609),
.B(n_1544),
.C(n_1541),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1621),
.B(n_1605),
.C(n_1545),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1542),
.Y(n_1627)
);

NAND5xp2_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1553),
.C(n_1546),
.D(n_1545),
.E(n_1544),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1617),
.B(n_1290),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1619),
.B(n_1472),
.Y(n_1630)
);

NOR2xp67_ASAP7_75t_L g1631 ( 
.A(n_1615),
.B(n_1548),
.Y(n_1631)
);

NOR2xp67_ASAP7_75t_L g1632 ( 
.A(n_1624),
.B(n_1548),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1626),
.A2(n_1625),
.B1(n_1623),
.B2(n_1618),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1631),
.B(n_1622),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1627),
.B(n_1485),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1629),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1630),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1632),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1628),
.B(n_1548),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1638),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1633),
.A2(n_1278),
.B(n_1195),
.Y(n_1641)
);

NOR3x1_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1257),
.C(n_1197),
.Y(n_1642)
);

NOR2xp67_ASAP7_75t_L g1643 ( 
.A(n_1636),
.B(n_1292),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1635),
.B(n_1292),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1640),
.B(n_1633),
.Y(n_1645)
);

AO22x2_ASAP7_75t_L g1646 ( 
.A1(n_1641),
.A2(n_1637),
.B1(n_1639),
.B2(n_1516),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1643),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1645),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_L g1649 ( 
.A(n_1648),
.B(n_1642),
.C(n_1647),
.D(n_1644),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1649),
.A2(n_1646),
.B1(n_1516),
.B2(n_1510),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1649),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1650),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1651),
.A2(n_1510),
.B1(n_1497),
.B2(n_1471),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1653),
.B(n_1197),
.Y(n_1654)
);

AO21x2_ASAP7_75t_L g1655 ( 
.A1(n_1652),
.A2(n_1197),
.B(n_1453),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1654),
.A2(n_1471),
.B(n_1470),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1656),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_R g1658 ( 
.A1(n_1657),
.A2(n_1655),
.B1(n_1463),
.B2(n_1457),
.C(n_1451),
.Y(n_1658)
);

AOI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1457),
.B(n_1463),
.C(n_1470),
.Y(n_1659)
);


endmodule