module fake_jpeg_12030_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AND2x2_ASAP7_75t_L g7 ( 
.A(n_6),
.B(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_5),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_3),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_17),
.B(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_1),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_4),
.B1(n_9),
.B2(n_15),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_21),
.A2(n_24),
.B(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_4),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_23),
.B(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_8),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_16),
.B1(n_11),
.B2(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_11),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.C(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_19),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_21),
.B1(n_11),
.B2(n_14),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_26),
.B(n_20),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.C(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_39),
.B(n_34),
.C(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_43),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_42),
.B(n_14),
.Y(n_46)
);


endmodule