module real_jpeg_4517_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_46),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_46),
.B1(n_52),
.B2(n_57),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_46),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_2),
.A2(n_243),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_2),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_2),
.A2(n_153),
.B1(n_280),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_2),
.A2(n_280),
.B1(n_380),
.B2(n_383),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_2),
.A2(n_170),
.B1(n_280),
.B2(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_119),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_4),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_4),
.A2(n_187),
.B1(n_229),
.B2(n_270),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_4),
.A2(n_187),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_4),
.A2(n_187),
.B1(n_450),
.B2(n_451),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_50),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_5),
.A2(n_50),
.B1(n_96),
.B2(n_100),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_5),
.A2(n_50),
.B1(n_259),
.B2(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_7),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_8),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_57),
.B1(n_133),
.B2(n_180),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_8),
.A2(n_96),
.B1(n_133),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_133),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_9),
.A2(n_123),
.B1(n_274),
.B2(n_277),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_9),
.A2(n_195),
.B1(n_277),
.B2(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_9),
.A2(n_57),
.B1(n_277),
.B2(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_9),
.A2(n_277),
.B1(n_407),
.B2(n_409),
.Y(n_406)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_12),
.Y(n_497)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_13),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_13),
.Y(n_120)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_13),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_13),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_13),
.Y(n_283)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_15),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_15),
.A2(n_87),
.B1(n_101),
.B2(n_123),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_15),
.A2(n_87),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_15),
.A2(n_87),
.B1(n_145),
.B2(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_16),
.B(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_16),
.A2(n_100),
.B(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_16),
.B(n_189),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_16),
.B(n_356),
.C(n_360),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_16),
.A2(n_366),
.B1(n_367),
.B2(n_370),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_16),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_16),
.B(n_150),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_16),
.A2(n_26),
.B1(n_406),
.B2(n_414),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_17),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_495),
.B(n_498),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_483),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_215),
.A3(n_233),
.B(n_480),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_197),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_22),
.B(n_197),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_126),
.C(n_161),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_23),
.B(n_126),
.CI(n_161),
.CON(n_343),
.SN(n_343)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_90),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_24),
.A2(n_25),
.B(n_92),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_47),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_25),
.A2(n_91),
.B1(n_92),
.B2(n_125),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_25),
.A2(n_47),
.B1(n_91),
.B2(n_335),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_39),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_26),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_26),
.A2(n_256),
.B1(n_262),
.B2(n_264),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_26),
.A2(n_264),
.B(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_26),
.A2(n_173),
.B(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_26),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_26),
.A2(n_396),
.B1(n_406),
.B2(n_410),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_26),
.A2(n_39),
.B(n_298),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_27),
.Y(n_397)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_29),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_31),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_31),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_32),
.B(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_32),
.A2(n_165),
.B(n_257),
.Y(n_319)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_34),
.Y(n_418)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_35),
.Y(n_400)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_39),
.Y(n_174)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_43),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_72)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_44),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_45),
.Y(n_391)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_45),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_47),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_59),
.B(n_79),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_49),
.A2(n_60),
.B1(n_80),
.B2(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_54),
.Y(n_181)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_54),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_54),
.Y(n_452)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_55),
.Y(n_370)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_55),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_55),
.Y(n_383)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_55),
.Y(n_443)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_58),
.A2(n_137),
.B1(n_138),
.B2(n_141),
.Y(n_136)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_58),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_59),
.B(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_59),
.A2(n_81),
.B(n_157),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_59),
.A2(n_79),
.B(n_157),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_59),
.A2(n_81),
.B1(n_159),
.B2(n_179),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_59),
.A2(n_464),
.B(n_465),
.Y(n_463)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_60),
.A2(n_80),
.B1(n_365),
.B2(n_371),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_60),
.A2(n_80),
.B1(n_371),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_60),
.A2(n_80),
.B1(n_379),
.B2(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_69),
.Y(n_359)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_81),
.B(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_89),
.Y(n_432)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_115),
.B(n_121),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_93),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_93),
.A2(n_189),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_93),
.A2(n_189),
.B1(n_273),
.B2(n_278),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_94),
.A2(n_184),
.B(n_188),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_94),
.A2(n_124),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_94),
.A2(n_124),
.B1(n_184),
.B2(n_279),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_94),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_107),
.Y(n_242)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_112),
.Y(n_271)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_113),
.Y(n_246)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_114),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_121),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_123),
.Y(n_210)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_123),
.Y(n_244)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_124),
.A2(n_208),
.B(n_211),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_155),
.B(n_160),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_155),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_135),
.B1(n_150),
.B2(n_151),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_129),
.A2(n_136),
.B(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_132),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_132),
.Y(n_436)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_135),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_135),
.A2(n_151),
.B(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_135),
.A2(n_226),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_135),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_135),
.A2(n_150),
.B1(n_324),
.B2(n_447),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_135),
.A2(n_150),
.B(n_488),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_136),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_136),
.A2(n_290),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_136),
.A2(n_290),
.B1(n_294),
.B2(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_140),
.Y(n_439)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_148),
.Y(n_248)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_149),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_193),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g447 ( 
.A1(n_152),
.A2(n_366),
.B(n_434),
.Y(n_447)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_156),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_198),
.CI(n_214),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_182),
.C(n_190),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_162),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_163),
.A2(n_176),
.B1(n_177),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_163),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_173),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_166),
.Y(n_299)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_172),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g430 ( 
.A1(n_195),
.A2(n_431),
.A3(n_433),
.B1(n_434),
.B2(n_437),
.Y(n_430)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_197),
.B(n_217),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_207),
.B2(n_213),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_206),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_201),
.B(n_223),
.C(n_230),
.Y(n_492)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_206),
.C(n_207),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_204),
.A2(n_227),
.B(n_294),
.Y(n_309)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_213),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_207),
.B(n_218),
.C(n_221),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_216),
.A2(n_481),
.B(n_482),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_227),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_232),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_344),
.B(n_474),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_329),
.C(n_341),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_313),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_236),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_301),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_237),
.B(n_301),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_284),
.C(n_296),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_238),
.B(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_267),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_268),
.C(n_272),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_255),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_240),
.B(n_255),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_243),
.A3(n_245),
.B1(n_247),
.B2(n_251),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_296),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.C(n_289),
.Y(n_284)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_285),
.B(n_286),
.CI(n_289),
.CON(n_315),
.SN(n_315)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_302),
.B(n_304),
.C(n_306),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_311),
.C(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_327),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_314),
.B(n_327),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.C(n_317),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_315),
.B(n_472),
.Y(n_471)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_315),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_316),
.B(n_317),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_320),
.C(n_322),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_318),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_459)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_322),
.B(n_459),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g474 ( 
.A1(n_329),
.A2(n_341),
.B(n_475),
.C(n_478),
.D(n_479),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_340),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_330),
.B(n_340),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_334),
.C(n_339),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_333)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_342),
.B(n_343),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_343),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_469),
.B(n_473),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_454),
.B(n_468),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_426),
.B(n_453),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_392),
.B(n_425),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_374),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_349),
.B(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_364),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_364),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_435),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_385),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_384),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_384),
.C(n_385),
.Y(n_427)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_378),
.Y(n_384)
);

INVx4_ASAP7_75t_SL g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_386),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_402),
.B(n_424),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_401),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_395),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_412),
.B(n_423),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_404),
.B(n_405),
.Y(n_423)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_428),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_445),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_446),
.C(n_448),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_444),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_444),
.Y(n_462)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_442),
.Y(n_450)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_448),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_456),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_463),
.C(n_466),
.Y(n_470)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_467),
.Y(n_461)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_462),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_471),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_493),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_486),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g503 ( 
.A(n_486),
.Y(n_503)
);

FAx1_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_489),
.CI(n_492),
.CON(n_486),
.SN(n_486)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_497),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);


endmodule