module fake_jpeg_30705_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_9),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_41),
.B1(n_26),
.B2(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_54),
.B1(n_59),
.B2(n_38),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_75),
.B1(n_65),
.B2(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_66),
.B(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_60),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_37),
.B1(n_21),
.B2(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_13),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_13),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_22),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_23),
.C(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_61),
.B1(n_58),
.B2(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_58),
.B1(n_56),
.B2(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_27),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR4xp25_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_98),
.C(n_83),
.D(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_47),
.C(n_49),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_72),
.B(n_97),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.C(n_108),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_110),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_87),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_96),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_92),
.B1(n_99),
.B2(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_119),
.A2(n_107),
.B1(n_81),
.B2(n_106),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_104),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_125),
.B(n_116),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.C(n_111),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_115),
.A3(n_78),
.B1(n_94),
.B2(n_27),
.C1(n_14),
.C2(n_23),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_98),
.B1(n_72),
.B2(n_67),
.Y(n_133)
);

AOI321xp33_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_115),
.A3(n_94),
.B1(n_127),
.B2(n_126),
.C(n_120),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_121),
.B(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_135),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_122),
.B1(n_84),
.B2(n_67),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_9),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_4),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_22),
.A3(n_10),
.B1(n_11),
.B2(n_5),
.C1(n_6),
.C2(n_4),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_4),
.B1(n_6),
.B2(n_22),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_22),
.Y(n_142)
);


endmodule