module fake_jpeg_31610_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_6),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_13),
.B(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_20),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_27),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_29),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_22),
.C(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_25),
.B1(n_21),
.B2(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_60),
.B(n_61),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_18),
.B1(n_24),
.B2(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_15),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_79),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_46),
.B1(n_51),
.B2(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_51),
.B1(n_52),
.B2(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_43),
.B1(n_37),
.B2(n_52),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_64),
.C(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_90),
.B(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_98),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_76),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_71),
.C(n_77),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_91),
.B1(n_81),
.B2(n_24),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_82),
.B1(n_87),
.B2(n_86),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_1),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_100),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_112),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_67),
.B1(n_72),
.B2(n_91),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_84),
.B(n_24),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_84),
.C(n_2),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_117),
.C(n_107),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_109),
.B1(n_108),
.B2(n_111),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_106),
.B(n_7),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_112),
.C(n_4),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_115),
.C(n_114),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_125),
.B(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_8),
.Y(n_128)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_5),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_9),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_11),
.Y(n_130)
);


endmodule