module fake_jpeg_15969_n_120 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_14),
.B1(n_21),
.B2(n_17),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_39),
.B1(n_29),
.B2(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_22),
.B1(n_18),
.B2(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_17),
.B1(n_21),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_10),
.B1(n_22),
.B2(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_24),
.B(n_28),
.C(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_60),
.B1(n_28),
.B2(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_15),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_32),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_12),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_31),
.B1(n_12),
.B2(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_46),
.B1(n_43),
.B2(n_50),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_1),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_80),
.B1(n_83),
.B2(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_46),
.B1(n_51),
.B2(n_56),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_46),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_70),
.B(n_69),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_90),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_72),
.C(n_69),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_89),
.C(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_80),
.B1(n_77),
.B2(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_96),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_107),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_100),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_111),
.Y(n_112)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_101),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_116),
.B(n_112),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_113),
.B(n_75),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_75),
.Y(n_120)
);


endmodule