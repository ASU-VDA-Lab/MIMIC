module fake_jpeg_16022_n_80 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_20),
.C(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_28),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_12),
.B1(n_16),
.B2(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_29),
.B1(n_14),
.B2(n_11),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_16),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_19),
.Y(n_36)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_26),
.CI(n_15),
.CON(n_44),
.SN(n_44)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_25),
.B1(n_11),
.B2(n_12),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_23),
.B1(n_18),
.B2(n_4),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_50),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_24),
.C(n_26),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_33),
.B1(n_23),
.B2(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_57),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_37),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_50),
.C(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.C(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_44),
.C(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_51),
.B1(n_52),
.B2(n_49),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_51),
.C(n_44),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_69),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_51),
.B(n_68),
.Y(n_73)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_67),
.A3(n_69),
.B1(n_37),
.B2(n_49),
.C(n_18),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_71),
.C(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_77),
.Y(n_80)
);


endmodule