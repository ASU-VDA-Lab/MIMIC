module fake_ibex_1266_n_2027 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_407, n_102, n_52, n_448, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2027);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2027;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_1930;
wire n_1234;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_1971;
wire n_879;
wire n_1957;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_1980;
wire n_462;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2006;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1982;
wire n_1334;
wire n_1963;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2010;
wire n_1470;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1967;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_1679;
wire n_1497;
wire n_2002;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_2000;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1976;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2012;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1961;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_753;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_1168;
wire n_865;
wire n_2013;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_955;
wire n_1333;
wire n_1916;
wire n_952;
wire n_1675;
wire n_1947;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_51),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_398),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_158),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_426),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_233),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_25),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_106),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_291),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_169),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_2),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_34),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_438),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_218),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_192),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_274),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_193),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_207),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_379),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_377),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_208),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_425),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_459),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_113),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_15),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_333),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_312),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_282),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_153),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_428),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_74),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_149),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_219),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_137),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_259),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_200),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_182),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_120),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_266),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_372),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_195),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_103),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_374),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_143),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_453),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_297),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_45),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_422),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_190),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_356),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_104),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_43),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_449),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_281),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_345),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_183),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_241),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_151),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_317),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_458),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_16),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_344),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_447),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_421),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_332),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_363),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_411),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_14),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_455),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_308),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_57),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_287),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_457),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_321),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_424),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_55),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_138),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_255),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_175),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_204),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_38),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_404),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_232),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_442),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_366),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_283),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_78),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_419),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_359),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_444),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_38),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_101),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_0),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_284),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_83),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_102),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_328),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_52),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_278),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_66),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_415),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_384),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_248),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_417),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_320),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_206),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g575 ( 
.A(n_72),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_342),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_434),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_413),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_407),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_341),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_77),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_268),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_93),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_91),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_32),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_111),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_405),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_215),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_152),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_136),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g591 ( 
.A(n_201),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_89),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_197),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_156),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_335),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_117),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_121),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_180),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_258),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_173),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_365),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_10),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_456),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_322),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_452),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_47),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_383),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_164),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_8),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_17),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_382),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_108),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_140),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_65),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_223),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_367),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_227),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_181),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_348),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_310),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_211),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_163),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_295),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_12),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_3),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_97),
.Y(n_627)
);

BUFx5_ASAP7_75t_L g628 ( 
.A(n_19),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_141),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_172),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_162),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_1),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_7),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_440),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_79),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_389),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_427),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_288),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_83),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_296),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_396),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_4),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_290),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_443),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_431),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_15),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_111),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_76),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_184),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_430),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_388),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_95),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_159),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_361),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_116),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_11),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_81),
.Y(n_657)
);

BUFx10_ASAP7_75t_L g658 ( 
.A(n_47),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_1),
.Y(n_659)
);

CKINVDCx12_ASAP7_75t_R g660 ( 
.A(n_66),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_330),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_86),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_96),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_78),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_331),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_349),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_106),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_67),
.Y(n_668)
);

BUFx5_ASAP7_75t_L g669 ( 
.A(n_107),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_18),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_51),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_294),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_133),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_44),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_420),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_338),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_307),
.Y(n_677)
);

BUFx6f_ASAP7_75t_SL g678 ( 
.A(n_221),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_26),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_329),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_179),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_353),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_85),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_454),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_399),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_311),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_116),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_166),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_20),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_416),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_124),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_293),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_48),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_441),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_118),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_148),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_93),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_237),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_378),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_168),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_235),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_306),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_275),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_276),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_189),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_257),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_450),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_325),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_36),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_313),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_214),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_410),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_44),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_16),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_402),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_408),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_423),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_68),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_397),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_157),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_304),
.Y(n_721)
);

CKINVDCx16_ASAP7_75t_R g722 ( 
.A(n_400),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_435),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_433),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_262),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_91),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_429),
.Y(n_727)
);

BUFx10_ASAP7_75t_L g728 ( 
.A(n_401),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_21),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_27),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_20),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_174),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_5),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_142),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_68),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_300),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_437),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_395),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_412),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_391),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_354),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_29),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_375),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_12),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_409),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_56),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_350),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_92),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_90),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_80),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_129),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_86),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_108),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_439),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_104),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_264),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_101),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_171),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_123),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_132),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_279),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_234),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_238),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_393),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_187),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_436),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_461),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_649),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_491),
.Y(n_769)
);

NOR2xp67_ASAP7_75t_L g770 ( 
.A(n_472),
.B(n_0),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_649),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_597),
.Y(n_772)
);

INVxp33_ASAP7_75t_SL g773 ( 
.A(n_597),
.Y(n_773)
);

CKINVDCx16_ASAP7_75t_R g774 ( 
.A(n_592),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_575),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_744),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_721),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_721),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_575),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_549),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_483),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_516),
.B(n_2),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_714),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_714),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_511),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_660),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_671),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_718),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_651),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_718),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_581),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_514),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_581),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_628),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_628),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_628),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_630),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_557),
.B(n_3),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_628),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_651),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_762),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_628),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_603),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_669),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_687),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_626),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_634),
.B(n_4),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_669),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_638),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_650),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_726),
.B(n_5),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_762),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_753),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_669),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_652),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_674),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_669),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_467),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_669),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_693),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_752),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_669),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_468),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_460),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_499),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_705),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_471),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_717),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_763),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_711),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_722),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_757),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_510),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_486),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_677),
.B(n_6),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_492),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_503),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_524),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_515),
.Y(n_841)
);

INVxp33_ASAP7_75t_SL g842 ( 
.A(n_535),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_532),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_465),
.B(n_6),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_591),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_591),
.Y(n_846)
);

INVxp67_ASAP7_75t_SL g847 ( 
.A(n_540),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_545),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_567),
.Y(n_849)
);

BUFx6f_ASAP7_75t_SL g850 ( 
.A(n_602),
.Y(n_850)
);

INVxp33_ASAP7_75t_L g851 ( 
.A(n_586),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_610),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_632),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_489),
.B(n_7),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_678),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_552),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_474),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_558),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_635),
.B(n_8),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_639),
.Y(n_860)
);

BUFx2_ASAP7_75t_SL g861 ( 
.A(n_678),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_642),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_559),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_485),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_560),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_646),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_562),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_470),
.Y(n_868)
);

INVxp33_ASAP7_75t_SL g869 ( 
.A(n_563),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_648),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_659),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_583),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_584),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_663),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_585),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_596),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_679),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_857),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_795),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_807),
.B(n_547),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_768),
.B(n_691),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_771),
.B(n_462),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_772),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_789),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_791),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_796),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_826),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_797),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_802),
.B(n_607),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_784),
.B(n_485),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_787),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_800),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_SL g893 ( 
.A(n_781),
.B(n_611),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_777),
.B(n_613),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_788),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_778),
.B(n_463),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_790),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_855),
.B(n_602),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_790),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_865),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_857),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_857),
.Y(n_902)
);

OA21x2_ASAP7_75t_L g903 ( 
.A1(n_801),
.A2(n_538),
.B(n_470),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_804),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_803),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_867),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_857),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_868),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_773),
.A2(n_615),
.B1(n_627),
.B2(n_625),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_803),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_821),
.B(n_633),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_814),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_851),
.B(n_658),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_783),
.B(n_695),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_814),
.B(n_525),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_806),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_810),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_851),
.B(n_658),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_816),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_782),
.B(n_525),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_850),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_819),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_824),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_815),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_874),
.B(n_655),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_868),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_825),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_845),
.B(n_656),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_827),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_835),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_829),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_794),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_841),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_785),
.B(n_644),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_854),
.Y(n_936)
);

OA21x2_ASAP7_75t_L g937 ( 
.A1(n_843),
.A2(n_543),
.B(n_538),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_848),
.Y(n_938)
);

CKINVDCx8_ASAP7_75t_R g939 ( 
.A(n_774),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_776),
.B(n_644),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_842),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_849),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_820),
.B(n_697),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_852),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_846),
.B(n_657),
.Y(n_945)
);

XOR2x2_ASAP7_75t_SL g946 ( 
.A(n_818),
.B(n_713),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_853),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_860),
.Y(n_948)
);

OAI21x1_ASAP7_75t_L g949 ( 
.A1(n_866),
.A2(n_654),
.B(n_543),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_869),
.B(n_728),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_870),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_859),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_871),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_877),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_873),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_847),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_862),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_876),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_844),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_844),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_728),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_782),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_799),
.Y(n_963)
);

BUFx8_ASAP7_75t_L g964 ( 
.A(n_850),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_836),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_856),
.B(n_742),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_861),
.B(n_662),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_799),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_770),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_875),
.B(n_748),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_832),
.B(n_664),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_833),
.B(n_667),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_809),
.B(n_668),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_838),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_809),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_813),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_837),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_837),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_786),
.B(n_683),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_767),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_775),
.B(n_750),
.Y(n_981)
);

INVx6_ASAP7_75t_L g982 ( 
.A(n_864),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_769),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_840),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_779),
.B(n_689),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_780),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_779),
.B(n_464),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_864),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_858),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_863),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_872),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_798),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_811),
.A2(n_730),
.B1(n_733),
.B2(n_709),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_812),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_828),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_830),
.B(n_469),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_831),
.B(n_735),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_818),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_793),
.B(n_746),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_805),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_834),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_808),
.B(n_749),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_817),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_822),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_823),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_789),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_802),
.B(n_473),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_772),
.B(n_751),
.Y(n_1008)
);

INVxp67_ASAP7_75t_L g1009 ( 
.A(n_826),
.Y(n_1009)
);

NAND2x1_ASAP7_75t_L g1010 ( 
.A(n_821),
.B(n_654),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_802),
.B(n_476),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_789),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_857),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_789),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_789),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_789),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_790),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_789),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_795),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_789),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_789),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_789),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_768),
.B(n_755),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_818),
.A2(n_647),
.B1(n_670),
.B2(n_565),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_767),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_795),
.Y(n_1026)
);

CKINVDCx16_ASAP7_75t_R g1027 ( 
.A(n_781),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_790),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_795),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_802),
.B(n_477),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_795),
.A2(n_754),
.B(n_719),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_772),
.B(n_759),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_795),
.A2(n_754),
.B(n_719),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_802),
.B(n_479),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_795),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_795),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_795),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_857),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_768),
.B(n_729),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_807),
.B(n_475),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_857),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_768),
.B(n_729),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_826),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_825),
.B(n_731),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_790),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_964),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_908),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_956),
.A2(n_729),
.B1(n_738),
.B2(n_478),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_L g1049 ( 
.A(n_920),
.B(n_480),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_921),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_883),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_982),
.B(n_729),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_978),
.A2(n_487),
.B1(n_502),
.B2(n_490),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_893),
.A2(n_507),
.B1(n_513),
.B2(n_506),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_908),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_927),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_964),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_963),
.B(n_481),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_927),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1039),
.Y(n_1061)
);

AND2x2_ASAP7_75t_SL g1062 ( 
.A(n_1027),
.B(n_517),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_913),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_1025),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_927),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_963),
.B(n_482),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_933),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1039),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_963),
.B(n_484),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_966),
.A2(n_520),
.B1(n_527),
.B2(n_518),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1042),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1042),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_914),
.B(n_548),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_SL g1074 ( 
.A(n_921),
.B(n_488),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_942),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_918),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_933),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_942),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_936),
.B(n_914),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_933),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_942),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_936),
.B(n_493),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_936),
.B(n_494),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_949),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_897),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_962),
.A2(n_550),
.B1(n_553),
.B2(n_541),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_1009),
.B(n_548),
.Y(n_1087)
);

AND3x2_ASAP7_75t_L g1088 ( 
.A(n_965),
.B(n_974),
.C(n_906),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_968),
.B(n_495),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1044),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_899),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_975),
.B(n_497),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_905),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_977),
.B(n_498),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_980),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_910),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_1017),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_957),
.A2(n_561),
.B1(n_564),
.B2(n_555),
.Y(n_1099)
);

INVx4_ASAP7_75t_L g1100 ( 
.A(n_955),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1017),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_941),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_973),
.B(n_466),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1028),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1031),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1028),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1045),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_912),
.Y(n_1108)
);

INVx4_ASAP7_75t_SL g1109 ( 
.A(n_915),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_959),
.A2(n_573),
.B1(n_574),
.B2(n_569),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_915),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_881),
.B(n_500),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1033),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_982),
.B(n_587),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_980),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_915),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_966),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_932),
.B(n_9),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_881),
.B(n_501),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1045),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_939),
.Y(n_1121)
);

BUFx10_ASAP7_75t_L g1122 ( 
.A(n_970),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_970),
.A2(n_890),
.B1(n_1023),
.B2(n_884),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_900),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_958),
.Y(n_1125)
);

INVxp67_ASAP7_75t_SL g1126 ( 
.A(n_1043),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_926),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_915),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1023),
.B(n_504),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_925),
.B(n_505),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_926),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1010),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_891),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_937),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_R g1135 ( 
.A(n_998),
.B(n_508),
.Y(n_1135)
);

OAI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_885),
.A2(n_590),
.B1(n_599),
.B2(n_593),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1004),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1006),
.A2(n_609),
.B1(n_612),
.B2(n_605),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_937),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_903),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_895),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_903),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_924),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_943),
.B(n_509),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_959),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_947),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_943),
.B(n_959),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1010),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_953),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1008),
.B(n_579),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1032),
.B(n_579),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_980),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_953),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_887),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_SL g1155 ( 
.A1(n_954),
.A2(n_616),
.B(n_614),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_960),
.B(n_512),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1012),
.A2(n_618),
.B1(n_620),
.B2(n_617),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_969),
.B(n_594),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_954),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_960),
.B(n_519),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_960),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_951),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1014),
.B(n_594),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_999),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1015),
.A2(n_623),
.B1(n_637),
.B2(n_621),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_928),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_930),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_983),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_920),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_931),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_934),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1007),
.B(n_521),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_938),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1011),
.B(n_522),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_929),
.B(n_945),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_944),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_894),
.B(n_523),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1016),
.B(n_643),
.Y(n_1178)
);

INVx6_ASAP7_75t_L g1179 ( 
.A(n_1004),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_920),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_948),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_961),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_889),
.B(n_496),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_879),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_981),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_917),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_952),
.Y(n_1187)
);

NAND2xp33_ASAP7_75t_SL g1188 ( 
.A(n_967),
.B(n_526),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_886),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1018),
.A2(n_680),
.B1(n_685),
.B2(n_682),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_920),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_888),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_952),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_892),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1030),
.B(n_528),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_979),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1020),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1021),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1022),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_976),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_904),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_911),
.B(n_571),
.Y(n_1202)
);

CKINVDCx16_ASAP7_75t_R g1203 ( 
.A(n_940),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_1034),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_878),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_916),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_983),
.B(n_686),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1002),
.B(n_9),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_882),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_896),
.B(n_1040),
.Y(n_1210)
);

INVx8_ASAP7_75t_L g1211 ( 
.A(n_1004),
.Y(n_1211)
);

OR2x6_ASAP7_75t_L g1212 ( 
.A(n_983),
.B(n_688),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1000),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_880),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_922),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_919),
.B(n_529),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_971),
.B(n_595),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1019),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1026),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_923),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1029),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1035),
.A2(n_702),
.B1(n_708),
.B2(n_701),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_972),
.B(n_530),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1036),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1037),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_935),
.B(n_643),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_950),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_909),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_986),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_878),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_878),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_898),
.B(n_531),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_997),
.B(n_533),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_986),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_986),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_981),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_992),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_993),
.B(n_715),
.C(n_710),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_992),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_901),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_L g1241 ( 
.A(n_985),
.B(n_727),
.C(n_723),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_994),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_992),
.Y(n_1243)
);

XNOR2xp5_ASAP7_75t_L g1244 ( 
.A(n_984),
.B(n_10),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_996),
.B(n_534),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_987),
.B(n_536),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_995),
.B(n_619),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_901),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_946),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_988),
.B(n_537),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1041),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1024),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_901),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_991),
.B(n_736),
.C(n_732),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_902),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_902),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_989),
.B(n_539),
.Y(n_1257)
);

AND2x6_ASAP7_75t_L g1258 ( 
.A(n_990),
.B(n_712),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1000),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_902),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1000),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1001),
.B(n_542),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1003),
.B(n_544),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_907),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_907),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_998),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1005),
.B(n_712),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_907),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1013),
.B(n_546),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1013),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1013),
.B(n_551),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_1038),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1038),
.A2(n_743),
.B1(n_756),
.B2(n_745),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1038),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1041),
.B(n_556),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1041),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_949),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_914),
.B(n_737),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1039),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_936),
.B(n_566),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1171),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1204),
.B(n_568),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1161),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1209),
.B(n_570),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1252),
.A2(n_758),
.B(n_765),
.C(n_760),
.Y(n_1285)
);

AO221x1_ASAP7_75t_L g1286 ( 
.A1(n_1054),
.A2(n_1154),
.B1(n_1138),
.B2(n_1190),
.C(n_1136),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1051),
.B(n_1126),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1123),
.A2(n_572),
.B1(n_578),
.B2(n_577),
.C(n_576),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1161),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1171),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1175),
.B(n_580),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1117),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1161),
.Y(n_1293)
);

INVxp67_ASAP7_75t_SL g1294 ( 
.A(n_1124),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1117),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1176),
.B(n_582),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1074),
.B(n_588),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1063),
.B(n_589),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1176),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1122),
.B(n_598),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1125),
.B(n_11),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1067),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1067),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1067),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1122),
.B(n_600),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1181),
.B(n_601),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1164),
.B(n_13),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1181),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1182),
.B(n_604),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1102),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1196),
.B(n_606),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1058),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1210),
.B(n_608),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1091),
.B(n_622),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1180),
.B(n_624),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1180),
.B(n_629),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1046),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1143),
.B(n_631),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1052),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_L g1320 ( 
.A(n_1134),
.B(n_636),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1194),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1145),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1197),
.B(n_640),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1194),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1145),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1153),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1052),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1228),
.A2(n_645),
.B1(n_653),
.B2(n_641),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1114),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1100),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1198),
.B(n_1199),
.Y(n_1332)
);

NOR3xp33_ASAP7_75t_L g1333 ( 
.A(n_1203),
.B(n_665),
.C(n_661),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1076),
.B(n_666),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1227),
.B(n_672),
.Y(n_1335)
);

BUFx5_ASAP7_75t_L g1336 ( 
.A(n_1113),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1114),
.B(n_13),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1144),
.B(n_675),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1050),
.B(n_1100),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1159),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1215),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1173),
.B(n_676),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1166),
.B(n_681),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1167),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1170),
.B(n_684),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1220),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1073),
.B(n_690),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1073),
.B(n_692),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1278),
.B(n_694),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1186),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1050),
.B(n_737),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1112),
.B(n_1119),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1185),
.B(n_14),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1211),
.Y(n_1354)
);

OR2x6_ASAP7_75t_L g1355 ( 
.A(n_1211),
.B(n_766),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1278),
.B(n_1214),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1129),
.B(n_696),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1150),
.B(n_698),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1151),
.B(n_699),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1118),
.B(n_1064),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1185),
.B(n_700),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1186),
.A2(n_704),
.B1(n_706),
.B2(n_703),
.Y(n_1362)
);

BUFx5_ASAP7_75t_L g1363 ( 
.A(n_1113),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1147),
.A2(n_766),
.B(n_19),
.C(n_17),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1133),
.B(n_707),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1141),
.B(n_716),
.Y(n_1366)
);

AOI221xp5_ASAP7_75t_L g1367 ( 
.A1(n_1165),
.A2(n_725),
.B1(n_734),
.B2(n_724),
.C(n_720),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1134),
.Y(n_1368)
);

BUFx8_ASAP7_75t_L g1369 ( 
.A(n_1266),
.Y(n_1369)
);

BUFx10_ASAP7_75t_L g1370 ( 
.A(n_1088),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1215),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1259),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1148),
.B(n_1132),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1061),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1207),
.Y(n_1375)
);

AND2x6_ASAP7_75t_SL g1376 ( 
.A(n_1207),
.B(n_18),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1068),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1071),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1072),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1279),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1236),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1084),
.A2(n_740),
.B(n_739),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_L g1383 ( 
.A(n_1134),
.B(n_741),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1162),
.B(n_747),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1236),
.B(n_761),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1148),
.B(n_474),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1148),
.B(n_474),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1146),
.Y(n_1388)
);

AND2x6_ASAP7_75t_SL g1389 ( 
.A(n_1212),
.B(n_21),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1087),
.B(n_22),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1079),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1183),
.B(n_22),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1105),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1132),
.B(n_474),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1242),
.B(n_1257),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1238),
.A2(n_673),
.B1(n_554),
.B2(n_764),
.C(n_25),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1070),
.B(n_23),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1262),
.B(n_1263),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1116),
.B(n_554),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1103),
.B(n_23),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1131),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1131),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1155),
.A2(n_764),
.B(n_673),
.C(n_554),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1085),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1202),
.B(n_24),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1250),
.B(n_24),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1116),
.B(n_554),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1078),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1212),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1187),
.B(n_26),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1193),
.B(n_27),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1139),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1226),
.B(n_28),
.Y(n_1413)
);

AND2x4_ASAP7_75t_SL g1414 ( 
.A(n_1229),
.B(n_673),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1105),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1053),
.B(n_28),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1092),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1217),
.B(n_29),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_SL g1419 ( 
.A(n_1128),
.B(n_673),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1128),
.B(n_1111),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1247),
.B(n_764),
.C(n_30),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1139),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1062),
.A2(n_764),
.B1(n_32),
.B2(n_30),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1090),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1246),
.B(n_31),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1049),
.B(n_31),
.C(n_33),
.Y(n_1426)
);

AOI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1241),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1163),
.B(n_35),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1097),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1178),
.B(n_36),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1261),
.B(n_37),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1229),
.B(n_37),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1086),
.B(n_39),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1200),
.B(n_39),
.Y(n_1434)
);

NOR2xp67_ASAP7_75t_L g1435 ( 
.A(n_1121),
.B(n_40),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1089),
.B(n_40),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1179),
.Y(n_1437)
);

CKINVDCx11_ASAP7_75t_R g1438 ( 
.A(n_1249),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1094),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_SL g1440 ( 
.A(n_1152),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1105),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1101),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1093),
.B(n_41),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1095),
.B(n_41),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1099),
.B(n_42),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1137),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1234),
.B(n_42),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1111),
.B(n_1169),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1104),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1108),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1106),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1135),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1224),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1157),
.B(n_43),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1130),
.B(n_45),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1234),
.B(n_1243),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1225),
.B(n_46),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1267),
.B(n_46),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1078),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1107),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1267),
.B(n_1172),
.Y(n_1461)
);

INVx8_ASAP7_75t_L g1462 ( 
.A(n_1213),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1127),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1111),
.B(n_48),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1208),
.B(n_49),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1258),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1174),
.B(n_50),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1120),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1098),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_SL g1470 ( 
.A(n_1169),
.B(n_53),
.Y(n_1470)
);

NOR2xp67_ASAP7_75t_SL g1471 ( 
.A(n_1179),
.B(n_53),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1277),
.A2(n_134),
.B(n_131),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1158),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1195),
.B(n_54),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1258),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1475)
);

CKINVDCx11_ASAP7_75t_R g1476 ( 
.A(n_1168),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1294),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1287),
.B(n_1158),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1281),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1319),
.B(n_1375),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1332),
.B(n_1222),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1330),
.B(n_1243),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1397),
.A2(n_1048),
.B(n_1239),
.C(n_1177),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1290),
.A2(n_1140),
.B1(n_1142),
.B2(n_1110),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1331),
.B(n_1292),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_SL g1486 ( 
.A1(n_1403),
.A2(n_1277),
.B(n_1191),
.C(n_1081),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1386),
.A2(n_1387),
.B(n_1394),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1398),
.A2(n_1216),
.B(n_1280),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1344),
.B(n_1254),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1412),
.A2(n_1422),
.B(n_1308),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1400),
.A2(n_1191),
.B(n_1066),
.C(n_1069),
.Y(n_1491)
);

NOR2xp67_ASAP7_75t_L g1492 ( 
.A(n_1312),
.B(n_1244),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1461),
.A2(n_1059),
.B(n_1233),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1331),
.B(n_1096),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1331),
.B(n_1235),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1299),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1408),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1350),
.A2(n_1160),
.B(n_1156),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_L g1499 ( 
.A(n_1336),
.B(n_1258),
.Y(n_1499)
);

CKINVDCx6p67_ASAP7_75t_R g1500 ( 
.A(n_1354),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1339),
.B(n_1237),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1369),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1346),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1404),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1295),
.B(n_1096),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1286),
.B(n_1258),
.Y(n_1506)
);

AO21x1_ASAP7_75t_L g1507 ( 
.A1(n_1472),
.A2(n_1075),
.B(n_1082),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1462),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1417),
.B(n_1223),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1369),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1296),
.A2(n_1083),
.B(n_1184),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1306),
.A2(n_1192),
.B(n_1189),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1439),
.B(n_1098),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1450),
.B(n_1201),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1307),
.B(n_1337),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1326),
.B(n_1327),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1395),
.A2(n_1218),
.B(n_1206),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1340),
.B(n_1219),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1453),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1356),
.B(n_1115),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1388),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1393),
.A2(n_1221),
.B(n_1055),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1374),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1393),
.A2(n_1056),
.B(n_1047),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1465),
.B(n_1245),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1328),
.B(n_1339),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1393),
.A2(n_1077),
.B(n_1057),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1291),
.A2(n_1273),
.B1(n_1115),
.B2(n_1065),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1409),
.B(n_1188),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1413),
.A2(n_1065),
.B1(n_1060),
.B2(n_1232),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1436),
.A2(n_1080),
.B(n_1060),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1313),
.B(n_1109),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1377),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1378),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_SL g1535 ( 
.A(n_1370),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1462),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1476),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1418),
.A2(n_1269),
.B(n_1275),
.C(n_1271),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1379),
.B(n_1109),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1428),
.A2(n_1251),
.B1(n_1231),
.B2(n_1240),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1415),
.A2(n_1231),
.B(n_1253),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1380),
.B(n_1251),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1415),
.A2(n_1274),
.B(n_1270),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1473),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1468),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1415),
.A2(n_1256),
.B(n_1230),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1301),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1317),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1406),
.A2(n_1425),
.B(n_1364),
.C(n_1467),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1298),
.B(n_1352),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1454),
.A2(n_1264),
.B(n_1276),
.C(n_1240),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1441),
.A2(n_1265),
.B(n_1260),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1424),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1441),
.A2(n_1264),
.B(n_1276),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1441),
.A2(n_1248),
.B(n_1205),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1282),
.B(n_57),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1430),
.B(n_58),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1343),
.A2(n_1248),
.B(n_1205),
.Y(n_1558)
);

NOR2xp67_ASAP7_75t_L g1559 ( 
.A(n_1452),
.B(n_58),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1368),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1284),
.B(n_1353),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1390),
.A2(n_1458),
.B1(n_1360),
.B2(n_1416),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1345),
.A2(n_1248),
.B(n_1205),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1310),
.B(n_59),
.Y(n_1564)
);

AO21x1_ASAP7_75t_L g1565 ( 
.A1(n_1470),
.A2(n_139),
.B(n_135),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1365),
.A2(n_1268),
.B(n_1255),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1368),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1433),
.A2(n_1268),
.B1(n_1255),
.B2(n_61),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1366),
.A2(n_1268),
.B(n_1255),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1391),
.B(n_59),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1410),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1285),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1358),
.B(n_60),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1373),
.A2(n_1272),
.B(n_145),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1318),
.A2(n_1272),
.B(n_146),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1372),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1359),
.B(n_62),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1288),
.B(n_1381),
.Y(n_1578)
);

AOI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1399),
.A2(n_147),
.B(n_144),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1445),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1355),
.B(n_63),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1443),
.A2(n_154),
.B(n_150),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1474),
.A2(n_160),
.B(n_155),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1355),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1411),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1457),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1362),
.B(n_64),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1347),
.B(n_67),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1323),
.B(n_69),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1455),
.A2(n_165),
.B(n_161),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1405),
.B(n_69),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1309),
.B(n_70),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1392),
.B(n_70),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1466),
.A2(n_1475),
.B1(n_1444),
.B2(n_1423),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1335),
.B(n_71),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1434),
.A2(n_1431),
.B(n_1447),
.C(n_1432),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1384),
.A2(n_170),
.B(n_167),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1463),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1351),
.B(n_71),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1367),
.B(n_72),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1429),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1351),
.B(n_1348),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1283),
.A2(n_177),
.B(n_176),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1349),
.B(n_73),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1289),
.A2(n_185),
.B(n_178),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1437),
.B(n_73),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1336),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1338),
.B(n_1357),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1293),
.A2(n_188),
.B(n_186),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1311),
.B(n_74),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1342),
.B(n_75),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1382),
.A2(n_194),
.B(n_191),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1333),
.B(n_75),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_SL g1614 ( 
.A1(n_1407),
.A2(n_1419),
.B(n_1464),
.C(n_1420),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1334),
.B(n_76),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1300),
.B(n_77),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1361),
.B(n_79),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1305),
.B(n_80),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1376),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1385),
.B(n_81),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1321),
.B(n_82),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1324),
.B(n_82),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1446),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1442),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1449),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1396),
.A2(n_87),
.B(n_84),
.C(n_85),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_R g1627 ( 
.A(n_1500),
.B(n_1389),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1562),
.A2(n_1329),
.B(n_1421),
.C(n_1314),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1549),
.A2(n_1368),
.B(n_1320),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1581),
.B(n_1370),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1488),
.A2(n_1426),
.B(n_1427),
.C(n_1471),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1503),
.B(n_1341),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1504),
.Y(n_1633)
);

OR2x2_ASAP7_75t_SL g1634 ( 
.A(n_1584),
.B(n_1438),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1479),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1502),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1508),
.B(n_1322),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1478),
.A2(n_1414),
.B1(n_1322),
.B2(n_1325),
.Y(n_1638)
);

CKINVDCx11_ASAP7_75t_R g1639 ( 
.A(n_1510),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1481),
.A2(n_1325),
.B1(n_1456),
.B2(n_1297),
.Y(n_1640)
);

NOR3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1537),
.B(n_1316),
.C(n_1315),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1519),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1496),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1516),
.B(n_1371),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1581),
.B(n_1336),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1594),
.A2(n_1435),
.B1(n_1440),
.B2(n_1451),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1477),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1440),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1486),
.A2(n_1383),
.B(n_1303),
.Y(n_1649)
);

A2O1A1Ixp33_ASAP7_75t_SL g1650 ( 
.A1(n_1615),
.A2(n_1459),
.B(n_1408),
.C(n_1304),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_SL g1651 ( 
.A(n_1616),
.B(n_1448),
.C(n_84),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1550),
.A2(n_1402),
.B1(n_1469),
.B2(n_1401),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1596),
.A2(n_1302),
.B(n_1460),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1578),
.B(n_1459),
.Y(n_1654)
);

OAI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1619),
.A2(n_1363),
.B1(n_1336),
.B2(n_89),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1545),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1515),
.B(n_1336),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1495),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1558),
.A2(n_1363),
.B(n_198),
.Y(n_1659)
);

INVxp67_ASAP7_75t_SL g1660 ( 
.A(n_1484),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1547),
.B(n_87),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1533),
.Y(n_1662)
);

AO21x1_ASAP7_75t_L g1663 ( 
.A1(n_1506),
.A2(n_1363),
.B(n_88),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1508),
.B(n_88),
.Y(n_1664)
);

BUFx12f_ASAP7_75t_L g1665 ( 
.A(n_1548),
.Y(n_1665)
);

NOR3xp33_ASAP7_75t_L g1666 ( 
.A(n_1572),
.B(n_90),
.C(n_92),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1523),
.B(n_1363),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1598),
.Y(n_1668)
);

AOI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1507),
.A2(n_1363),
.B(n_199),
.Y(n_1669)
);

O2A1O1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1561),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1576),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_SL g1672 ( 
.A(n_1607),
.B(n_94),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1571),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1563),
.A2(n_1569),
.B(n_1566),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1499),
.A2(n_202),
.B(n_196),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1585),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1495),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1607),
.A2(n_1586),
.B1(n_1556),
.B2(n_1518),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1606),
.B(n_100),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1535),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1602),
.B(n_102),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1534),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1526),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_1683)
);

O2A1O1Ixp5_ASAP7_75t_SL g1684 ( 
.A1(n_1587),
.A2(n_1485),
.B(n_1582),
.C(n_1505),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1520),
.B(n_105),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1538),
.A2(n_205),
.B(n_203),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1525),
.B(n_109),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1522),
.A2(n_210),
.B(n_209),
.Y(n_1688)
);

CKINVDCx8_ASAP7_75t_R g1689 ( 
.A(n_1606),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1480),
.B(n_1526),
.Y(n_1690)
);

OAI22x1_ASAP7_75t_L g1691 ( 
.A1(n_1613),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1501),
.B(n_110),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1521),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1512),
.A2(n_213),
.B(n_212),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1489),
.B(n_112),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1511),
.A2(n_217),
.B(n_216),
.Y(n_1696)
);

AOI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1555),
.A2(n_222),
.B(n_220),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1588),
.B(n_113),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1553),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1544),
.B(n_114),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1494),
.B(n_114),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1623),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1514),
.B(n_115),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1618),
.B(n_115),
.C(n_117),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_SL g1705 ( 
.A(n_1610),
.B(n_118),
.C(n_119),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1509),
.B(n_119),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1564),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1560),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1592),
.B(n_120),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_SL g1710 ( 
.A(n_1617),
.B(n_121),
.C(n_122),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1501),
.B(n_122),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1626),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1601),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1624),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1517),
.A2(n_125),
.B(n_126),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1536),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1600),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1513),
.B(n_127),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1483),
.A2(n_128),
.B(n_130),
.C(n_224),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1679),
.A2(n_1620),
.B(n_1595),
.C(n_1604),
.Y(n_1720)
);

AO31x2_ASAP7_75t_L g1721 ( 
.A1(n_1674),
.A2(n_1565),
.A3(n_1568),
.B(n_1583),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1633),
.B(n_1625),
.Y(n_1722)
);

AO31x2_ASAP7_75t_L g1723 ( 
.A1(n_1663),
.A2(n_1590),
.A3(n_1597),
.B(n_1593),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1629),
.A2(n_1567),
.B(n_1560),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1689),
.A2(n_1599),
.B1(n_1559),
.B2(n_1589),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1647),
.Y(n_1726)
);

AO31x2_ASAP7_75t_L g1727 ( 
.A1(n_1678),
.A2(n_1591),
.A3(n_1612),
.B(n_1605),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1647),
.B(n_1492),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1642),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1682),
.B(n_1482),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1668),
.Y(n_1731)
);

AO31x2_ASAP7_75t_L g1732 ( 
.A1(n_1719),
.A2(n_1631),
.A3(n_1649),
.B(n_1686),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1645),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1655),
.B(n_1646),
.Y(n_1734)
);

INVx3_ASAP7_75t_SL g1735 ( 
.A(n_1636),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1659),
.A2(n_1567),
.B(n_1560),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1665),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1669),
.A2(n_1541),
.B(n_1543),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1697),
.A2(n_1490),
.B(n_1546),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1630),
.B(n_1529),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1646),
.A2(n_1611),
.B1(n_1557),
.B2(n_1577),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1656),
.B(n_1573),
.Y(n_1742)
);

BUFx12f_ASAP7_75t_L g1743 ( 
.A(n_1639),
.Y(n_1743)
);

AO22x2_ASAP7_75t_L g1744 ( 
.A1(n_1683),
.A2(n_1497),
.B1(n_1570),
.B2(n_1498),
.Y(n_1744)
);

BUFx3_ASAP7_75t_L g1745 ( 
.A(n_1671),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_SL g1746 ( 
.A1(n_1715),
.A2(n_1628),
.B(n_1670),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1653),
.A2(n_1567),
.B(n_1575),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1650),
.A2(n_1614),
.B(n_1551),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1657),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1662),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1637),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1681),
.B(n_1493),
.Y(n_1752)
);

A2O1A1Ixp33_ASAP7_75t_L g1753 ( 
.A1(n_1666),
.A2(n_1580),
.B(n_1491),
.C(n_1532),
.Y(n_1753)
);

AO31x2_ASAP7_75t_L g1754 ( 
.A1(n_1667),
.A2(n_1609),
.A3(n_1603),
.B(n_1540),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1658),
.B(n_1497),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1637),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1713),
.B(n_1621),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1661),
.B(n_130),
.Y(n_1758)
);

AO31x2_ASAP7_75t_L g1759 ( 
.A1(n_1675),
.A2(n_1530),
.A3(n_1622),
.B(n_1574),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1660),
.A2(n_1694),
.B(n_1696),
.Y(n_1760)
);

INVx3_ASAP7_75t_SL g1761 ( 
.A(n_1680),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1635),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1684),
.A2(n_1490),
.B(n_1552),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1643),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1701),
.B(n_1528),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1688),
.A2(n_1579),
.B(n_1524),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1714),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1707),
.B(n_1542),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1749),
.A2(n_1734),
.B1(n_1726),
.B2(n_1731),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1729),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1741),
.A2(n_1710),
.B1(n_1691),
.B2(n_1654),
.Y(n_1771)
);

AND2x4_ASAP7_75t_SL g1772 ( 
.A(n_1755),
.B(n_1680),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1729),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1761),
.B(n_1627),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1746),
.A2(n_1664),
.B1(n_1712),
.B2(n_1676),
.Y(n_1775)
);

INVxp67_ASAP7_75t_L g1776 ( 
.A(n_1745),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1731),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

INVx6_ASAP7_75t_L g1779 ( 
.A(n_1743),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1735),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1751),
.Y(n_1781)
);

BUFx2_ASAP7_75t_L g1782 ( 
.A(n_1756),
.Y(n_1782)
);

CKINVDCx11_ASAP7_75t_R g1783 ( 
.A(n_1737),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1752),
.A2(n_1673),
.B1(n_1664),
.B2(n_1705),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1725),
.A2(n_1701),
.B1(n_1690),
.B2(n_1692),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1755),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1728),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1762),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1762),
.Y(n_1789)
);

AOI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1765),
.A2(n_1672),
.B(n_1709),
.Y(n_1790)
);

INVx6_ASAP7_75t_L g1791 ( 
.A(n_1758),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1750),
.A2(n_1717),
.B1(n_1634),
.B2(n_1704),
.Y(n_1792)
);

CKINVDCx11_ASAP7_75t_R g1793 ( 
.A(n_1764),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1733),
.Y(n_1794)
);

BUFx10_ASAP7_75t_L g1795 ( 
.A(n_1740),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1733),
.B(n_1658),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1722),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1757),
.A2(n_1717),
.B1(n_1651),
.B2(n_1695),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1768),
.B(n_1693),
.Y(n_1799)
);

INVx8_ASAP7_75t_L g1800 ( 
.A(n_1730),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1744),
.A2(n_1698),
.B1(n_1687),
.B2(n_1648),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1744),
.A2(n_1702),
.B1(n_1677),
.B2(n_1716),
.Y(n_1802)
);

INVx5_ASAP7_75t_L g1803 ( 
.A(n_1781),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1788),
.B(n_1742),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1770),
.Y(n_1805)
);

AO21x2_ASAP7_75t_L g1806 ( 
.A1(n_1790),
.A2(n_1748),
.B(n_1763),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_SL g1807 ( 
.A(n_1769),
.B(n_1708),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1773),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1777),
.Y(n_1809)
);

NAND2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1781),
.B(n_1708),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1782),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1787),
.Y(n_1812)
);

OAI21x1_ASAP7_75t_L g1813 ( 
.A1(n_1801),
.A2(n_1739),
.B(n_1766),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1789),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1778),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1794),
.A2(n_1747),
.B(n_1738),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1797),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1799),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1800),
.B(n_1769),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1792),
.B(n_1711),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1793),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1800),
.B(n_1699),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1800),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1794),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1796),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1792),
.B(n_1798),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1791),
.Y(n_1827)
);

OR2x6_ASAP7_75t_L g1828 ( 
.A(n_1786),
.B(n_1724),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1796),
.B(n_1732),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1802),
.B(n_1732),
.Y(n_1830)
);

AO21x2_ASAP7_75t_L g1831 ( 
.A1(n_1784),
.A2(n_1760),
.B(n_1753),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1721),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1803),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1818),
.B(n_1817),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1832),
.B(n_1772),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1805),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1826),
.A2(n_1791),
.B1(n_1798),
.B2(n_1795),
.Y(n_1837)
);

AND2x4_ASAP7_75t_SL g1838 ( 
.A(n_1827),
.B(n_1795),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1832),
.B(n_1776),
.Y(n_1839)
);

AND2x4_ASAP7_75t_L g1840 ( 
.A(n_1832),
.B(n_1784),
.Y(n_1840)
);

A2O1A1Ixp33_ASAP7_75t_L g1841 ( 
.A1(n_1826),
.A2(n_1774),
.B(n_1785),
.C(n_1771),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1812),
.Y(n_1842)
);

OAI21x1_ASAP7_75t_SL g1843 ( 
.A1(n_1807),
.A2(n_1819),
.B(n_1804),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_SL g1844 ( 
.A(n_1803),
.B(n_1638),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1820),
.A2(n_1720),
.B(n_1780),
.C(n_1640),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1825),
.B(n_1815),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1825),
.B(n_1779),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1809),
.B(n_1700),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1822),
.B(n_1779),
.Y(n_1850)
);

A2O1A1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1820),
.A2(n_1677),
.B(n_1641),
.C(n_1685),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1821),
.A2(n_1703),
.B(n_1706),
.C(n_1718),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1814),
.B(n_1783),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1823),
.A2(n_1644),
.B(n_1632),
.C(n_1652),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1808),
.B(n_1721),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_L g1856 ( 
.A1(n_1830),
.A2(n_1736),
.B(n_1531),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1833),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1855),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1840),
.B(n_1829),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1842),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1847),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1836),
.B(n_1808),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1840),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1839),
.B(n_1829),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1839),
.B(n_1824),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1833),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1848),
.B(n_1830),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1853),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1833),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1835),
.B(n_1813),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1837),
.A2(n_1831),
.B1(n_1828),
.B2(n_1803),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1843),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1869),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1862),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1869),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1862),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1858),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1858),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1861),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1870),
.B(n_1835),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1870),
.B(n_1844),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1861),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1861),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1863),
.B(n_1831),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1871),
.A2(n_1841),
.B1(n_1851),
.B2(n_1845),
.C(n_1852),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1869),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1860),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1857),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1867),
.B(n_1831),
.Y(n_1889)
);

INVx6_ASAP7_75t_L g1890 ( 
.A(n_1886),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1888),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1888),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1881),
.B(n_1872),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1880),
.B(n_1867),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1877),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1895),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1893),
.B(n_1880),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1891),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1891),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1892),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1900),
.B(n_1896),
.Y(n_1901)
);

INVxp33_ASAP7_75t_L g1902 ( 
.A(n_1897),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1898),
.B(n_1893),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1903),
.B(n_1893),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1901),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1902),
.B(n_1898),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1901),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1901),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1905),
.B(n_1899),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1907),
.A2(n_1885),
.B1(n_1890),
.B2(n_1881),
.Y(n_1910)
);

NAND3xp33_ASAP7_75t_L g1911 ( 
.A(n_1906),
.B(n_1872),
.C(n_1887),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1908),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1889),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1906),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1905),
.A2(n_1889),
.B1(n_1884),
.B2(n_1881),
.C(n_1878),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1914),
.B(n_1868),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1912),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1910),
.B(n_1878),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1909),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1911),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1913),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1915),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1914),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_SL g1924 ( 
.A1(n_1914),
.A2(n_1535),
.B1(n_1863),
.B2(n_1869),
.C1(n_1876),
.C2(n_1866),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1914),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

INVxp67_ASAP7_75t_SL g1927 ( 
.A(n_1914),
.Y(n_1927)
);

NAND3xp33_ASAP7_75t_SL g1928 ( 
.A(n_1926),
.B(n_1846),
.C(n_1894),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1925),
.B(n_1880),
.Y(n_1929)
);

NOR3xp33_ASAP7_75t_L g1930 ( 
.A(n_1927),
.B(n_1875),
.C(n_1873),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1916),
.B(n_1922),
.Y(n_1931)
);

NAND3xp33_ASAP7_75t_SL g1932 ( 
.A(n_1923),
.B(n_1866),
.C(n_1849),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1922),
.B(n_1890),
.Y(n_1933)
);

NOR2xp67_ASAP7_75t_L g1934 ( 
.A(n_1920),
.B(n_1873),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_L g1935 ( 
.A(n_1917),
.B(n_1875),
.C(n_1539),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1921),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1919),
.B(n_1890),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1918),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1924),
.B(n_1876),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1925),
.B(n_1874),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1927),
.Y(n_1941)
);

O2A1O1Ixp33_ASAP7_75t_L g1942 ( 
.A1(n_1927),
.A2(n_1850),
.B(n_1886),
.C(n_1883),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1927),
.Y(n_1943)
);

O2A1O1Ixp33_ASAP7_75t_L g1944 ( 
.A1(n_1941),
.A2(n_1850),
.B(n_1854),
.C(n_1874),
.Y(n_1944)
);

AOI21xp33_ASAP7_75t_SL g1945 ( 
.A1(n_1931),
.A2(n_1879),
.B(n_1882),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1937),
.Y(n_1946)
);

AOI221x1_ASAP7_75t_L g1947 ( 
.A1(n_1943),
.A2(n_1882),
.B1(n_1870),
.B2(n_1856),
.C(n_1859),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1933),
.A2(n_1870),
.B(n_1859),
.Y(n_1948)
);

NAND5xp2_ASAP7_75t_L g1949 ( 
.A(n_1938),
.B(n_1942),
.C(n_1939),
.D(n_1930),
.E(n_1935),
.Y(n_1949)
);

AOI32xp33_ASAP7_75t_L g1950 ( 
.A1(n_1936),
.A2(n_1838),
.A3(n_1859),
.B1(n_1865),
.B2(n_1864),
.Y(n_1950)
);

OAI211xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1929),
.A2(n_1844),
.B(n_226),
.C(n_228),
.Y(n_1951)
);

AOI222xp33_ASAP7_75t_L g1952 ( 
.A1(n_1934),
.A2(n_1859),
.B1(n_1865),
.B2(n_1864),
.C1(n_1803),
.C2(n_1813),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1940),
.B(n_1806),
.Y(n_1953)
);

NOR3xp33_ASAP7_75t_L g1954 ( 
.A(n_1932),
.B(n_1487),
.C(n_1554),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1928),
.A2(n_1708),
.B(n_1816),
.C(n_1527),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1933),
.A2(n_1806),
.B1(n_1810),
.B2(n_1828),
.C(n_1723),
.Y(n_1956)
);

AOI21xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1931),
.A2(n_225),
.B(n_229),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1937),
.Y(n_1958)
);

OAI211xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1941),
.A2(n_230),
.B(n_231),
.C(n_236),
.Y(n_1959)
);

OAI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1931),
.A2(n_1816),
.B(n_240),
.C(n_242),
.Y(n_1960)
);

AOI222xp33_ASAP7_75t_L g1961 ( 
.A1(n_1946),
.A2(n_1806),
.B1(n_1810),
.B2(n_1723),
.C1(n_1828),
.C2(n_1727),
.Y(n_1961)
);

NAND4xp25_ASAP7_75t_L g1962 ( 
.A(n_1949),
.B(n_239),
.C(n_243),
.D(n_244),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1958),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1953),
.Y(n_1964)
);

AND3x1_ASAP7_75t_L g1965 ( 
.A(n_1944),
.B(n_1828),
.C(n_245),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1955),
.B(n_246),
.Y(n_1966)
);

AOI221xp5_ASAP7_75t_L g1967 ( 
.A1(n_1957),
.A2(n_1723),
.B1(n_1727),
.B2(n_1721),
.C(n_251),
.Y(n_1967)
);

NAND2x1p5_ASAP7_75t_L g1968 ( 
.A(n_1959),
.B(n_247),
.Y(n_1968)
);

XNOR2xp5_ASAP7_75t_L g1969 ( 
.A(n_1960),
.B(n_249),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1948),
.A2(n_1732),
.B1(n_1727),
.B2(n_1759),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1945),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.C(n_254),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_SL g1972 ( 
.A(n_1954),
.B(n_256),
.Y(n_1972)
);

O2A1O1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1951),
.A2(n_260),
.B(n_261),
.C(n_263),
.Y(n_1973)
);

AOI222xp33_ASAP7_75t_L g1974 ( 
.A1(n_1956),
.A2(n_265),
.B1(n_267),
.B2(n_269),
.C1(n_270),
.C2(n_271),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1950),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1947),
.Y(n_1976)
);

AOI222xp33_ASAP7_75t_L g1977 ( 
.A1(n_1952),
.A2(n_272),
.B1(n_273),
.B2(n_277),
.C1(n_280),
.C2(n_285),
.Y(n_1977)
);

OAI221xp5_ASAP7_75t_SL g1978 ( 
.A1(n_1958),
.A2(n_1759),
.B1(n_289),
.B2(n_292),
.C(n_298),
.Y(n_1978)
);

OAI211xp5_ASAP7_75t_L g1979 ( 
.A1(n_1958),
.A2(n_286),
.B(n_299),
.C(n_301),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1963),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1976),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1975),
.A2(n_1759),
.B1(n_1754),
.B2(n_305),
.Y(n_1982)
);

INVxp67_ASAP7_75t_SL g1983 ( 
.A(n_1968),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1965),
.B(n_302),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1969),
.B(n_303),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1962),
.B(n_309),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1964),
.Y(n_1987)
);

AOI31xp33_ASAP7_75t_L g1988 ( 
.A1(n_1971),
.A2(n_314),
.A3(n_315),
.B(n_316),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_L g1989 ( 
.A(n_1974),
.B(n_318),
.C(n_319),
.Y(n_1989)
);

AO22x2_ASAP7_75t_L g1990 ( 
.A1(n_1979),
.A2(n_323),
.B1(n_324),
.B2(n_326),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1966),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1980),
.B(n_1964),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1983),
.B(n_1987),
.Y(n_1993)
);

O2A1O1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1981),
.A2(n_1972),
.B(n_1973),
.C(n_1977),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1986),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1990),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1984),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1991),
.A2(n_1978),
.B1(n_1967),
.B2(n_1970),
.C(n_1961),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1985),
.A2(n_1754),
.B1(n_334),
.B2(n_336),
.Y(n_1999)
);

NAND3x1_ASAP7_75t_L g2000 ( 
.A(n_1989),
.B(n_327),
.C(n_337),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_1982),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_L g2002 ( 
.A(n_1993),
.B(n_1988),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1995),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1992),
.A2(n_339),
.B(n_340),
.Y(n_2004)
);

AND3x1_ASAP7_75t_L g2005 ( 
.A(n_1994),
.B(n_343),
.C(n_346),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1997),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_2001),
.A2(n_1754),
.B1(n_351),
.B2(n_352),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1996),
.B(n_347),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1999),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2003),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2002),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2006),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_2005),
.A2(n_2000),
.B1(n_1998),
.B2(n_358),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_SL g2014 ( 
.A(n_2012),
.B(n_2008),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2010),
.Y(n_2015)
);

OAI22xp5_ASAP7_75t_SL g2016 ( 
.A1(n_2013),
.A2(n_2009),
.B1(n_2007),
.B2(n_2004),
.Y(n_2016)
);

OAI22x1_ASAP7_75t_L g2017 ( 
.A1(n_2015),
.A2(n_2011),
.B1(n_357),
.B2(n_360),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2014),
.B(n_355),
.Y(n_2018)
);

XNOR2xp5_ASAP7_75t_L g2019 ( 
.A(n_2017),
.B(n_2016),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2018),
.B(n_362),
.C(n_364),
.Y(n_2020)
);

OAI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_2018),
.A2(n_368),
.B(n_369),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_2019),
.A2(n_2021),
.B(n_2020),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2019),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_2023),
.B(n_370),
.Y(n_2024)
);

OAI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_2024),
.A2(n_2022),
.B1(n_373),
.B2(n_376),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_2025),
.A2(n_371),
.B1(n_380),
.B2(n_381),
.C(n_385),
.Y(n_2026)
);

AOI211xp5_ASAP7_75t_L g2027 ( 
.A1(n_2026),
.A2(n_386),
.B(n_387),
.C(n_390),
.Y(n_2027)
);


endmodule