module fake_jpeg_3042_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_23),
.A2(n_7),
.B(n_11),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_2),
.B(n_3),
.Y(n_97)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_19),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_63),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_4),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_61),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_30),
.B(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_69),
.Y(n_88)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_65),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_9),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_30),
.B(n_8),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_8),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_27),
.B1(n_14),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_75),
.B1(n_79),
.B2(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_69),
.B1(n_67),
.B2(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_27),
.B1(n_14),
.B2(n_26),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_26),
.B1(n_15),
.B2(n_33),
.Y(n_82)
);

NAND2x1_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_15),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_38),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_35),
.B1(n_28),
.B2(n_18),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_57),
.B1(n_43),
.B2(n_35),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_36),
.B1(n_24),
.B2(n_0),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_36),
.B1(n_1),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_12),
.B1(n_103),
.B2(n_89),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_37),
.B(n_1),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_60),
.A2(n_2),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_114),
.Y(n_135)
);

INVx2_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_12),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_92),
.B1(n_102),
.B2(n_70),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_98),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_108),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_95),
.C(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_93),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_137),
.B(n_139),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_73),
.B(n_82),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_129),
.B(n_152),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_70),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_132),
.B1(n_134),
.B2(n_121),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_79),
.B1(n_96),
.B2(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_96),
.B1(n_94),
.B2(n_72),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_90),
.C(n_71),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_125),
.C(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_131),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_160),
.B(n_168),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_125),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_172),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_167),
.B1(n_149),
.B2(n_151),
.Y(n_173)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_151),
.A2(n_122),
.B1(n_125),
.B2(n_128),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_111),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_142),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_184),
.B1(n_165),
.B2(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_149),
.C(n_155),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_181),
.C(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_139),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_137),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_110),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_114),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_140),
.B1(n_138),
.B2(n_136),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_164),
.B1(n_157),
.B2(n_168),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_144),
.B1(n_128),
.B2(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_191),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_195),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_158),
.A3(n_168),
.B1(n_163),
.B2(n_160),
.Y(n_190)
);

OAI322xp33_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_135),
.A3(n_161),
.B1(n_160),
.B2(n_159),
.C1(n_111),
.C2(n_145),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_135),
.A3(n_161),
.B1(n_166),
.B2(n_120),
.C(n_124),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_162),
.B1(n_143),
.B2(n_133),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_148),
.C(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_198),
.C(n_192),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_130),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_205),
.C(n_198),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_201),
.B(n_175),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_181),
.C(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_200),
.A2(n_189),
.B1(n_184),
.B2(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_213),
.B1(n_200),
.B2(n_202),
.Y(n_214)
);

OA21x2_ASAP7_75t_SL g211 ( 
.A1(n_204),
.A2(n_190),
.B(n_186),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_212),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_203),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_217),
.B1(n_209),
.B2(n_210),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_209),
.C(n_211),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_205),
.B1(n_175),
.B2(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_215),
.A2(n_207),
.B1(n_213),
.B2(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_218),
.B(n_214),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_216),
.C(n_217),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_222),
.B1(n_219),
.B2(n_210),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_72),
.A3(n_143),
.B1(n_153),
.B2(n_176),
.C1(n_224),
.C2(n_218),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_227),
.CI(n_176),
.CON(n_230),
.SN(n_230)
);


endmodule