module real_jpeg_33636_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_1),
.B(n_37),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_1),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_1),
.B(n_163),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_2),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_4),
.B(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_5),
.Y(n_113)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_6),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_6),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_11),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_12),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_13),
.B(n_37),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_136),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_100),
.B(n_135),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_72),
.B(n_99),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_54),
.B(n_71),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_21),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_21),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_43),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_44),
.C(n_49),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_35),
.B(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_37),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_39),
.B(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_45),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_64),
.B(n_70),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_74),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_88),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_89),
.C(n_92),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_85),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.C(n_85),
.Y(n_121)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_96),
.B(n_162),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_102),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_122),
.B1(n_133),
.B2(n_134),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_120),
.B2(n_121),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_121),
.C(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_114),
.C(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_125),
.C(n_129),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_186),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_185),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_185),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_169),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_156),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_152),
.B2(n_155),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_152),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_165),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);


endmodule