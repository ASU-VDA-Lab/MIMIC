module fake_jpeg_10332_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_17),
.B1(n_24),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_65),
.B1(n_34),
.B2(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_57),
.Y(n_70)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_22),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_17),
.B1(n_24),
.B2(n_20),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_52),
.A2(n_23),
.B1(n_21),
.B2(n_29),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_33),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_19),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_17),
.B1(n_20),
.B2(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_27),
.Y(n_90)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_68),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_17),
.B1(n_34),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_83),
.B1(n_100),
.B2(n_59),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_79),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_78),
.B(n_33),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_31),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_30),
.B1(n_60),
.B2(n_58),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_22),
.B1(n_43),
.B2(n_38),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_103),
.B1(n_61),
.B2(n_45),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_31),
.B1(n_34),
.B2(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_28),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_97),
.B1(n_61),
.B2(n_45),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_33),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_27),
.B1(n_28),
.B2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_39),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_101),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_105),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_65),
.C(n_48),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_59),
.B(n_33),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_25),
.C(n_19),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_113),
.Y(n_147)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_101),
.B1(n_70),
.B2(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_119),
.A2(n_70),
.B1(n_75),
.B2(n_69),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_129),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_75),
.B1(n_69),
.B2(n_84),
.Y(n_143)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_92),
.Y(n_135)
);

OAI22x1_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_86),
.B1(n_68),
.B2(n_67),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_132),
.B(n_138),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_111),
.B1(n_159),
.B2(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_152),
.C(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_124),
.B1(n_126),
.B2(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_151),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_84),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_161),
.B(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_77),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_148),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_89),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_99),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_98),
.C(n_102),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_91),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_104),
.B1(n_116),
.B2(n_107),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_121),
.B1(n_106),
.B2(n_113),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_93),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_48),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_157),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_96),
.B1(n_81),
.B2(n_103),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_25),
.B1(n_19),
.B2(n_43),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_0),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_168),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_142),
.A3(n_141),
.B1(n_151),
.B2(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_105),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_170),
.B1(n_180),
.B2(n_185),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_129),
.B1(n_110),
.B2(n_127),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_174),
.A2(n_187),
.B1(n_188),
.B2(n_2),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_178),
.B(n_183),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_179),
.A2(n_161),
.B(n_136),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_186),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_111),
.B1(n_25),
.B2(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_55),
.B1(n_25),
.B2(n_3),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_55),
.B1(n_2),
.B2(n_4),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_1),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_198),
.C(n_199),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_152),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_148),
.C(n_145),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_211),
.B1(n_175),
.B2(n_178),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_132),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_208),
.C(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_139),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_187),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_2),
.C(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_5),
.C(n_7),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_177),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_172),
.B(n_168),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_170),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_164),
.B1(n_175),
.B2(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_232),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_220),
.B(n_227),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_169),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_9),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_180),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_231),
.C(n_233),
.Y(n_235)
);

OA21x2_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_194),
.B(n_199),
.Y(n_227)
);

OR2x6_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_174),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_229),
.A2(n_193),
.B(n_201),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_181),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_211),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_197),
.C(n_202),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_247),
.C(n_228),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_183),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_243),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_241),
.A2(n_250),
.B(n_222),
.C(n_224),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_225),
.A2(n_193),
.B(n_182),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_244),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_200),
.B(n_201),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_173),
.B(n_212),
.Y(n_245)
);

HAxp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_248),
.CON(n_262),
.SN(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_210),
.C(n_8),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_226),
.A2(n_7),
.B(n_8),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_8),
.B(n_9),
.Y(n_249)
);

AOI21x1_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_11),
.B(n_12),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_219),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_215),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_228),
.C(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_259),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_233),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_263),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_10),
.C(n_11),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_11),
.B(n_12),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_248),
.B(n_245),
.Y(n_264)
);

AOI31xp67_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_262),
.A3(n_249),
.B(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_271),
.Y(n_276)
);

XOR2x1_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_246),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_241),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_246),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_273),
.A2(n_261),
.B(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_255),
.B(n_256),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_251),
.B(n_254),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_268),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_267),
.A2(n_247),
.B1(n_14),
.B2(n_15),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.C(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_274),
.B(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_276),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_289),
.B(n_290),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_13),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_279),
.B(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_13),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_16),
.B(n_292),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_16),
.Y(n_294)
);


endmodule