module fake_jpeg_20881_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_32),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_64),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_50),
.B(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_24),
.B1(n_29),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_19),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_40),
.B1(n_38),
.B2(n_18),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_74),
.B(n_85),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_94),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_84),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_97),
.B1(n_21),
.B2(n_26),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_39),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_40),
.B1(n_41),
.B2(n_37),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_17),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_17),
.B1(n_43),
.B2(n_40),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_25),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_98),
.B1(n_35),
.B2(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_26),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_106),
.B(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_80),
.B1(n_75),
.B2(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_101),
.B(n_30),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2x1_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_37),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_37),
.B1(n_35),
.B2(n_38),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_118),
.B1(n_71),
.B2(n_93),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_1),
.B(n_2),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_21),
.B(n_31),
.Y(n_114)
);

NOR2xp67_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_32),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_96),
.B1(n_66),
.B2(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_76),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_125),
.B(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_137),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_86),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_28),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_132),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_86),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_143),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_142),
.Y(n_168)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_100),
.B1(n_99),
.B2(n_114),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_150),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_115),
.B1(n_80),
.B2(n_79),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_94),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_28),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_15),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_124),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_152),
.B(n_146),
.Y(n_175)
);

OAI21x1_ASAP7_75t_R g153 ( 
.A1(n_129),
.A2(n_117),
.B(n_110),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_69),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_124),
.A3(n_103),
.B1(n_123),
.B2(n_110),
.C1(n_67),
.C2(n_90),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_30),
.B1(n_27),
.B2(n_140),
.C(n_75),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_123),
.C(n_70),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_30),
.C(n_27),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_103),
.B1(n_119),
.B2(n_89),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_136),
.B1(n_133),
.B2(n_139),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_167),
.A2(n_32),
.B(n_115),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_143),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_127),
.B1(n_126),
.B2(n_133),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_187),
.B1(n_171),
.B2(n_157),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_182),
.B1(n_184),
.B2(n_170),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_152),
.B(n_150),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_191),
.C(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_192),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_139),
.B1(n_143),
.B2(n_136),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_183),
.A2(n_185),
.B(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_140),
.B1(n_142),
.B2(n_98),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_161),
.B(n_165),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_69),
.B1(n_75),
.B2(n_15),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_14),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_205),
.B1(n_174),
.B2(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_203),
.B1(n_206),
.B2(n_178),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_202),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_182),
.B1(n_177),
.B2(n_155),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_2),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_168),
.B1(n_172),
.B2(n_166),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_151),
.B1(n_158),
.B2(n_172),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_196),
.B(n_175),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_215),
.C(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_193),
.B(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_214),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_183),
.C(n_181),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_210),
.B1(n_198),
.B2(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_13),
.C(n_12),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_203),
.C(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_3),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_201),
.B1(n_207),
.B2(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_207),
.B1(n_198),
.B2(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_216),
.B(n_227),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_234),
.B1(n_228),
.B2(n_220),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_217),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_222),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_237),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_222),
.B(n_225),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_238),
.B(n_234),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_223),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_7),
.C(n_8),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_239),
.B(n_8),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_245),
.A2(n_243),
.B(n_9),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_7),
.Y(n_247)
);


endmodule