module real_jpeg_28312_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_1),
.A2(n_10),
.B(n_92),
.C(n_94),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_42),
.B1(n_94),
.B2(n_95),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_66),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_66),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_5),
.A2(n_37),
.B1(n_94),
.B2(n_95),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_7),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_9),
.B(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_29),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_10),
.A2(n_29),
.B(n_59),
.C(n_68),
.D(n_124),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_26),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_10),
.A2(n_51),
.B(n_136),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_22),
.B(n_32),
.C(n_74),
.D(n_164),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_113)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_118),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_18),
.B(n_82),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_57),
.C(n_71),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_19),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_39),
.C(n_44),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_31),
.Y(n_20)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_23),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_22),
.A2(n_42),
.B(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_23),
.A2(n_29),
.A3(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_25),
.B(n_36),
.Y(n_164)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_26),
.A2(n_32),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_28),
.B(n_30),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g123 ( 
.A1(n_28),
.A2(n_46),
.A3(n_61),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_29),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_41),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_41),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_46),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_47),
.B(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_51),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_56),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_56),
.A2(n_87),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_57),
.B(n_71),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_67),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_59),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_69),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_70),
.A2(n_114),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_70),
.B(n_93),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_72),
.B(n_76),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_79),
.A2(n_142),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_81),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_98),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_154),
.Y(n_153)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B(n_103),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_169),
.B(n_173),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_159),
.B(n_168),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_138),
.B(n_158),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_135),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_145),
.B(n_157),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_156),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_161),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);


endmodule