module fake_jpeg_4878_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_27),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_30),
.C(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_28),
.B1(n_30),
.B2(n_25),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_28),
.B1(n_24),
.B2(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_16),
.B(n_24),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_17),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_17),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_37),
.B1(n_36),
.B2(n_39),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_74),
.B1(n_48),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_18),
.B1(n_36),
.B2(n_55),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_28),
.B1(n_38),
.B2(n_39),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_72),
.C(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_38),
.B1(n_36),
.B2(n_22),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_90),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_104),
.B(n_15),
.Y(n_135)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_101),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_45),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_77),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_54),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_18),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_59),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_60),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_65),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_63),
.C(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_107),
.B(n_73),
.Y(n_120)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_111),
.B1(n_76),
.B2(n_79),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_64),
.B1(n_55),
.B2(n_62),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_72),
.B(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_91),
.C(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_120),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_124),
.Y(n_142)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_80),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_130),
.B(n_134),
.Y(n_143)
);

INVxp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.Y(n_127)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_53),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_109),
.B1(n_103),
.B2(n_90),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_135),
.B1(n_106),
.B2(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_78),
.B1(n_70),
.B2(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_110),
.B1(n_106),
.B2(n_78),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_18),
.B(n_15),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_144),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_105),
.B1(n_97),
.B2(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_92),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_146),
.B(n_134),
.Y(n_173)
);

BUFx12f_ASAP7_75t_SL g146 ( 
.A(n_135),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_15),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_153),
.C(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_159),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_15),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_152),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_15),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_71),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_15),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_167),
.C(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_123),
.C(n_112),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_158),
.A2(n_132),
.B1(n_113),
.B2(n_122),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_169),
.B1(n_174),
.B2(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_119),
.B1(n_133),
.B2(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_155),
.B(n_128),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_113),
.B1(n_133),
.B2(n_116),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_112),
.B1(n_115),
.B2(n_61),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_23),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_154),
.B(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_26),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_116),
.B1(n_120),
.B2(n_119),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_190),
.C(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_145),
.B(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_179),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_149),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_139),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_200),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_143),
.C(n_128),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_129),
.B1(n_124),
.B2(n_37),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_201),
.B1(n_172),
.B2(n_162),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_129),
.C(n_71),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_173),
.C(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_129),
.B1(n_37),
.B2(n_29),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_181),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_208),
.B1(n_210),
.B2(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_213),
.C(n_217),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_163),
.B1(n_171),
.B2(n_177),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_214),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_178),
.B1(n_174),
.B2(n_162),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_195),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_215),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_182),
.C(n_37),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_218),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_230),
.B(n_233),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_186),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_23),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_212),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_197),
.B1(n_185),
.B2(n_199),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_224),
.B1(n_231),
.B2(n_227),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_219),
.B(n_188),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_213),
.C(n_217),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_190),
.C(n_192),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_215),
.C(n_204),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_29),
.B1(n_1),
.B2(n_0),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_20),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_238),
.C(n_240),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_229),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_222),
.Y(n_247)
);

AO221x1_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_23),
.B1(n_20),
.B2(n_0),
.C(n_1),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_242),
.B(n_245),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_10),
.C(n_14),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_23),
.C(n_20),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_5),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_0),
.B1(n_1),
.B2(n_23),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_245),
.C(n_244),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_2),
.B(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_253),
.B(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_26),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_23),
.Y(n_259)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_4),
.B(n_5),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_261),
.B1(n_6),
.B2(n_9),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_4),
.C(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_258),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_259),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_252),
.C(n_254),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_20),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_20),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_261),
.A2(n_249),
.B1(n_9),
.B2(n_10),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_265),
.B(n_11),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_263),
.B(n_266),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_269),
.B(n_11),
.C(n_13),
.D(n_14),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_6),
.B(n_11),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_13),
.C(n_26),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_272),
.B(n_271),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_20),
.Y(n_274)
);


endmodule