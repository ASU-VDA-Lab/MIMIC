module fake_jpeg_11271_n_185 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_10),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx8_ASAP7_75t_SL g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_25),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_9),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_92),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_73),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_64),
.B1(n_69),
.B2(n_60),
.Y(n_102)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_73),
.B1(n_72),
.B2(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_94),
.A2(n_106),
.B1(n_107),
.B2(n_81),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_55),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_1),
.C(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_72),
.B1(n_78),
.B2(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_70),
.B1(n_80),
.B2(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_57),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_67),
.B1(n_74),
.B2(n_79),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_67),
.B1(n_79),
.B2(n_65),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_116),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_71),
.B(n_58),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_75),
.B1(n_68),
.B2(n_56),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_124),
.B(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_76),
.B(n_3),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_119),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_126),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_29),
.B1(n_53),
.B2(n_51),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_21),
.B1(n_46),
.B2(n_45),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_19),
.B(n_48),
.C(n_47),
.Y(n_124)
);

CKINVDCx9p33_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_93),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_4),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_4),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_137),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_145),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_7),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_36),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_122),
.B(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_13),
.B(n_16),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_18),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_165),
.C(n_138),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_159),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_136),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_38),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_40),
.Y(n_161)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_162),
.A3(n_164),
.B1(n_140),
.B2(n_137),
.C1(n_135),
.C2(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_54),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_171),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_177),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_143),
.B1(n_151),
.B2(n_169),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_175),
.A2(n_169),
.B1(n_156),
.B2(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_178),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_158),
.C(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_150),
.B1(n_176),
.B2(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_157),
.Y(n_185)
);


endmodule