module fake_jpeg_1299_n_682 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_682);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_682;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_58),
.B(n_63),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_61),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_66),
.Y(n_189)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_67),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_74),
.Y(n_167)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_77),
.B(n_81),
.Y(n_175)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_79),
.B(n_111),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_37),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_82),
.B(n_90),
.Y(n_181)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_43),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_91),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_93),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_94),
.B(n_97),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_95),
.Y(n_211)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_99),
.A2(n_36),
.B1(n_48),
.B2(n_47),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_39),
.Y(n_101)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_23),
.B(n_9),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_102),
.B(n_104),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_39),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_105),
.B(n_106),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_23),
.B(n_18),
.C(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_31),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_109),
.B(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_11),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_119),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_33),
.B(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_120),
.B(n_125),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_27),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_122),
.B(n_74),
.Y(n_228)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_9),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_130),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_35),
.Y(n_129)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_28),
.Y(n_131)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_72),
.B1(n_116),
.B2(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_134),
.A2(n_149),
.B1(n_182),
.B2(n_218),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_85),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_136),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_59),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_139),
.B(n_151),
.Y(n_262)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_142),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g273 ( 
.A(n_144),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_78),
.A2(n_30),
.B1(n_51),
.B2(n_49),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_60),
.Y(n_151)
);

INVx2_ASAP7_75t_R g153 ( 
.A(n_75),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_153),
.B(n_229),
.Y(n_237)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_178),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_83),
.A2(n_36),
.B1(n_51),
.B2(n_49),
.Y(n_182)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_69),
.B(n_45),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_186),
.Y(n_259)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_190),
.Y(n_310)
);

BUFx12_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_191),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_62),
.Y(n_196)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_196),
.Y(n_318)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

CKINVDCx6p67_ASAP7_75t_R g270 ( 
.A(n_200),
.Y(n_270)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_96),
.Y(n_203)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_66),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_206),
.B(n_231),
.Y(n_282)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_73),
.Y(n_210)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_76),
.Y(n_213)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_84),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_65),
.Y(n_219)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_100),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_80),
.Y(n_227)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_38),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_92),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_238),
.Y(n_322)
);

INVx5_ASAP7_75t_SL g235 ( 
.A(n_153),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_235),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_188),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_236),
.A2(n_253),
.B1(n_271),
.B2(n_155),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_237),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_106),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_150),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_240),
.B(n_276),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_150),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_243),
.B(n_258),
.Y(n_340)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_245),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_86),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_246),
.B(n_257),
.Y(n_319)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_248),
.Y(n_326)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_249),
.Y(n_323)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_208),
.A2(n_212),
.B1(n_215),
.B2(n_193),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_186),
.A2(n_45),
.B1(n_39),
.B2(n_44),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_143),
.B(n_0),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_175),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_175),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_261),
.B(n_265),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_184),
.B(n_103),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

CKINVDCx12_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_186),
.A2(n_98),
.B1(n_95),
.B2(n_93),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_195),
.B(n_16),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_181),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_289),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_181),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_173),
.B(n_0),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_0),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_224),
.B(n_16),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_294),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_183),
.A2(n_99),
.B1(n_45),
.B2(n_44),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_285),
.A2(n_296),
.B1(n_311),
.B2(n_227),
.Y(n_362)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_176),
.Y(n_287)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_187),
.Y(n_288)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_145),
.B(n_15),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_137),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_147),
.B(n_15),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_292),
.B(n_298),
.Y(n_363)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_141),
.Y(n_293)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_157),
.B(n_209),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_140),
.Y(n_295)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_149),
.A2(n_45),
.B1(n_44),
.B2(n_52),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_52),
.C(n_42),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_137),
.C(n_207),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_180),
.B(n_205),
.Y(n_298)
);

BUFx16f_ASAP7_75t_L g299 ( 
.A(n_230),
.Y(n_299)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_205),
.B(n_14),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_300),
.B(n_301),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_132),
.B(n_14),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_156),
.Y(n_304)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_133),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_305),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_219),
.A2(n_44),
.B1(n_42),
.B2(n_52),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_306),
.A2(n_314),
.B1(n_160),
.B2(n_194),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_148),
.B(n_7),
.Y(n_307)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_182),
.A2(n_42),
.B1(n_34),
.B2(n_27),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_138),
.B(n_6),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_312),
.B(n_315),
.Y(n_343)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_198),
.Y(n_313)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_163),
.A2(n_34),
.B1(n_2),
.B2(n_3),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_152),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_217),
.B(n_169),
.Y(n_316)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_174),
.B(n_6),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_317),
.A2(n_146),
.B1(n_192),
.B2(n_189),
.Y(n_348)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_259),
.A2(n_134),
.B(n_191),
.C(n_230),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g425 ( 
.A1(n_324),
.A2(n_362),
.B1(n_232),
.B2(n_242),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_246),
.B(n_152),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_325),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_204),
.B(n_216),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_333),
.A2(n_372),
.B1(n_379),
.B2(n_299),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_267),
.A2(n_225),
.B1(n_189),
.B2(n_222),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_334),
.A2(n_368),
.B1(n_270),
.B2(n_263),
.Y(n_416)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_337),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_348),
.B(n_299),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_257),
.B(n_281),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_364),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_358),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_271),
.A2(n_198),
.B1(n_155),
.B2(n_222),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_354),
.A2(n_270),
.B1(n_249),
.B2(n_250),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_258),
.A2(n_159),
.B1(n_146),
.B2(n_211),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_359),
.Y(n_419)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

A2O1A1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_280),
.A2(n_204),
.B(n_216),
.C(n_172),
.Y(n_361)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_365),
.B(n_378),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_309),
.B(n_262),
.Y(n_364)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_263),
.Y(n_366)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_237),
.A2(n_159),
.B1(n_207),
.B2(n_201),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_254),
.B(n_203),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_296),
.A2(n_196),
.B1(n_179),
.B2(n_164),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_247),
.Y(n_374)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_374),
.Y(n_407)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_248),
.Y(n_376)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_285),
.A2(n_172),
.B(n_34),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_311),
.A2(n_211),
.B1(n_201),
.B2(n_192),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_319),
.B(n_297),
.C(n_288),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_381),
.B(n_418),
.C(n_342),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_244),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_SL g455 ( 
.A(n_382),
.B(n_420),
.C(n_424),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_244),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_385),
.A2(n_387),
.B(n_425),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_329),
.A2(n_304),
.B1(n_254),
.B2(n_303),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_386),
.A2(n_414),
.B1(n_423),
.B2(n_427),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_282),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_392),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_234),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_399),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_319),
.B(n_350),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_398),
.Y(n_432)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

OR2x4_ASAP7_75t_L g397 ( 
.A(n_356),
.B(n_235),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_SL g457 ( 
.A1(n_397),
.A2(n_371),
.B(n_343),
.C(n_353),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_309),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_286),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_274),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_400),
.B(n_409),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_340),
.B(n_303),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_408),
.B(n_412),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_274),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_336),
.B(n_287),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_349),
.B(n_268),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_413),
.B(n_417),
.Y(n_436)
);

INVx5_ASAP7_75t_SL g415 ( 
.A(n_331),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_415),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_347),
.B(n_290),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_339),
.B(n_273),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_270),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_344),
.A2(n_232),
.B1(n_242),
.B2(n_266),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_422),
.A2(n_255),
.B(n_371),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_362),
.A2(n_290),
.B1(n_252),
.B2(n_239),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_324),
.B(n_270),
.Y(n_424)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_378),
.A2(n_252),
.B1(n_239),
.B2(n_241),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_266),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_428),
.B(n_353),
.Y(n_462)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_332),
.Y(n_429)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_429),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_395),
.Y(n_433)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_429),
.Y(n_437)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_390),
.A2(n_325),
.B1(n_328),
.B2(n_358),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_446),
.B1(n_468),
.B2(n_406),
.Y(n_473)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_441),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_394),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_453),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_391),
.A2(n_339),
.B(n_325),
.C(n_361),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_447),
.B(n_448),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_390),
.A2(n_365),
.B1(n_348),
.B2(n_328),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_324),
.B(n_331),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_383),
.A2(n_332),
.B(n_341),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_408),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g495 ( 
.A(n_449),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_343),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_457),
.B(n_463),
.Y(n_482)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_406),
.A2(n_341),
.B1(n_354),
.B2(n_337),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

INVx5_ASAP7_75t_SL g474 ( 
.A(n_460),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_374),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_462),
.B(n_323),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_398),
.B(n_342),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_407),
.Y(n_466)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_417),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_470),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_401),
.A2(n_336),
.B1(n_335),
.B2(n_320),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_424),
.A2(n_255),
.B(n_245),
.Y(n_470)
);

BUFx24_ASAP7_75t_SL g471 ( 
.A(n_382),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_381),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_462),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_472),
.B(n_480),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_473),
.A2(n_494),
.B1(n_499),
.B2(n_504),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_443),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_491),
.Y(n_515)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_479),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_335),
.C(n_425),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_487),
.C(n_488),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_485),
.B(n_496),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_411),
.Y(n_486)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_486),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_425),
.C(n_376),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_446),
.A2(n_406),
.B1(n_423),
.B2(n_427),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_430),
.B1(n_457),
.B2(n_436),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_445),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_442),
.B(n_425),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_507),
.C(n_448),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_465),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_493),
.B(n_430),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_459),
.A2(n_420),
.B1(n_414),
.B2(n_422),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_338),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_405),
.Y(n_498)
);

AOI21xp33_ASAP7_75t_L g513 ( 
.A1(n_498),
.A2(n_468),
.B(n_447),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_451),
.A2(n_386),
.B1(n_402),
.B2(n_421),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_402),
.Y(n_500)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_500),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_456),
.A2(n_402),
.B1(n_403),
.B2(n_405),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_467),
.B(n_403),
.Y(n_505)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_505),
.Y(n_527)
);

MAJx2_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_415),
.C(n_323),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_457),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_367),
.C(n_327),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_388),
.Y(n_508)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_508),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_456),
.A2(n_388),
.B1(n_419),
.B2(n_359),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_511),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_470),
.A2(n_419),
.B1(n_330),
.B2(n_410),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_495),
.B(n_486),
.Y(n_512)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_513),
.A2(n_474),
.B(n_497),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_518),
.A2(n_521),
.B1(n_535),
.B2(n_511),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_519),
.B(n_532),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_477),
.A2(n_440),
.B1(n_464),
.B2(n_433),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_487),
.A2(n_455),
.B1(n_444),
.B2(n_431),
.Y(n_522)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_522),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_524),
.B(n_529),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_525),
.B(n_503),
.Y(n_576)
);

NOR4xp25_ASAP7_75t_L g526 ( 
.A(n_478),
.B(n_457),
.C(n_437),
.D(n_435),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g568 ( 
.A(n_526),
.B(n_499),
.CI(n_510),
.CON(n_568),
.SN(n_568)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_476),
.B(n_438),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_488),
.B(n_435),
.C(n_466),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_537),
.C(n_540),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_457),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_543),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_458),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_375),
.Y(n_533)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_508),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_534),
.B(n_484),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_494),
.A2(n_452),
.B1(n_460),
.B2(n_454),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_481),
.B(n_469),
.C(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_538),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_507),
.B(n_434),
.C(n_327),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_483),
.B(n_352),
.Y(n_541)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_541),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_482),
.C(n_492),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_475),
.C(n_509),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_473),
.A2(n_434),
.B1(n_452),
.B2(n_450),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_490),
.A2(n_450),
.B1(n_330),
.B2(n_389),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_548),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_482),
.B(n_404),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_546),
.B(n_502),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_352),
.Y(n_547)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_547),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_505),
.A2(n_502),
.B1(n_489),
.B2(n_509),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_475),
.B(n_404),
.Y(n_549)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_549),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_551),
.A2(n_539),
.B1(n_515),
.B2(n_527),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_526),
.A2(n_501),
.B(n_504),
.Y(n_552)
);

XOR2x1_ASAP7_75t_L g605 ( 
.A(n_552),
.B(n_273),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_530),
.Y(n_554)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_554),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_557),
.B(n_562),
.Y(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_563),
.A2(n_527),
.B1(n_523),
.B2(n_538),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_536),
.A2(n_474),
.B1(n_497),
.B2(n_489),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_564),
.A2(n_580),
.B1(n_545),
.B2(n_543),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_514),
.B(n_479),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_568),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_516),
.B(n_484),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_578),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_544),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_570),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_516),
.B(n_268),
.C(n_426),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_572),
.B(n_574),
.C(n_577),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_389),
.C(n_503),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g597 ( 
.A(n_576),
.B(n_548),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_540),
.B(n_519),
.C(n_542),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_518),
.B(n_321),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_512),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_579),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_536),
.A2(n_370),
.B1(n_360),
.B2(n_346),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_546),
.C(n_522),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_589),
.C(n_591),
.Y(n_607)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_584),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_564),
.A2(n_556),
.B1(n_565),
.B2(n_555),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_585),
.A2(n_598),
.B1(n_604),
.B2(n_562),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_586),
.A2(n_585),
.B(n_584),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_587),
.A2(n_555),
.B1(n_552),
.B2(n_578),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_550),
.B(n_515),
.C(n_525),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_550),
.B(n_532),
.C(n_523),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_572),
.B(n_528),
.C(n_520),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_596),
.C(n_600),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_528),
.C(n_520),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_599),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_573),
.A2(n_558),
.B1(n_517),
.B2(n_553),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_561),
.B(n_557),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_577),
.B(n_531),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_563),
.B(n_514),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_241),
.C(n_321),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_556),
.A2(n_539),
.B1(n_544),
.B2(n_370),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_576),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_553),
.A2(n_346),
.B1(n_345),
.B2(n_326),
.Y(n_604)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_605),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_601),
.Y(n_609)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_610),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_611),
.A2(n_582),
.B1(n_592),
.B2(n_599),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_590),
.B(n_559),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_612),
.B(n_616),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_588),
.A2(n_566),
.B1(n_571),
.B2(n_575),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_613),
.A2(n_617),
.B1(n_589),
.B2(n_600),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_614),
.A2(n_606),
.B1(n_611),
.B2(n_622),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_574),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_SL g617 ( 
.A(n_595),
.B(n_568),
.C(n_570),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_594),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_619),
.B(n_620),
.Y(n_635)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_588),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_580),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_621),
.B(n_626),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_602),
.A2(n_568),
.B1(n_273),
.B2(n_326),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_622),
.A2(n_582),
.B1(n_275),
.B2(n_260),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_623),
.A2(n_251),
.B(n_310),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_593),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_624),
.B(n_284),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_345),
.Y(n_625)
);

NOR2xp67_ASAP7_75t_SL g644 ( 
.A(n_625),
.B(n_277),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_627),
.A2(n_628),
.B1(n_629),
.B2(n_631),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_606),
.A2(n_583),
.B1(n_605),
.B2(n_581),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_624),
.B(n_581),
.C(n_592),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_630),
.B(n_632),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_607),
.B(n_264),
.C(n_277),
.Y(n_632)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_633),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_608),
.A2(n_275),
.B1(n_260),
.B2(n_251),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_637),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_638),
.A2(n_625),
.B(n_626),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_620),
.A2(n_619),
.B1(n_609),
.B2(n_608),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_640),
.B(n_623),
.Y(n_645)
);

FAx1_ASAP7_75t_SL g642 ( 
.A(n_617),
.B(n_310),
.CI(n_284),
.CON(n_642),
.SN(n_642)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_642),
.B(n_644),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_645),
.B(n_646),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_607),
.C(n_615),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_647),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_639),
.B(n_615),
.C(n_618),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_650),
.B(n_657),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_636),
.B(n_618),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_651),
.B(n_653),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_636),
.A2(n_284),
.B(n_264),
.Y(n_652)
);

OA21x2_ASAP7_75t_L g658 ( 
.A1(n_652),
.A2(n_635),
.B(n_641),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_629),
.B(n_308),
.C(n_272),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_633),
.B(n_308),
.C(n_272),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_658),
.A2(n_661),
.B1(n_7),
.B2(n_2),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_SL g660 ( 
.A1(n_648),
.A2(n_641),
.B1(n_631),
.B2(n_643),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_660),
.B(n_662),
.Y(n_667)
);

AOI31xp67_ASAP7_75t_L g661 ( 
.A1(n_646),
.A2(n_635),
.A3(n_642),
.B(n_640),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_654),
.B(n_632),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_649),
.B(n_637),
.C(n_644),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_665),
.B(n_657),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_664),
.B(n_653),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_669),
.Y(n_674)
);

AOI322xp5_ASAP7_75t_L g670 ( 
.A1(n_659),
.A2(n_642),
.A3(n_655),
.B1(n_656),
.B2(n_652),
.C1(n_34),
.C2(n_7),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_670),
.B(n_671),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_658),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_672),
.A2(n_665),
.B1(n_663),
.B2(n_666),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_675),
.B(n_13),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_671),
.B(n_667),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_676),
.A2(n_677),
.B(n_673),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_678),
.B(n_3),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_679),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_SL g681 ( 
.A1(n_680),
.A2(n_4),
.B(n_17),
.C(n_18),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_681),
.A2(n_17),
.B1(n_0),
.B2(n_34),
.Y(n_682)
);


endmodule