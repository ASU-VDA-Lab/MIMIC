module real_aes_15553_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_733;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g863 ( .A(n_0), .B(n_864), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_1), .A2(n_4), .B1(n_261), .B2(n_262), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_2), .A2(n_43), .B1(n_132), .B2(n_161), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_3), .A2(n_24), .B1(n_161), .B2(n_242), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_5), .A2(n_16), .B1(n_522), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_6), .A2(n_119), .B1(n_120), .B2(n_834), .Y(n_118) );
INVx1_ASAP7_75t_L g834 ( .A(n_6), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_7), .A2(n_59), .B1(n_169), .B2(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_8), .A2(n_17), .B1(n_132), .B2(n_134), .Y(n_131) );
INVx1_ASAP7_75t_L g864 ( .A(n_9), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_10), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_11), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_12), .A2(n_18), .B1(n_543), .B2(n_544), .Y(n_542) );
OR2x2_ASAP7_75t_L g108 ( .A(n_13), .B(n_37), .Y(n_108) );
BUFx2_ASAP7_75t_L g869 ( .A(n_13), .Y(n_869) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_14), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_15), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_19), .A2(n_97), .B1(n_262), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_20), .A2(n_38), .B1(n_204), .B2(n_579), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_21), .B(n_203), .Y(n_576) );
OAI21x1_ASAP7_75t_L g144 ( .A1(n_22), .A2(n_57), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_23), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_25), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_26), .B(n_137), .Y(n_217) );
INVx4_ASAP7_75t_R g185 ( .A(n_27), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_28), .A2(n_46), .B1(n_139), .B2(n_259), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_29), .A2(n_53), .B1(n_139), .B2(n_522), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_30), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_31), .B(n_579), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_32), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_33), .B(n_161), .Y(n_224) );
INVx1_ASAP7_75t_L g266 ( .A(n_34), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_SL g239 ( .A1(n_35), .A2(n_132), .B(n_136), .C(n_240), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_36), .A2(n_54), .B1(n_132), .B2(n_139), .Y(n_248) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_37), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_39), .A2(n_84), .B1(n_132), .B2(n_588), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_40), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_41), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_42), .A2(n_45), .B1(n_132), .B2(n_134), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_44), .A2(n_58), .B1(n_522), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g221 ( .A(n_47), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_48), .B(n_132), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_49), .Y(n_159) );
INVx2_ASAP7_75t_L g114 ( .A(n_50), .Y(n_114) );
INVx1_ASAP7_75t_L g106 ( .A(n_51), .Y(n_106) );
BUFx3_ASAP7_75t_L g117 ( .A(n_51), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_52), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_55), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_56), .A2(n_86), .B1(n_132), .B2(n_139), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_60), .A2(n_73), .B1(n_259), .B2(n_524), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_61), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_62), .A2(n_76), .B1(n_132), .B2(n_134), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_63), .A2(n_95), .B1(n_522), .B2(n_544), .Y(n_565) );
INVx1_ASAP7_75t_L g145 ( .A(n_64), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_65), .B(n_148), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_66), .A2(n_510), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_66), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_67), .A2(n_88), .B1(n_139), .B2(n_259), .Y(n_258) );
AO22x1_ASAP7_75t_L g201 ( .A1(n_68), .A2(n_74), .B1(n_202), .B2(n_204), .Y(n_201) );
INVx1_ASAP7_75t_L g148 ( .A(n_69), .Y(n_148) );
AND2x2_ASAP7_75t_L g243 ( .A(n_70), .B(n_155), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_71), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_72), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_75), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g137 ( .A(n_77), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_78), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_79), .B(n_155), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_80), .A2(n_96), .B1(n_139), .B2(n_169), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_81), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_82), .B(n_143), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_83), .Y(n_560) );
INVx1_ASAP7_75t_L g871 ( .A(n_85), .Y(n_871) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_87), .B(n_155), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_89), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_90), .B(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_91), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g509 ( .A(n_91), .Y(n_509) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_92), .B(n_203), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_93), .A2(n_141), .B(n_169), .C(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g189 ( .A(n_94), .B(n_190), .Y(n_189) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_98), .B(n_167), .Y(n_166) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_858), .B(n_870), .Y(n_99) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_110), .Y(n_100) );
INVxp67_ASAP7_75t_L g849 ( .A(n_101), .Y(n_849) );
NOR2xp33_ASAP7_75t_SL g101 ( .A(n_102), .B(n_109), .Y(n_101) );
INVx5_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x6_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
HB1xp67_ASAP7_75t_L g848 ( .A(n_106), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_107), .B(n_116), .Y(n_115) );
AND3x2_ASAP7_75t_L g847 ( .A(n_107), .B(n_833), .C(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_108), .B(n_117), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_118), .B(n_835), .Y(n_110) );
INVx6_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_SL g112 ( .A(n_113), .B(n_115), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx3_ASAP7_75t_L g838 ( .A(n_114), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_114), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22x1_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_506), .B1(n_510), .B2(n_831), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_415), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_331), .C(n_362), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_297), .Y(n_123) );
AOI211x1_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_209), .B(n_252), .C(n_283), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_173), .Y(n_126) );
AND2x2_ASAP7_75t_L g438 ( .A(n_127), .B(n_313), .Y(n_438) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_152), .Y(n_127) );
INVx1_ASAP7_75t_L g323 ( .A(n_128), .Y(n_323) );
OR2x2_ASAP7_75t_L g444 ( .A(n_128), .B(n_295), .Y(n_444) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g280 ( .A(n_129), .B(n_153), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_129), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g312 ( .A(n_129), .Y(n_312) );
OR2x2_ASAP7_75t_L g343 ( .A(n_129), .B(n_174), .Y(n_343) );
AND2x2_ASAP7_75t_L g357 ( .A(n_129), .B(n_174), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_129), .B(n_350), .Y(n_394) );
AO31x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_142), .A3(n_146), .B(n_149), .Y(n_129) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B1(n_138), .B2(n_140), .Y(n_130) );
INVx4_ASAP7_75t_L g134 ( .A(n_132), .Y(n_134) );
INVx1_ASAP7_75t_L g524 ( .A(n_132), .Y(n_524) );
INVx1_ASAP7_75t_L g544 ( .A(n_132), .Y(n_544) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
INVx1_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
INVx1_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_133), .Y(n_205) );
INVx1_ASAP7_75t_L g236 ( .A(n_133), .Y(n_236) );
INVx2_ASAP7_75t_L g242 ( .A(n_133), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_134), .A2(n_159), .B(n_160), .C(n_162), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g574 ( .A1(n_134), .A2(n_136), .B(n_575), .C(n_576), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_135), .A2(n_195), .B1(n_247), .B2(n_248), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_135), .A2(n_140), .B1(n_258), .B2(n_260), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_135), .A2(n_521), .B1(n_523), .B2(n_525), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_135), .A2(n_525), .B1(n_531), .B2(n_532), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_135), .A2(n_542), .B1(n_545), .B2(n_546), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_135), .A2(n_525), .B1(n_557), .B2(n_558), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_135), .A2(n_546), .B1(n_565), .B2(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_135), .A2(n_578), .B(n_580), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_135), .A2(n_140), .B1(n_587), .B2(n_589), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_135), .A2(n_525), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_136), .A2(n_166), .B(n_168), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_136), .B(n_201), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_136), .A2(n_194), .B(n_201), .C(n_207), .Y(n_296) );
BUFx8_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g141 ( .A(n_137), .Y(n_141) );
INVx2_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
INVx1_ASAP7_75t_L g220 ( .A(n_137), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_139), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g261 ( .A(n_139), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_140), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_SL g546 ( .A(n_141), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_142), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_142), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx2_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
OAI21xp33_ASAP7_75t_L g207 ( .A1(n_143), .A2(n_199), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_144), .Y(n_156) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_146), .A2(n_230), .A3(n_541), .B(n_547), .Y(n_540) );
AO31x2_ASAP7_75t_L g555 ( .A1(n_146), .A2(n_249), .A3(n_556), .B(n_559), .Y(n_555) );
AO31x2_ASAP7_75t_L g601 ( .A1(n_146), .A2(n_585), .A3(n_602), .B(n_606), .Y(n_601) );
BUFx10_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx10_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
INVx1_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
INVx1_ASAP7_75t_L g264 ( .A(n_147), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx2_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
BUFx2_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_151), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_151), .B(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g274 ( .A(n_152), .Y(n_274) );
AND2x2_ASAP7_75t_L g325 ( .A(n_152), .B(n_191), .Y(n_325) );
AND2x2_ASAP7_75t_L g468 ( .A(n_152), .B(n_174), .Y(n_468) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g292 ( .A(n_153), .Y(n_292) );
AND2x2_ASAP7_75t_L g311 ( .A(n_153), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g348 ( .A(n_153), .Y(n_348) );
AND2x2_ASAP7_75t_L g372 ( .A(n_153), .B(n_174), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g153 ( .A(n_154), .B(n_157), .Y(n_153) );
NOR2x1_ASAP7_75t_L g170 ( .A(n_155), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g249 ( .A(n_155), .Y(n_249) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g225 ( .A(n_156), .B(n_172), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_156), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_156), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g572 ( .A(n_156), .Y(n_572) );
BUFx3_ASAP7_75t_L g585 ( .A(n_156), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_156), .B(n_607), .Y(n_606) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_165), .B(n_170), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_161), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx3_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g259 ( .A(n_167), .Y(n_259) );
INVx1_ASAP7_75t_L g579 ( .A(n_167), .Y(n_579) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AO31x2_ASAP7_75t_L g245 ( .A1(n_172), .A2(n_246), .A3(n_249), .B(n_250), .Y(n_245) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_173), .Y(n_272) );
AND2x2_ASAP7_75t_L g333 ( .A(n_173), .B(n_322), .Y(n_333) );
INVx2_ASAP7_75t_L g465 ( .A(n_173), .Y(n_465) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_191), .Y(n_173) );
INVx1_ASAP7_75t_L g270 ( .A(n_174), .Y(n_270) );
AND2x4_ASAP7_75t_L g282 ( .A(n_174), .B(n_192), .Y(n_282) );
INVx2_ASAP7_75t_L g350 ( .A(n_174), .Y(n_350) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_189), .Y(n_174) );
AO31x2_ASAP7_75t_L g518 ( .A1(n_175), .A2(n_519), .A3(n_520), .B(n_526), .Y(n_518) );
AO31x2_ASAP7_75t_L g529 ( .A1(n_175), .A2(n_263), .A3(n_530), .B(n_533), .Y(n_529) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g547 ( .A(n_177), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_177), .B(n_591), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_183), .B(n_188), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx2_ASAP7_75t_L g198 ( .A(n_181), .Y(n_198) );
INVx1_ASAP7_75t_L g605 ( .A(n_186), .Y(n_605) );
INVx1_ASAP7_75t_L g519 ( .A(n_188), .Y(n_519) );
AND2x2_ASAP7_75t_L g349 ( .A(n_191), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g356 ( .A(n_191), .Y(n_356) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g434 ( .A(n_192), .B(n_350), .Y(n_434) );
AOI21x1_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_200), .B(n_206), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_199), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_195), .A2(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g525 ( .A(n_196), .Y(n_525) );
INVx1_ASAP7_75t_L g543 ( .A(n_198), .Y(n_543) );
INVxp67_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g522 ( .A(n_203), .Y(n_522) );
OAI21xp33_ASAP7_75t_SL g216 ( .A1(n_204), .A2(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_208), .A2(n_232), .B(n_239), .Y(n_231) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_226), .Y(n_210) );
OR2x2_ASAP7_75t_L g339 ( .A(n_211), .B(n_227), .Y(n_339) );
AND2x2_ASAP7_75t_L g477 ( .A(n_211), .B(n_421), .Y(n_477) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x4_ASAP7_75t_L g254 ( .A(n_212), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g359 ( .A(n_212), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_212), .B(n_301), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_212), .B(n_277), .Y(n_414) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g271 ( .A(n_213), .Y(n_271) );
AND2x2_ASAP7_75t_L g287 ( .A(n_213), .B(n_288), .Y(n_287) );
NAND2x1p5_ASAP7_75t_SL g300 ( .A(n_213), .B(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_213), .B(n_277), .Y(n_379) );
AND2x2_ASAP7_75t_L g427 ( .A(n_213), .B(n_256), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_213), .B(n_255), .Y(n_470) );
BUFx2_ASAP7_75t_L g489 ( .A(n_213), .Y(n_489) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_225), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
BUFx4f_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g273 ( .A(n_227), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g386 ( .A(n_227), .Y(n_386) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_244), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_228), .B(n_256), .Y(n_289) );
INVx2_ASAP7_75t_L g301 ( .A(n_228), .Y(n_301) );
AND2x2_ASAP7_75t_L g337 ( .A(n_228), .B(n_245), .Y(n_337) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g277 ( .A(n_229), .Y(n_277) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_243), .Y(n_229) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_230), .A2(n_257), .A3(n_263), .B(n_265), .Y(n_256) );
AO31x2_ASAP7_75t_L g563 ( .A1(n_230), .A2(n_519), .A3(n_564), .B(n_567), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_235), .B(n_238), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g262 ( .A(n_236), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_SL g588 ( .A(n_242), .Y(n_588) );
INVx1_ASAP7_75t_L g361 ( .A(n_244), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_244), .B(n_256), .Y(n_378) );
INVx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
BUFx2_ASAP7_75t_L g288 ( .A(n_245), .Y(n_288) );
OR2x2_ASAP7_75t_L g320 ( .A(n_245), .B(n_256), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_245), .B(n_256), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_273), .B1(n_275), .B2(n_279), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_267), .B1(n_271), .B2(n_272), .Y(n_253) );
INVx2_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_254), .B(n_337), .Y(n_351) );
AND2x2_ASAP7_75t_L g385 ( .A(n_254), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx1_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_263), .A2(n_585), .A3(n_586), .B(n_590), .Y(n_584) );
INVx2_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_SL g581 ( .A(n_264), .Y(n_581) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g443 ( .A(n_269), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g324 ( .A(n_270), .Y(n_324) );
AND3x1_ASAP7_75t_L g428 ( .A(n_270), .B(n_291), .C(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g384 ( .A(n_271), .Y(n_384) );
AND2x4_ASAP7_75t_L g420 ( .A(n_271), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g458 ( .A(n_274), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_275), .Y(n_462) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
OR2x2_ASAP7_75t_L g435 ( .A(n_276), .B(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_276), .Y(n_483) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g383 ( .A(n_277), .B(n_361), .Y(n_383) );
AND2x2_ASAP7_75t_L g425 ( .A(n_277), .B(n_292), .Y(n_425) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_277), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_280), .B(n_281), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_280), .A2(n_281), .B(n_345), .C(n_351), .Y(n_344) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_280), .B(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_280), .B(n_438), .Y(n_484) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_282), .B(n_311), .Y(n_330) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_285), .B(n_290), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_289), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_290), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g340 ( .A(n_291), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_291), .B(n_357), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_291), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_291), .B(n_349), .Y(n_505) );
INVx3_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx2_ASAP7_75t_L g488 ( .A(n_292), .Y(n_488) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g314 ( .A(n_295), .Y(n_314) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_310), .B(n_315), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_304), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
OAI33xp33_ASAP7_75t_L g364 ( .A1(n_300), .A2(n_305), .A3(n_365), .B1(n_366), .B2(n_368), .B3(n_369), .Y(n_364) );
OR2x2_ASAP7_75t_L g496 ( .A(n_300), .B(n_320), .Y(n_496) );
INVx2_ASAP7_75t_L g498 ( .A(n_300), .Y(n_498) );
INVx1_ASAP7_75t_L g319 ( .A(n_301), .Y(n_319) );
OR2x2_ASAP7_75t_L g360 ( .A(n_301), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g368 ( .A(n_305), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g486 ( .A(n_305), .B(n_487), .C(n_489), .Y(n_486) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_306), .B(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_306), .B(n_470), .Y(n_474) );
AND2x4_ASAP7_75t_L g503 ( .A(n_306), .B(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g329 ( .A(n_308), .Y(n_329) );
OR2x2_ASAP7_75t_L g335 ( .A(n_308), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g448 ( .A(n_308), .B(n_383), .Y(n_448) );
INVx1_ASAP7_75t_L g504 ( .A(n_308), .Y(n_504) );
AND2x4_ASAP7_75t_SL g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g327 ( .A(n_311), .Y(n_327) );
INVx1_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
AND2x2_ASAP7_75t_L g411 ( .A(n_312), .B(n_314), .Y(n_411) );
INVx1_ASAP7_75t_L g451 ( .A(n_313), .Y(n_451) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_321), .B1(n_328), .B2(n_330), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g407 ( .A(n_320), .Y(n_407) );
INVx2_ASAP7_75t_L g421 ( .A(n_320), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_325), .C(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_323), .B(n_348), .Y(n_450) );
OR2x2_ASAP7_75t_L g466 ( .A(n_323), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g479 ( .A(n_323), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_325), .B(n_393), .Y(n_454) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_332), .B(n_352), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B1(n_338), .B2(n_340), .C(n_344), .Y(n_332) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI32xp33_ASAP7_75t_L g501 ( .A1(n_335), .A2(n_432), .A3(n_450), .B1(n_502), .B2(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g471 ( .A(n_337), .Y(n_471) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g352 ( .A1(n_340), .A2(n_353), .B(n_358), .Y(n_352) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_341), .B(n_488), .Y(n_500) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AND2x2_ASAP7_75t_L g494 ( .A(n_347), .B(n_375), .Y(n_494) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
INVx2_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
AND2x2_ASAP7_75t_L g371 ( .A(n_355), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g390 ( .A(n_356), .Y(n_390) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_380), .C(n_391), .D(n_402), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_371), .B1(n_373), .B2(n_376), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_365), .A2(n_493), .B1(n_495), .B2(n_496), .Y(n_492) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g475 ( .A(n_370), .B(n_434), .Y(n_475) );
AND2x2_ASAP7_75t_L g478 ( .A(n_372), .B(n_479), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_392), .B1(n_396), .B2(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
OR2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g397 ( .A(n_379), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_385), .B(n_387), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_381), .A2(n_486), .B(n_490), .C(n_492), .Y(n_485) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g460 ( .A(n_383), .Y(n_460) );
AND2x4_ASAP7_75t_L g453 ( .A(n_386), .B(n_427), .Y(n_453) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g418 ( .A1(n_393), .A2(n_419), .B(n_422), .Y(n_418) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g424 ( .A(n_394), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_394), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g400 ( .A(n_398), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_400), .A2(n_431), .B1(n_435), .B2(n_437), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_409), .B2(n_412), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_407), .Y(n_423) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_480), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_417), .B(n_439), .C(n_455), .D(n_472), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_430), .Y(n_417) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g482 ( .A(n_420), .B(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_426), .B2(n_428), .Y(n_422) );
INVxp67_ASAP7_75t_L g446 ( .A(n_426), .Y(n_446) );
BUFx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g436 ( .A(n_427), .Y(n_436) );
AND2x2_ASAP7_75t_L g459 ( .A(n_427), .B(n_460), .Y(n_459) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_445), .B(n_447), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g464 ( .A(n_442), .B(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g461 ( .A(n_443), .Y(n_461) );
OAI32xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .A3(n_451), .B1(n_452), .B2(n_454), .Y(n_447) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B1(n_461), .B2(n_462), .C(n_463), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B(n_469), .Y(n_463) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g495 ( .A(n_474), .Y(n_495) );
INVx1_ASAP7_75t_L g491 ( .A(n_475), .Y(n_491) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
OAI211xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_484), .B(n_485), .C(n_497), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_501), .Y(n_497) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
BUFx8_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g856 ( .A(n_508), .B(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g833 ( .A(n_509), .Y(n_833) );
INVx2_ASAP7_75t_L g841 ( .A(n_510), .Y(n_841) );
AND3x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_693), .C(n_747), .Y(n_510) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_653), .Y(n_511) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_592), .C(n_635), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_535), .B(n_550), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g685 ( .A(n_516), .B(n_596), .Y(n_685) );
INVx2_ASAP7_75t_L g711 ( .A(n_516), .Y(n_711) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
INVx1_ASAP7_75t_L g610 ( .A(n_517), .Y(n_610) );
INVx2_ASAP7_75t_L g725 ( .A(n_517), .Y(n_725) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g538 ( .A(n_518), .Y(n_538) );
AND2x4_ASAP7_75t_L g668 ( .A(n_518), .B(n_630), .Y(n_668) );
INVx1_ASAP7_75t_L g721 ( .A(n_528), .Y(n_721) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g549 ( .A(n_529), .Y(n_549) );
AND2x4_ASAP7_75t_L g599 ( .A(n_529), .B(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_529), .Y(n_627) );
INVx2_ASAP7_75t_L g630 ( .A(n_529), .Y(n_630) );
OR2x2_ASAP7_75t_L g644 ( .A(n_529), .B(n_601), .Y(n_644) );
AND2x2_ASAP7_75t_L g746 ( .A(n_529), .B(n_540), .Y(n_746) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_536), .B(n_802), .Y(n_801) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
OR2x2_ASAP7_75t_L g628 ( .A(n_537), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_537), .B(n_647), .Y(n_692) );
AND2x2_ASAP7_75t_L g757 ( .A(n_537), .B(n_733), .Y(n_757) );
INVx4_ASAP7_75t_L g791 ( .A(n_537), .Y(n_791) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g626 ( .A(n_538), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_538), .B(n_598), .Y(n_664) );
AND2x2_ASAP7_75t_L g774 ( .A(n_538), .B(n_601), .Y(n_774) );
AND2x2_ASAP7_75t_L g808 ( .A(n_538), .B(n_630), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
INVx4_ASAP7_75t_SL g598 ( .A(n_540), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_540), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g709 ( .A(n_540), .B(n_601), .Y(n_709) );
BUFx2_ASAP7_75t_L g727 ( .A(n_540), .Y(n_727) );
AOI222xp33_ASAP7_75t_L g635 ( .A1(n_549), .A2(n_636), .B1(n_641), .B2(n_642), .C1(n_645), .C2(n_649), .Y(n_635) );
INVx1_ASAP7_75t_L g766 ( .A(n_549), .Y(n_766) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_561), .Y(n_550) );
AND2x2_ASAP7_75t_L g803 ( .A(n_551), .B(n_615), .Y(n_803) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g824 ( .A(n_552), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g633 ( .A(n_553), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_553), .B(n_616), .Y(n_772) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_554), .B(n_620), .Y(n_662) );
AND2x2_ASAP7_75t_L g690 ( .A(n_554), .B(n_570), .Y(n_690) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g619 ( .A(n_555), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g652 ( .A(n_555), .B(n_584), .Y(n_652) );
INVx1_ASAP7_75t_L g680 ( .A(n_555), .Y(n_680) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_555), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_561), .A2(n_678), .B1(n_736), .B2(n_737), .C1(n_739), .C2(n_741), .Y(n_735) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g670 ( .A(n_562), .Y(n_670) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g616 ( .A(n_563), .Y(n_616) );
AND2x2_ASAP7_75t_L g621 ( .A(n_563), .B(n_584), .Y(n_621) );
AND2x2_ASAP7_75t_L g681 ( .A(n_563), .B(n_583), .Y(n_681) );
AND2x2_ASAP7_75t_L g669 ( .A(n_569), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g764 ( .A(n_569), .B(n_680), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_569), .B(n_771), .Y(n_770) );
AND3x1_ASAP7_75t_L g829 ( .A(n_569), .B(n_599), .C(n_830), .Y(n_829) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_583), .Y(n_569) );
AND2x2_ASAP7_75t_L g650 ( .A(n_570), .B(n_616), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_570), .B(n_752), .Y(n_799) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx2_ASAP7_75t_L g613 ( .A(n_571), .Y(n_613) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B(n_582), .Y(n_571) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_572), .A2(n_573), .B(n_582), .Y(n_620) );
OAI21x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .B(n_581), .Y(n_573) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g615 ( .A(n_584), .B(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g648 ( .A(n_584), .B(n_634), .Y(n_648) );
INVx1_ASAP7_75t_L g658 ( .A(n_584), .Y(n_658) );
BUFx2_ASAP7_75t_L g752 ( .A(n_584), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_611), .B(n_617), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2x1_ASAP7_75t_L g594 ( .A(n_595), .B(n_608), .Y(n_594) );
AOI221xp5_ASAP7_75t_SL g675 ( .A1(n_595), .A2(n_676), .B1(n_682), .B2(n_686), .C(n_691), .Y(n_675) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_597), .B(n_610), .Y(n_796) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_598), .B(n_630), .Y(n_629) );
AND2x4_ASAP7_75t_L g638 ( .A(n_598), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g674 ( .A(n_598), .Y(n_674) );
INVx1_ASAP7_75t_L g684 ( .A(n_598), .Y(n_684) );
AND2x2_ASAP7_75t_L g703 ( .A(n_598), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g715 ( .A(n_598), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_598), .B(n_721), .Y(n_828) );
INVx2_ASAP7_75t_L g663 ( .A(n_599), .Y(n_663) );
AND2x2_ASAP7_75t_L g673 ( .A(n_599), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_599), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_599), .B(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g624 ( .A(n_601), .Y(n_624) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_601), .Y(n_667) );
INVx1_ASAP7_75t_L g704 ( .A(n_601), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_601), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g643 ( .A(n_609), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_609), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_610), .Y(n_702) );
NOR2xp33_ASAP7_75t_R g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_613), .B(n_683), .C(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g714 ( .A(n_613), .B(n_621), .Y(n_714) );
AND2x2_ASAP7_75t_L g743 ( .A(n_613), .B(n_713), .Y(n_743) );
OR2x2_ASAP7_75t_L g810 ( .A(n_613), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_L g736 ( .A(n_615), .B(n_619), .Y(n_736) );
INVx2_ASAP7_75t_SL g820 ( .A(n_615), .Y(n_820) );
INVx2_ASAP7_75t_L g647 ( .A(n_616), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_616), .B(n_661), .Y(n_660) );
INVx3_ASAP7_75t_L g689 ( .A(n_616), .Y(n_689) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_616), .Y(n_762) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_622), .A3(n_625), .B1(n_628), .B2(n_631), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g641 ( .A(n_619), .B(n_621), .Y(n_641) );
AND2x2_ASAP7_75t_L g699 ( .A(n_619), .B(n_681), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_619), .B(n_681), .Y(n_707) );
INVx1_ASAP7_75t_L g634 ( .A(n_620), .Y(n_634) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_621), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g776 ( .A(n_621), .Y(n_776) );
INVx2_ASAP7_75t_L g811 ( .A(n_621), .Y(n_811) );
AND2x2_ASAP7_75t_L g823 ( .A(n_621), .B(n_690), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_622), .B(n_744), .C(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g639 ( .A(n_624), .Y(n_639) );
AOI321xp33_ASAP7_75t_L g822 ( .A1(n_625), .A2(n_684), .A3(n_823), .B1(n_824), .B2(n_826), .C(n_829), .Y(n_822) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g640 ( .A(n_627), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_629), .A2(n_648), .B1(n_827), .B2(n_828), .Y(n_826) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g729 ( .A(n_633), .B(n_688), .Y(n_729) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g763 ( .A(n_638), .Y(n_763) );
NAND2x1_ASAP7_75t_L g790 ( .A(n_638), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_638), .B(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g788 ( .A(n_640), .B(n_774), .Y(n_788) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g728 ( .A(n_644), .Y(n_728) );
OR2x2_ASAP7_75t_L g795 ( .A(n_644), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_647), .B(n_648), .Y(n_672) );
NOR2x1p5_ASAP7_75t_L g713 ( .A(n_647), .B(n_652), .Y(n_713) );
INVx1_ASAP7_75t_L g783 ( .A(n_647), .Y(n_783) );
NOR2x1_ASAP7_75t_L g784 ( .A(n_648), .B(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVxp67_ASAP7_75t_SL g827 ( .A(n_650), .Y(n_827) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_665), .C(n_675), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_663), .C(n_664), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g805 ( .A(n_659), .Y(n_805) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g697 ( .A(n_662), .Y(n_697) );
INVx1_ASAP7_75t_L g733 ( .A(n_662), .Y(n_733) );
NAND2xp33_ASAP7_75t_L g737 ( .A(n_663), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g741 ( .A(n_663), .Y(n_741) );
INVx1_ASAP7_75t_L g767 ( .A(n_664), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B(n_671), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx3_ASAP7_75t_L g716 ( .A(n_668), .Y(n_716) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g793 ( .A(n_680), .B(n_783), .Y(n_793) );
AND2x2_ASAP7_75t_L g696 ( .A(n_681), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g761 ( .A(n_681), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
OR2x2_ASAP7_75t_L g719 ( .A(n_684), .B(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g698 ( .A(n_685), .Y(n_698) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g732 ( .A(n_689), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g821 ( .A(n_690), .Y(n_821) );
NOR2xp67_ASAP7_75t_L g693 ( .A(n_694), .B(n_730), .Y(n_693) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_705), .C(n_717), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g738 ( .A(n_703), .Y(n_738) );
AND2x2_ASAP7_75t_L g813 ( .A(n_703), .B(n_724), .Y(n_813) );
INVx1_ASAP7_75t_L g760 ( .A(n_704), .Y(n_760) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI32xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .A3(n_710), .B1(n_712), .B2(n_715), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g740 ( .A(n_709), .Y(n_740) );
NAND2x1_ASAP7_75t_L g778 ( .A(n_709), .B(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g739 ( .A(n_711), .B(n_740), .Y(n_739) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
OAI211xp5_ASAP7_75t_SL g765 ( .A1(n_716), .A2(n_759), .B(n_766), .C(n_767), .Y(n_765) );
INVx2_ASAP7_75t_L g779 ( .A(n_716), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .B(n_729), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_723), .Y(n_734) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx2_ASAP7_75t_L g817 ( .A(n_724), .Y(n_817) );
INVx3_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g825 ( .A(n_725), .B(n_760), .Y(n_825) );
AND2x2_ASAP7_75t_L g830 ( .A(n_725), .B(n_786), .Y(n_830) );
AND2x4_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g755 ( .A(n_728), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_734), .B(n_735), .C(n_742), .Y(n_730) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
NAND2x1p5_ASAP7_75t_L g749 ( .A(n_732), .B(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx2_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_780), .C(n_809), .Y(n_747) );
OAI211xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_753), .B(n_756), .C(n_768), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_754), .A2(n_793), .B1(n_794), .B2(n_797), .Y(n_792) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B1(n_764), .B2(n_765), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_759), .B(n_791), .Y(n_802) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g773 ( .A(n_766), .B(n_774), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_773), .B1(n_775), .B2(n_777), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g798 ( .A(n_772), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI211xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_787), .B(n_792), .C(n_800), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_SL g797 ( .A(n_798), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B1(n_804), .B2(n_806), .Y(n_800) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI211xp5_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_812), .B(n_814), .C(n_822), .Y(n_809) );
INVxp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
INVx4_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_833), .B(n_863), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_839), .B(n_850), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
BUFx8_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
OAI21xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_843), .B(n_849), .Y(n_839) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx4_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NOR2x1p5_ASAP7_75t_L g861 ( .A(n_848), .B(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx10_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx11_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
OR2x6_ASAP7_75t_L g859 ( .A(n_860), .B(n_865), .Y(n_859) );
OR2x6_ASAP7_75t_L g873 ( .A(n_860), .B(n_865), .Y(n_873) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NOR2x1p5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx5_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
endmodule