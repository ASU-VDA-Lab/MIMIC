module fake_jpeg_17873_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_59),
.B1(n_70),
.B2(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

OR2x4_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_36),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_66),
.B(n_21),
.C(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_19),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_24),
.B1(n_28),
.B2(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_60),
.B(n_64),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_33),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_22),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_45),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_24),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_44),
.B(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_35),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_28),
.B1(n_34),
.B2(n_29),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_43),
.B1(n_41),
.B2(n_20),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_34),
.B(n_1),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_75),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_43),
.B1(n_41),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_81),
.B1(n_88),
.B2(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_74),
.A2(n_86),
.B1(n_23),
.B2(n_26),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_43),
.B1(n_41),
.B2(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_104),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_0),
.B1(n_69),
.B2(n_48),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_44),
.B1(n_20),
.B2(n_32),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_97),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_44),
.B1(n_21),
.B2(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_31),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_63),
.A3(n_49),
.B1(n_59),
.B2(n_51),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_78),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_63),
.C(n_53),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_113),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_52),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_91),
.B1(n_88),
.B2(n_74),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_70),
.A3(n_65),
.B1(n_31),
.B2(n_30),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_129),
.B1(n_72),
.B2(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_80),
.B(n_30),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_0),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_130),
.B(n_96),
.Y(n_134)
);

OA22x2_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_68),
.B1(n_50),
.B2(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_1),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_18),
.C(n_50),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_87),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_26),
.C(n_18),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_18),
.C(n_2),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_134),
.B(n_137),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_135),
.A2(n_144),
.B(n_148),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_96),
.B(n_79),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_123),
.B(n_130),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_102),
.B1(n_77),
.B2(n_69),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_95),
.B1(n_90),
.B2(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_151),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_48),
.B1(n_68),
.B2(n_67),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_97),
.B(n_76),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_5),
.C(n_6),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_89),
.B1(n_78),
.B2(n_105),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_93),
.B(n_2),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_153),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_93),
.B(n_92),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_150),
.A2(n_157),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_1),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_93),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_3),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_4),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_106),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_154),
.Y(n_199)
);

AOI221xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_175),
.B1(n_183),
.B2(n_145),
.C(n_161),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_113),
.C(n_123),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_189),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_132),
.C(n_110),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_179),
.C(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_130),
.B(n_117),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_110),
.C(n_124),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_124),
.C(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_136),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_142),
.C(n_134),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_159),
.C(n_146),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_138),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_121),
.Y(n_189)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_199),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_197),
.A2(n_191),
.B(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_169),
.B(n_145),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_209),
.Y(n_227)
);

OA21x2_ASAP7_75t_SL g223 ( 
.A1(n_202),
.A2(n_185),
.B(n_168),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_137),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_210),
.C(n_5),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_152),
.C(n_153),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_152),
.B1(n_150),
.B2(n_139),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_214),
.B1(n_187),
.B2(n_191),
.Y(n_217)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_150),
.B1(n_155),
.B2(n_148),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_203),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_230),
.B1(n_204),
.B2(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_164),
.B1(n_179),
.B2(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_223),
.B1(n_225),
.B2(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_229),
.C(n_233),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_194),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_164),
.B1(n_178),
.B2(n_190),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_180),
.B(n_178),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_231),
.B(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_173),
.B1(n_163),
.B2(n_192),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_167),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_192),
.B1(n_162),
.B2(n_116),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_116),
.B(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_6),
.C(n_7),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_208),
.C(n_233),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

INVx11_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_231),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_207),
.C(n_210),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_243),
.C(n_226),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_242),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_198),
.C(n_212),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_7),
.Y(n_246)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_230),
.Y(n_247)
);

NAND4xp25_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_249),
.C(n_9),
.D(n_10),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_8),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_252),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_222),
.B(n_225),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_253),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_228),
.CI(n_219),
.CON(n_255),
.SN(n_255)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_232),
.B1(n_224),
.B2(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_261),
.B1(n_12),
.B2(n_15),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_260),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_270),
.B1(n_271),
.B2(n_250),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_237),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_265),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_241),
.B1(n_235),
.B2(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_256),
.B(n_252),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_10),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_16),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_254),
.B(n_259),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_250),
.B(n_255),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_255),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_278),
.B(n_271),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_280),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_275),
.A2(n_267),
.B(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

AO22x1_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_268),
.B1(n_251),
.B2(n_256),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_286),
.B(n_283),
.CI(n_16),
.CON(n_288),
.SN(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_284),
.C(n_287),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_288),
.Y(n_290)
);


endmodule