module fake_jpeg_2268_n_528 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_528);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_7),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_26),
.A2(n_7),
.B1(n_1),
.B2(n_2),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_17),
.B1(n_52),
.B2(n_46),
.Y(n_126)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_72),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_28),
.B(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_8),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_50),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_93),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_28),
.B(n_11),
.C(n_4),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_17),
.C(n_52),
.Y(n_166)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_11),
.Y(n_93)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_99),
.Y(n_155)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_44),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_37),
.C(n_41),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_123),
.C(n_19),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_130),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_45),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_73),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_124),
.B(n_139),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_166),
.Y(n_221)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_67),
.B(n_35),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_65),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_92),
.B1(n_75),
.B2(n_83),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_143),
.A2(n_172),
.B1(n_159),
.B2(n_167),
.Y(n_224)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_160),
.Y(n_214)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_54),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_101),
.Y(n_181)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_59),
.Y(n_170)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_98),
.A2(n_52),
.B1(n_53),
.B2(n_47),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_178),
.Y(n_235)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_60),
.B1(n_99),
.B2(n_66),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_115),
.B(n_108),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_179),
.B(n_184),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_180),
.A2(n_222),
.B1(n_160),
.B2(n_164),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_181),
.B(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_108),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_84),
.C(n_97),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_131),
.B(n_37),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_187),
.B(n_193),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_189),
.Y(n_228)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_118),
.B(n_64),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_114),
.A2(n_61),
.B1(n_36),
.B2(n_53),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_203),
.B1(n_212),
.B2(n_42),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_94),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_202),
.B(n_204),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_114),
.A2(n_34),
.B1(n_53),
.B2(n_36),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_120),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_207),
.B(n_223),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_91),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_136),
.Y(n_245)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_119),
.A2(n_38),
.B1(n_34),
.B2(n_47),
.Y(n_212)
);

BUFx4f_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_148),
.Y(n_219)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_134),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_123),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_145),
.B1(n_154),
.B2(n_159),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_131),
.B(n_48),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_226),
.B(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_130),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_250),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_143),
.B1(n_147),
.B2(n_133),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_241),
.A2(n_249),
.B1(n_257),
.B2(n_263),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_224),
.B1(n_195),
.B2(n_183),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_245),
.B(n_200),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_144),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_214),
.B1(n_112),
.B2(n_220),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_177),
.B(n_157),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_171),
.B1(n_149),
.B2(n_167),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_226),
.A2(n_140),
.B1(n_122),
.B2(n_145),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_SL g264 ( 
.A(n_189),
.B(n_95),
.C(n_150),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_218),
.Y(n_291)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_224),
.B1(n_186),
.B2(n_154),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_272),
.A2(n_284),
.B1(n_287),
.B2(n_290),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_191),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_275),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_274),
.A2(n_286),
.B1(n_288),
.B2(n_238),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_227),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_214),
.B1(n_190),
.B2(n_215),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_277),
.A2(n_291),
.B(n_233),
.Y(n_325)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_202),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_279),
.B(n_281),
.Y(n_322)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_178),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_282),
.Y(n_308)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_185),
.B1(n_122),
.B2(n_140),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_294),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_185),
.B1(n_217),
.B2(n_208),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_128),
.B1(n_132),
.B2(n_217),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_242),
.A2(n_208),
.B1(n_205),
.B2(n_213),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_241),
.A2(n_128),
.B1(n_132),
.B2(n_205),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_240),
.B1(n_235),
.B2(n_262),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_281),
.B1(n_269),
.B2(n_279),
.Y(n_307)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_231),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_298),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_255),
.B(n_236),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_192),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_211),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_235),
.B(n_215),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_300),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_235),
.B(n_206),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_264),
.C(n_266),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_310),
.C(n_317),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_330),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_288),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_266),
.C(n_259),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_234),
.B1(n_213),
.B2(n_238),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_316),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_292),
.A2(n_229),
.B1(n_237),
.B2(n_210),
.Y(n_312)
);

HAxp5_ASAP7_75t_SL g313 ( 
.A(n_273),
.B(n_251),
.CON(n_313),
.SN(n_313)
);

INVx2_ASAP7_75t_R g332 ( 
.A(n_313),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_229),
.B1(n_237),
.B2(n_261),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_272),
.A2(n_253),
.B1(n_259),
.B2(n_260),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_248),
.C(n_261),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_284),
.A2(n_260),
.B1(n_246),
.B2(n_243),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_327),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_325),
.A2(n_291),
.B(n_277),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_246),
.B1(n_243),
.B2(n_247),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_247),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_254),
.C(n_290),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_298),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_325),
.A2(n_291),
.B(n_289),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_334),
.A2(n_345),
.B(n_347),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_300),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_310),
.C(n_317),
.Y(n_364)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

INVx13_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_352),
.B1(n_222),
.B2(n_188),
.Y(n_377)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_322),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_343),
.A2(n_357),
.B(n_287),
.Y(n_387)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_344),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_350),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_285),
.B(n_299),
.Y(n_347)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_270),
.A3(n_276),
.B1(n_294),
.B2(n_280),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_316),
.B(n_286),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_321),
.Y(n_351)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_351),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_326),
.A2(n_283),
.B1(n_278),
.B2(n_268),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_354),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_296),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_302),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_329),
.C(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_295),
.B(n_282),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_359),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_282),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_306),
.B1(n_320),
.B2(n_311),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_377),
.B1(n_333),
.B2(n_353),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_303),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_363),
.B(n_371),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_343),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_328),
.C(n_308),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_375),
.C(n_379),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_312),
.B(n_318),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_370),
.B(n_378),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_233),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_373),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_254),
.C(n_196),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_216),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_135),
.C(n_197),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_346),
.A2(n_309),
.B1(n_314),
.B2(n_306),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_381),
.A2(n_384),
.B1(n_350),
.B2(n_333),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_346),
.A2(n_323),
.B1(n_327),
.B2(n_290),
.Y(n_384)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_350),
.Y(n_400)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_334),
.C(n_359),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_342),
.C(n_341),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_390),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_390),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_392),
.B(n_404),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_393),
.A2(n_409),
.B1(n_381),
.B2(n_380),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_405),
.Y(n_438)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_376),
.Y(n_395)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_382),
.B1(n_367),
.B2(n_385),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_400),
.B(n_387),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_386),
.A2(n_332),
.B(n_336),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_402),
.A2(n_412),
.B(n_417),
.Y(n_428)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_383),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_332),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_408),
.B(n_379),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_336),
.B1(n_344),
.B2(n_331),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_413),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_360),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_374),
.A2(n_339),
.B(n_174),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_415),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_268),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_416),
.B(n_38),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_168),
.B(n_225),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_365),
.A2(n_112),
.B(n_155),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_419),
.A2(n_201),
.B(n_96),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_409),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_407),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_426),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_423),
.A2(n_431),
.B1(n_433),
.B2(n_435),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_389),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_429),
.C(n_436),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_375),
.C(n_366),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_393),
.A2(n_380),
.B1(n_384),
.B2(n_364),
.Y(n_431)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_432),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_406),
.A2(n_369),
.B1(n_382),
.B2(n_367),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_155),
.C(n_201),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_419),
.B(n_403),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_400),
.C(n_414),
.Y(n_459)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_418),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_442),
.B(n_396),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_421),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_445),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_425),
.A2(n_406),
.B1(n_412),
.B2(n_416),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_451),
.B1(n_455),
.B2(n_461),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_421),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_410),
.Y(n_446)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_434),
.A2(n_397),
.B1(n_407),
.B2(n_411),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_454),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_423),
.A2(n_413),
.B1(n_417),
.B2(n_395),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_458),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_453),
.Y(n_471)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_14),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_431),
.A2(n_42),
.B1(n_38),
.B2(n_36),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_457),
.A2(n_434),
.B1(n_428),
.B2(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_462),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_429),
.C(n_422),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_463),
.B(n_468),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_457),
.A2(n_428),
.B1(n_441),
.B2(n_439),
.Y(n_465)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_438),
.C(n_427),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_L g470 ( 
.A1(n_459),
.A2(n_426),
.B(n_437),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_470),
.A2(n_152),
.B(n_95),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_468),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_454),
.A2(n_438),
.B1(n_436),
.B2(n_42),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_475),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_449),
.B(n_22),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_476),
.B(n_477),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_446),
.B(n_451),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_456),
.B(n_22),
.Y(n_478)
);

NAND3xp33_ASAP7_75t_SL g489 ( 
.A(n_478),
.B(n_21),
.C(n_29),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_444),
.B(n_455),
.Y(n_480)
);

AOI21xp33_ASAP7_75t_L g502 ( 
.A1(n_480),
.A2(n_492),
.B(n_470),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_493),
.Y(n_496)
);

MAJx2_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_453),
.C(n_458),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_491),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_461),
.C(n_448),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_488),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_448),
.C(n_460),
.Y(n_488)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_489),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_462),
.A2(n_19),
.B(n_46),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_48),
.C(n_71),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_485),
.B(n_472),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_494),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_473),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_501),
.Y(n_513)
);

OAI211xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_467),
.B(n_466),
.C(n_474),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_497),
.A2(n_502),
.B(n_503),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_490),
.B(n_486),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_481),
.B(n_41),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_505),
.Y(n_514)
);

INVx6_ASAP7_75t_L g505 ( 
.A(n_488),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_484),
.A2(n_29),
.B1(n_48),
.B2(n_71),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_5),
.C(n_6),
.Y(n_512)
);

AOI322xp5_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_487),
.A3(n_483),
.B1(n_493),
.B2(n_492),
.C1(n_491),
.C2(n_96),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_510),
.Y(n_515)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_90),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_12),
.Y(n_510)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_90),
.C(n_4),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_7),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_512),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_516),
.B(n_518),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_498),
.B(n_496),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_498),
.C(n_499),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_514),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_515),
.B(n_509),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_522),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_514),
.C(n_517),
.Y(n_523)
);

NOR3xp33_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_13),
.C(n_15),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_524),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_0),
.B1(n_13),
.B2(n_524),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_13),
.B(n_0),
.Y(n_528)
);


endmodule