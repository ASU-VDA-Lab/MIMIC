module fake_netlist_6_1759_n_1073 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1073);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1073;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_955;
wire n_284;
wire n_400;
wire n_337;
wire n_739;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_989;
wire n_843;
wire n_772;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_982;
wire n_831;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_993;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_33),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_76),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_103),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_153),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_51),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_140),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_105),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_156),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_116),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_102),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_119),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_68),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_64),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_31),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_182),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_145),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_190),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_131),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_50),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_41),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_75),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_13),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_57),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_86),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_73),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_146),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_25),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_60),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_78),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_117),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_59),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_11),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_82),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_84),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_122),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_101),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_109),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_98),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_237),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_263),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_258),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_231),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_263),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_205),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_206),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_208),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_214),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_204),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_222),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_272),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_225),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_225),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_230),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_210),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_230),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_296),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_207),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_283),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_209),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_273),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_320),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_316),
.B(n_314),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_213),
.B1(n_268),
.B2(n_267),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_212),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_320),
.B(n_288),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

BUFx8_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_309),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_283),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_226),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_309),
.Y(n_352)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_226),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_269),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_215),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_218),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_219),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_291),
.A2(n_241),
.B1(n_261),
.B2(n_257),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_293),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_236),
.B1(n_256),
.B2(n_223),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_318),
.A2(n_239),
.B1(n_224),
.B2(n_252),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_220),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_300),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_277),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_280),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_228),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_318),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_287),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_324),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_345),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_324),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_359),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_352),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_338),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_338),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_376),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_376),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_299),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_375),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_299),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_375),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_364),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_R g396 ( 
.A(n_371),
.B(n_279),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_364),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_344),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_344),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_366),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_340),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_336),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_333),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_333),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_369),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_373),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_368),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_373),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_357),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_341),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_341),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_331),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_328),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_337),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_342),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_337),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_356),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_370),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_329),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_354),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_325),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_325),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_361),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_355),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_362),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_355),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_R g442 ( 
.A(n_339),
.B(n_298),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_374),
.B(n_306),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_327),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_327),
.Y(n_448)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_386),
.B(n_377),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_416),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_395),
.B1(n_397),
.B2(n_403),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_435),
.B(n_312),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_440),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_441),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_418),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_404),
.B(n_315),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_438),
.B(n_377),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_405),
.B(n_391),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_414),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_382),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_420),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_449),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_310),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_382),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_339),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_439),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_392),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_279),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_437),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_428),
.B(n_363),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_388),
.B(n_363),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_412),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_429),
.B(n_339),
.Y(n_489)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_422),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_229),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_407),
.B(n_232),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_417),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_393),
.B(n_444),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_425),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_444),
.B(n_367),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx8_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_367),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_372),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_389),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_447),
.B(n_353),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_430),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_448),
.B(n_289),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_421),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_353),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_409),
.B(n_234),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_396),
.B(n_372),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_384),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_385),
.B(n_235),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_390),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_442),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_387),
.B(n_326),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_378),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_380),
.Y(n_527)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_398),
.B(n_290),
.C(n_335),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_381),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_414),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_458),
.B(n_343),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_460),
.B(n_242),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_452),
.B(n_244),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_519),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_465),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_458),
.B(n_343),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_476),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_456),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_474),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_462),
.Y(n_543)
);

AOI211xp5_ASAP7_75t_L g544 ( 
.A1(n_491),
.A2(n_245),
.B(n_334),
.C(n_346),
.Y(n_544)
);

OAI221xp5_ASAP7_75t_L g545 ( 
.A1(n_523),
.A2(n_334),
.B1(n_346),
.B2(n_2),
.C(n_3),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_455),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_462),
.B(n_334),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_523),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_483),
.B(n_334),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_524),
.B(n_353),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_450),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_459),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_524),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_480),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_482),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_467),
.Y(n_561)
);

OR2x2_ASAP7_75t_SL g562 ( 
.A(n_517),
.B(n_518),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_471),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_477),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_502),
.B(n_346),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_503),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_530),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_494),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_516),
.A2(n_489),
.B1(n_509),
.B2(n_501),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_468),
.B(n_346),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_484),
.B(n_28),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_486),
.B(n_4),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_499),
.B(n_353),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_483),
.B(n_29),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_454),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_478),
.B(n_4),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_473),
.A2(n_499),
.B1(n_514),
.B2(n_510),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_453),
.B(n_5),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_486),
.B(n_5),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_495),
.B(n_349),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_506),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_503),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_483),
.B(n_504),
.Y(n_590)
);

BUFx6f_ASAP7_75t_SL g591 ( 
.A(n_520),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_567),
.B(n_493),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_582),
.A2(n_481),
.B(n_515),
.C(n_464),
.Y(n_593)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_536),
.A2(n_521),
.B(n_513),
.C(n_504),
.Y(n_594)
);

AO21x2_ASAP7_75t_L g595 ( 
.A1(n_587),
.A2(n_507),
.B(n_525),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_536),
.A2(n_505),
.B(n_531),
.C(n_466),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_534),
.B(n_479),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_591),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_534),
.B(n_510),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_577),
.A2(n_492),
.B(n_461),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_541),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_579),
.B(n_512),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_582),
.A2(n_522),
.B(n_528),
.C(n_457),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_550),
.A2(n_470),
.B(n_349),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_557),
.B(n_470),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_533),
.B(n_512),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_550),
.A2(n_508),
.B(n_470),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_558),
.B(n_470),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_537),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_512),
.C(n_520),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_533),
.B(n_511),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_580),
.A2(n_498),
.B(n_8),
.C(n_9),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_581),
.A2(n_349),
.B(n_527),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_566),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_559),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_574),
.B(n_490),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_570),
.B(n_543),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_573),
.B(n_520),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_545),
.A2(n_527),
.B1(n_526),
.B2(n_529),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_538),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_546),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_L g623 ( 
.A(n_535),
.B(n_502),
.C(n_526),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_547),
.B(n_526),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_541),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_553),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_573),
.A2(n_32),
.B(n_30),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_572),
.B(n_349),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_545),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_541),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_554),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

NOR2x1_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_529),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_561),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_563),
.Y(n_635)
);

OR2x2_ASAP7_75t_SL g636 ( 
.A(n_589),
.B(n_529),
.Y(n_636)
);

NAND2x1p5_ASAP7_75t_L g637 ( 
.A(n_560),
.B(n_35),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_552),
.A2(n_38),
.B(n_37),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_572),
.B(n_250),
.Y(n_639)
);

BUFx4f_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_549),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_40),
.B(n_39),
.Y(n_642)
);

OAI321xp33_ASAP7_75t_L g643 ( 
.A1(n_576),
.A2(n_7),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_643)
);

AND2x4_ASAP7_75t_SL g644 ( 
.A(n_565),
.B(n_42),
.Y(n_644)
);

AOI21x1_ASAP7_75t_L g645 ( 
.A1(n_588),
.A2(n_253),
.B(n_250),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_572),
.B(n_571),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_592),
.B(n_586),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_597),
.B(n_590),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_625),
.Y(n_649)
);

O2A1O1Ixp33_ASAP7_75t_L g650 ( 
.A1(n_593),
.A2(n_583),
.B(n_584),
.C(n_585),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_612),
.B(n_562),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_SL g652 ( 
.A1(n_599),
.A2(n_544),
.B(n_540),
.C(n_564),
.Y(n_652)
);

OAI22x1_ASAP7_75t_L g653 ( 
.A1(n_611),
.A2(n_578),
.B1(n_575),
.B2(n_556),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_598),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_640),
.B(n_578),
.Y(n_656)
);

CKINVDCx14_ASAP7_75t_R g657 ( 
.A(n_607),
.Y(n_657)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_628),
.A2(n_568),
.B(n_542),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_532),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_625),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_605),
.A2(n_539),
.B(n_569),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_640),
.A2(n_591),
.B1(n_556),
.B2(n_548),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_641),
.B(n_548),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_645),
.A2(n_556),
.B(n_548),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_605),
.A2(n_45),
.B(n_43),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_616),
.B(n_250),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_619),
.A2(n_118),
.B(n_203),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_618),
.B(n_265),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_613),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_669)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_633),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_15),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_594),
.A2(n_265),
.B(n_253),
.C(n_250),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_615),
.B(n_250),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_621),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_626),
.Y(n_675)
);

NOR3xp33_ASAP7_75t_SL g676 ( 
.A(n_620),
.B(n_16),
.C(n_17),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_641),
.B(n_253),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_620),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_603),
.A2(n_629),
.B(n_602),
.C(n_596),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_617),
.B(n_265),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

OAI22x1_ASAP7_75t_L g682 ( 
.A1(n_646),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_600),
.A2(n_123),
.B(n_202),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_614),
.A2(n_121),
.B(n_200),
.Y(n_684)
);

O2A1O1Ixp5_ASAP7_75t_L g685 ( 
.A1(n_639),
.A2(n_265),
.B(n_253),
.C(n_21),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_634),
.B(n_19),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_635),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_614),
.A2(n_120),
.B(n_198),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_610),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_622),
.B(n_20),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_644),
.B(n_24),
.Y(n_691)
);

AND2x2_ASAP7_75t_SL g692 ( 
.A(n_623),
.B(n_26),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_606),
.A2(n_26),
.B(n_27),
.C(n_46),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_625),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_595),
.B(n_27),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_636),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_609),
.A2(n_49),
.B(n_52),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_637),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_630),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_660),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_658),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_649),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_654),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_700),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_695),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_660),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_655),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_671),
.A2(n_637),
.B1(n_642),
.B2(n_638),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

INVx6_ASAP7_75t_SL g711 ( 
.A(n_657),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_649),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_647),
.B(n_632),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_697),
.Y(n_714)
);

CKINVDCx16_ASAP7_75t_R g715 ( 
.A(n_670),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_651),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_648),
.B(n_601),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_659),
.B(n_630),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_656),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_692),
.A2(n_627),
.B1(n_630),
.B2(n_608),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_700),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_691),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_674),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_696),
.Y(n_725)
);

AO21x1_ASAP7_75t_L g726 ( 
.A1(n_678),
.A2(n_643),
.B(n_58),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_663),
.Y(n_727)
);

INVx6_ASAP7_75t_L g728 ( 
.A(n_673),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_689),
.Y(n_729)
);

AND2x6_ASAP7_75t_L g730 ( 
.A(n_694),
.B(n_643),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_663),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_675),
.B(n_56),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_681),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_687),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_676),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_677),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_686),
.Y(n_738)
);

BUFx12f_ASAP7_75t_L g739 ( 
.A(n_668),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_664),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_690),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_666),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_679),
.B(n_199),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_685),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_650),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_680),
.B(n_61),
.Y(n_746)
);

INVx5_ASAP7_75t_SL g747 ( 
.A(n_699),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_197),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_653),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_652),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_662),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_62),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_699),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_661),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_693),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_667),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_698),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_683),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_684),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_688),
.Y(n_760)
);

AO21x2_ASAP7_75t_L g761 ( 
.A1(n_702),
.A2(n_665),
.B(n_65),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_702),
.A2(n_63),
.B(n_66),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_722),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_758),
.A2(n_67),
.B(n_69),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_721),
.B(n_70),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_753),
.A2(n_71),
.B(n_72),
.C(n_74),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_713),
.B(n_77),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_754),
.A2(n_79),
.B(n_80),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_760),
.A2(n_81),
.B(n_83),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_747),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_736),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_758),
.A2(n_92),
.B(n_93),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_725),
.B(n_94),
.Y(n_773)
);

BUFx4f_ASAP7_75t_L g774 ( 
.A(n_719),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_756),
.A2(n_95),
.B(n_96),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_719),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_725),
.B(n_97),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_753),
.B(n_99),
.Y(n_778)
);

OAI21x1_ASAP7_75t_L g779 ( 
.A1(n_756),
.A2(n_100),
.B(n_104),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_750),
.A2(n_108),
.B(n_110),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_708),
.B(n_111),
.Y(n_781)
);

OAI21x1_ASAP7_75t_L g782 ( 
.A1(n_750),
.A2(n_112),
.B(n_113),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_708),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_740),
.A2(n_114),
.B(n_115),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_740),
.A2(n_124),
.B(n_125),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_757),
.A2(n_126),
.B(n_127),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_735),
.B(n_128),
.C(n_130),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_716),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_788)
);

AO21x2_ASAP7_75t_L g789 ( 
.A1(n_744),
.A2(n_137),
.B(n_142),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_753),
.B(n_144),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_709),
.A2(n_147),
.B(n_148),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_720),
.A2(n_150),
.B(n_151),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_743),
.A2(n_152),
.B(n_154),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_727),
.A2(n_155),
.B(n_157),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_719),
.Y(n_795)
);

CKINVDCx6p67_ASAP7_75t_R g796 ( 
.A(n_715),
.Y(n_796)
);

AND2x4_ASAP7_75t_SL g797 ( 
.A(n_721),
.B(n_741),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_SL g798 ( 
.A1(n_736),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_723),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_733),
.Y(n_800)
);

AO21x2_ASAP7_75t_L g801 ( 
.A1(n_726),
.A2(n_165),
.B(n_166),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_738),
.B(n_167),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_735),
.A2(n_196),
.B1(n_170),
.B2(n_171),
.Y(n_803)
);

OAI21x1_ASAP7_75t_L g804 ( 
.A1(n_752),
.A2(n_737),
.B(n_724),
.Y(n_804)
);

OA21x2_ASAP7_75t_L g805 ( 
.A1(n_727),
.A2(n_168),
.B(n_173),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_747),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_724),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_704),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_745),
.B(n_178),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_701),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_731),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_807),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_800),
.B(n_741),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_778),
.A2(n_755),
.B1(n_748),
.B2(n_751),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_807),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_763),
.Y(n_816)
);

AOI21x1_ASAP7_75t_L g817 ( 
.A1(n_809),
.A2(n_742),
.B(n_717),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_783),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_811),
.Y(n_819)
);

BUFx4f_ASAP7_75t_SL g820 ( 
.A(n_808),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_804),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_799),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_794),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_762),
.Y(n_824)
);

AO21x2_ASAP7_75t_L g825 ( 
.A1(n_791),
.A2(n_731),
.B(n_746),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_809),
.A2(n_745),
.B(n_718),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_749),
.Y(n_827)
);

INVxp33_ASAP7_75t_L g828 ( 
.A(n_763),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_762),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_794),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_794),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_771),
.A2(n_759),
.B1(n_749),
.B2(n_728),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_773),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_797),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_805),
.B(n_749),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_805),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_805),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_781),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_789),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_797),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_767),
.B(n_741),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_789),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_781),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_808),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_776),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_773),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_777),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_776),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_777),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_761),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_761),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_801),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_801),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_833),
.B(n_734),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_846),
.B(n_796),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_812),
.B(n_795),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_844),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_822),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_812),
.Y(n_859)
);

AND2x2_ASAP7_75t_SL g860 ( 
.A(n_835),
.B(n_771),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_822),
.B(n_795),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_812),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_848),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_848),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_820),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_841),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_815),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_817),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_SL g870 ( 
.A(n_832),
.B(n_798),
.C(n_769),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_846),
.B(n_802),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_815),
.B(n_792),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_818),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_847),
.B(n_723),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_R g875 ( 
.A(n_835),
.B(n_827),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_818),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_818),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_825),
.A2(n_798),
.B1(n_778),
.B2(n_790),
.Y(n_878)
);

CKINVDCx16_ASAP7_75t_R g879 ( 
.A(n_841),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_828),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_R g881 ( 
.A(n_817),
.B(n_715),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_814),
.A2(n_803),
.B1(n_778),
.B2(n_790),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_857),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_873),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_876),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_854),
.B(n_847),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_859),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_876),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_867),
.B(n_819),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_819),
.Y(n_890)
);

OR2x2_ASAP7_75t_L g891 ( 
.A(n_864),
.B(n_837),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_859),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_869),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_870),
.A2(n_825),
.B1(n_803),
.B2(n_770),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_877),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_874),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_877),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_863),
.B(n_819),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_862),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_862),
.B(n_837),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_868),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_858),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_868),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_871),
.B(n_849),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_865),
.B(n_821),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_902),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_904),
.B(n_849),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_884),
.Y(n_908)
);

AO31x2_ASAP7_75t_L g909 ( 
.A1(n_902),
.A2(n_826),
.A3(n_850),
.B(n_824),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_905),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_894),
.A2(n_860),
.B(n_882),
.Y(n_911)
);

AOI211xp5_ASAP7_75t_L g912 ( 
.A1(n_896),
.A2(n_826),
.B(n_806),
.C(n_881),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_905),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_886),
.A2(n_878),
.B1(n_881),
.B2(n_769),
.C(n_869),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_889),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_883),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_893),
.A2(n_860),
.B1(n_825),
.B2(n_790),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_885),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_889),
.B(n_861),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_891),
.B(n_856),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_906),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_908),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_916),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_915),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_920),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_919),
.B(n_890),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_919),
.B(n_890),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_911),
.A2(n_827),
.B1(n_869),
.B2(n_855),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_911),
.B(n_880),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_910),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_913),
.B(n_898),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_921),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_921),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_922),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_924),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_930),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_931),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_926),
.B(n_898),
.Y(n_939)
);

INVxp33_ASAP7_75t_L g940 ( 
.A(n_932),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_932),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_933),
.B(n_929),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_933),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_935),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_934),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_937),
.B(n_923),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_941),
.Y(n_947)
);

INVxp67_ASAP7_75t_SL g948 ( 
.A(n_940),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_941),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_942),
.B(n_938),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_SL g951 ( 
.A(n_943),
.B(n_857),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_946),
.B(n_923),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_944),
.B(n_927),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_945),
.B(n_928),
.Y(n_954)
);

AOI222xp33_ASAP7_75t_SL g955 ( 
.A1(n_941),
.A2(n_928),
.B1(n_936),
.B2(n_816),
.C1(n_912),
.C2(n_914),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_941),
.B(n_939),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_941),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_SL g958 ( 
.A(n_947),
.B(n_866),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_948),
.B(n_918),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_957),
.B(n_907),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_949),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_956),
.B(n_866),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_956),
.B(n_907),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_950),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_953),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_952),
.B(n_866),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_965),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_961),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_966),
.B(n_951),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_962),
.A2(n_954),
.B(n_964),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_959),
.A2(n_914),
.B(n_955),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_958),
.B(n_955),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_960),
.Y(n_974)
);

OAI33xp33_ASAP7_75t_L g975 ( 
.A1(n_963),
.A2(n_891),
.A3(n_850),
.B1(n_852),
.B2(n_853),
.B3(n_900),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_967),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_970),
.B(n_714),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_968),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_969),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_974),
.B(n_917),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_972),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_973),
.B(n_711),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_971),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_975),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_977),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_976),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_978),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_981),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_979),
.B(n_711),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_980),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_983),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_984),
.B(n_909),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_L g994 ( 
.A(n_981),
.B(n_723),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_L g995 ( 
.A(n_990),
.B(n_787),
.C(n_766),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_989),
.B(n_917),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_986),
.B(n_768),
.C(n_786),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_991),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_993),
.B(n_869),
.Y(n_999)
);

NAND4xp25_ASAP7_75t_SL g1000 ( 
.A(n_987),
.B(n_788),
.C(n_768),
.D(n_705),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_985),
.B(n_992),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_988),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_909),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_998),
.A2(n_786),
.B1(n_706),
.B2(n_852),
.C(n_853),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_858),
.B1(n_765),
.B2(n_732),
.C(n_710),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_999),
.A2(n_996),
.B(n_1003),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1002),
.B(n_909),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_997),
.A2(n_765),
.B(n_732),
.C(n_703),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_995),
.Y(n_1009)
);

AOI211xp5_ASAP7_75t_L g1010 ( 
.A1(n_1006),
.A2(n_1000),
.B(n_793),
.C(n_780),
.Y(n_1010)
);

AOI21xp33_ASAP7_75t_SL g1011 ( 
.A1(n_1007),
.A2(n_1008),
.B(n_1009),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_1005),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_1004),
.A2(n_785),
.B(n_784),
.Y(n_1013)
);

NAND5xp2_ASAP7_75t_L g1014 ( 
.A(n_1006),
.B(n_813),
.C(n_839),
.D(n_842),
.E(n_872),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_1006),
.B(n_703),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1006),
.B(n_888),
.Y(n_1016)
);

AOI321xp33_ASAP7_75t_L g1017 ( 
.A1(n_1009),
.A2(n_861),
.A3(n_838),
.B1(n_843),
.B2(n_810),
.C(n_872),
.Y(n_1017)
);

AOI222xp33_ASAP7_75t_L g1018 ( 
.A1(n_1009),
.A2(n_739),
.B1(n_728),
.B2(n_823),
.C1(n_836),
.C2(n_851),
.Y(n_1018)
);

AOI221xp5_ASAP7_75t_L g1019 ( 
.A1(n_1006),
.A2(n_858),
.B1(n_701),
.B2(n_707),
.C(n_897),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_707),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1012),
.B(n_895),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_1014),
.A2(n_858),
.B(n_861),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_901),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_1016),
.B(n_865),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_1011),
.A2(n_1018),
.B(n_1010),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1013),
.B(n_1017),
.Y(n_1026)
);

AOI222xp33_ASAP7_75t_L g1027 ( 
.A1(n_1012),
.A2(n_823),
.B1(n_836),
.B2(n_829),
.C1(n_851),
.C2(n_839),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_1015),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_1020),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1024),
.B(n_903),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1021),
.Y(n_1031)
);

AND3x4_ASAP7_75t_L g1032 ( 
.A(n_1025),
.B(n_838),
.C(n_843),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1026),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_901),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_1023),
.B(n_834),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_1022),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1027),
.A2(n_764),
.B(n_772),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_1025),
.B(n_775),
.C(n_779),
.Y(n_1038)
);

NOR4xp75_ASAP7_75t_L g1039 ( 
.A(n_1025),
.B(n_810),
.C(n_180),
.D(n_181),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_1028),
.B(n_707),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_1020),
.A2(n_782),
.B(n_845),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_1039),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1036),
.B(n_1035),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_1029),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1030),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1033),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_1031),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_1034),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1032),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1047),
.Y(n_1051)
);

OA22x2_ASAP7_75t_L g1052 ( 
.A1(n_1045),
.A2(n_1038),
.B1(n_1041),
.B2(n_1037),
.Y(n_1052)
);

AO22x2_ASAP7_75t_L g1053 ( 
.A1(n_1042),
.A2(n_885),
.B1(n_903),
.B2(n_899),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_L g1054 ( 
.A(n_1046),
.B(n_701),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1043),
.Y(n_1055)
);

OA22x2_ASAP7_75t_L g1056 ( 
.A1(n_1048),
.A2(n_899),
.B1(n_892),
.B2(n_887),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1044),
.B(n_729),
.Y(n_1057)
);

XNOR2x2_ASAP7_75t_SL g1058 ( 
.A(n_1051),
.B(n_1050),
.Y(n_1058)
);

AND3x4_ASAP7_75t_L g1059 ( 
.A(n_1052),
.B(n_1049),
.C(n_1054),
.Y(n_1059)
);

OAI221xp5_ASAP7_75t_L g1060 ( 
.A1(n_1055),
.A2(n_712),
.B1(n_774),
.B2(n_875),
.C(n_900),
.Y(n_1060)
);

INVxp67_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1061),
.Y(n_1062)
);

XOR2xp5_ASAP7_75t_L g1063 ( 
.A(n_1062),
.B(n_1057),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1063),
.A2(n_1059),
.B1(n_1053),
.B2(n_1060),
.Y(n_1064)
);

OAI322xp33_ASAP7_75t_L g1065 ( 
.A1(n_1063),
.A2(n_1056),
.A3(n_875),
.B1(n_185),
.B2(n_186),
.C1(n_187),
.C2(n_191),
.Y(n_1065)
);

OR3x2_ASAP7_75t_L g1066 ( 
.A(n_1064),
.B(n_179),
.C(n_183),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_R g1067 ( 
.A1(n_1065),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1066),
.A2(n_712),
.B1(n_774),
.B2(n_887),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_SL g1069 ( 
.A1(n_1067),
.A2(n_195),
.B1(n_730),
.B2(n_712),
.Y(n_1069)
);

AO21x1_ASAP7_75t_L g1070 ( 
.A1(n_1068),
.A2(n_829),
.B(n_842),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_1069),
.A2(n_836),
.B(n_823),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1071),
.A2(n_840),
.B(n_892),
.Y(n_1072)
);

AOI211xp5_ASAP7_75t_L g1073 ( 
.A1(n_1072),
.A2(n_1070),
.B(n_831),
.C(n_830),
.Y(n_1073)
);


endmodule