module fake_jpeg_30377_n_529 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_529);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_529;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_57),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_59),
.Y(n_121)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_68),
.Y(n_118)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g125 ( 
.A(n_70),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_75),
.B(n_79),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_52),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_87),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_46),
.Y(n_117)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_95),
.B(n_99),
.Y(n_158)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_12),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_100),
.B(n_102),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_0),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_49),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_38),
.B1(n_44),
.B2(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_109),
.A2(n_111),
.B1(n_120),
.B2(n_140),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_110),
.B(n_132),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_38),
.B1(n_51),
.B2(n_34),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_40),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_17),
.B1(n_25),
.B2(n_40),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g124 ( 
.A(n_53),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_136),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_55),
.B(n_34),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_59),
.Y(n_138)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_54),
.A2(n_17),
.B1(n_25),
.B2(n_34),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_165),
.Y(n_191)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_73),
.A2(n_25),
.B1(n_17),
.B2(n_43),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_159),
.B1(n_97),
.B2(n_84),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_73),
.A2(n_43),
.B1(n_36),
.B2(n_50),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_70),
.Y(n_163)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_69),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_146),
.B(n_158),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_167),
.A2(n_183),
.B(n_145),
.Y(n_226)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_112),
.B(n_78),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_174),
.C(n_133),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_96),
.C(n_64),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_175),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_176),
.Y(n_235)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_181),
.B(n_206),
.Y(n_257)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_90),
.B(n_91),
.Y(n_183)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_125),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_185),
.A2(n_133),
.B1(n_145),
.B2(n_76),
.Y(n_249)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_30),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_195),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_134),
.A2(n_81),
.B1(n_83),
.B2(n_41),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_36),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_218),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_125),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_46),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_196),
.B(n_208),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_134),
.A2(n_81),
.B1(n_83),
.B2(n_41),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_111),
.A2(n_33),
.B1(n_20),
.B2(n_50),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_155),
.A2(n_33),
.B1(n_20),
.B2(n_67),
.Y(n_201)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_116),
.B(n_118),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_70),
.B(n_43),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_35),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_35),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_160),
.B(n_37),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_147),
.Y(n_213)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

CKINVDCx12_ASAP7_75t_R g214 ( 
.A(n_125),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_231)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_216),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_128),
.A2(n_101),
.B1(n_98),
.B2(n_63),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_173),
.B(n_123),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_224),
.B(n_255),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_167),
.B(n_37),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_225),
.B(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_226),
.A2(n_238),
.B1(n_240),
.B2(n_249),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_191),
.B(n_127),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_250),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_215),
.A2(n_157),
.B1(n_135),
.B2(n_93),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_171),
.A2(n_130),
.B1(n_162),
.B2(n_161),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_173),
.B(n_215),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_253),
.C(n_168),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_174),
.A2(n_194),
.B(n_188),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_203),
.A2(n_138),
.B1(n_148),
.B2(n_107),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_254),
.A2(n_199),
.B1(n_205),
.B2(n_107),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_135),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_203),
.B(n_127),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_259),
.B(n_178),
.Y(n_277)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_202),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_269),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_200),
.C(n_182),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_212),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_204),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_275),
.B(n_276),
.Y(n_328)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_277),
.B(n_287),
.Y(n_329)
);

OR2x4_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_163),
.Y(n_278)
);

NAND2x1_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_290),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_177),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_292),
.B(n_298),
.Y(n_309)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_285),
.B1(n_252),
.B2(n_235),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_222),
.B(n_189),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_226),
.A2(n_172),
.B1(n_218),
.B2(n_209),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_283),
.B1(n_261),
.B2(n_256),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_249),
.A2(n_130),
.B1(n_108),
.B2(n_162),
.Y(n_283)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_284),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.Y(n_301)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_187),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_244),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_256),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_170),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_296),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_239),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_295),
.B(n_221),
.Y(n_322)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_294),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_186),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_299),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_259),
.B(n_236),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_303),
.B(n_313),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_245),
.B1(n_240),
.B2(n_238),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_323),
.B1(n_331),
.B2(n_332),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_306),
.A2(n_315),
.B(n_316),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_270),
.A2(n_255),
.B(n_222),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_239),
.B(n_253),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_292),
.A2(n_277),
.B(n_278),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_322),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_223),
.B(n_229),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_319),
.B(n_324),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_229),
.B1(n_241),
.B2(n_244),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_320),
.A2(n_327),
.B1(n_297),
.B2(n_275),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_265),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_298),
.C(n_263),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_290),
.A2(n_231),
.B1(n_161),
.B2(n_108),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_242),
.B(n_233),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_241),
.B1(n_244),
.B2(n_141),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_281),
.B(n_242),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_330),
.B(n_264),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_279),
.A2(n_139),
.B1(n_115),
.B2(n_141),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_279),
.A2(n_139),
.B1(n_115),
.B2(n_219),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_298),
.B1(n_290),
.B2(n_291),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_333),
.A2(n_311),
.B(n_318),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_247),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_334),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_290),
.Y(n_337)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_247),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_342),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_357),
.C(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_312),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_364),
.B1(n_304),
.B2(n_308),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_311),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_299),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_284),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_352),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_350),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_305),
.A2(n_288),
.B1(n_287),
.B2(n_276),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_351),
.A2(n_310),
.B1(n_251),
.B2(n_269),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_280),
.Y(n_353)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_319),
.B(n_233),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_359),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_300),
.C(n_316),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_296),
.Y(n_358)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_237),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_314),
.B(n_237),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_360),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_320),
.B(n_243),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_363),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_321),
.B(n_251),
.C(n_216),
.Y(n_362)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_315),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_313),
.A2(n_303),
.B1(n_327),
.B2(n_302),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_317),
.C(n_304),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_175),
.C(n_190),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_335),
.A2(n_304),
.B1(n_332),
.B2(n_331),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_372),
.A2(n_383),
.B(n_384),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_373),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_243),
.Y(n_376)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_387),
.Y(n_398)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_301),
.Y(n_379)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_357),
.B(n_301),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_381),
.B(n_362),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_308),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_381),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_335),
.A2(n_299),
.B(n_312),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_336),
.B(n_318),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_385),
.B(n_388),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_335),
.A2(n_306),
.B(n_310),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_386),
.A2(n_390),
.B(n_333),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_358),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_340),
.B(n_285),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_397),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_176),
.B(n_178),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_351),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_289),
.Y(n_394)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_394),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_347),
.A2(n_268),
.B1(n_66),
.B2(n_86),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_401),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_386),
.B(n_391),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_368),
.B(n_344),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_405),
.B(n_413),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_343),
.C(n_354),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_406),
.B(n_416),
.C(n_417),
.Y(n_441)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_385),
.Y(n_409)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_348),
.Y(n_410)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_355),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_414),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_367),
.B(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_373),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_419),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_392),
.B(n_354),
.C(n_355),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_337),
.C(n_364),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_393),
.B(n_359),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_380),
.B(n_338),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_423),
.Y(n_435)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_339),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_425),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_383),
.B(n_339),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_384),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_426),
.B(n_438),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_399),
.A2(n_372),
.B1(n_391),
.B2(n_366),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_430),
.A2(n_403),
.B1(n_418),
.B2(n_420),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_422),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_437),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_409),
.A2(n_374),
.B1(n_402),
.B2(n_396),
.Y(n_436)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_436),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_410),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_399),
.A2(n_338),
.B(n_370),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_439),
.B(n_448),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_388),
.C(n_369),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_444),
.C(n_445),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_371),
.C(n_395),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_371),
.C(n_395),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_415),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_419),
.C(n_425),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_414),
.A2(n_396),
.B1(n_380),
.B2(n_370),
.Y(n_447)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_404),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_375),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_453),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_444),
.B(n_411),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_457),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_424),
.C(n_398),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_465),
.C(n_446),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_434),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_458),
.B(n_459),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_430),
.A2(n_421),
.B1(n_387),
.B2(n_398),
.Y(n_459)
);

OA22x2_ASAP7_75t_L g461 ( 
.A1(n_443),
.A2(n_349),
.B1(n_408),
.B2(n_397),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_466),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_428),
.B(n_412),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_463),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_440),
.A2(n_407),
.B1(n_390),
.B2(n_346),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_464),
.A2(n_432),
.B1(n_426),
.B2(n_438),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_389),
.C(n_407),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_440),
.A2(n_72),
.B1(n_179),
.B2(n_169),
.Y(n_466)
);

AO221x1_ASAP7_75t_L g467 ( 
.A1(n_431),
.A2(n_169),
.B1(n_179),
.B2(n_180),
.C(n_156),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_467),
.A2(n_434),
.B(n_435),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_473),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_451),
.A2(n_439),
.B(n_443),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_471),
.A2(n_466),
.B(n_1),
.Y(n_497)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_472),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_445),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_449),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_482),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_435),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_481),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_459),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_429),
.C(n_432),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_484),
.C(n_462),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_450),
.A2(n_429),
.B1(n_427),
.B2(n_94),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_427),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_18),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_461),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_18),
.C(n_1),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_486),
.B(n_496),
.Y(n_508)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_474),
.B(n_469),
.Y(n_487)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_487),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_493),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_475),
.B(n_460),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_464),
.C(n_461),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_498),
.C(n_499),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_476),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_497),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_18),
.C(n_1),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_0),
.C(n_2),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_494),
.A2(n_479),
.B(n_484),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_501),
.A2(n_507),
.B(n_485),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_489),
.B(n_482),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_506),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_490),
.B(n_0),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_492),
.A2(n_2),
.B(n_3),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_2),
.C(n_4),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_4),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_511),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_509),
.A2(n_486),
.B1(n_499),
.B2(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_513),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_488),
.C(n_6),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_516),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_501),
.B(n_8),
.C(n_9),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_SL g521 ( 
.A(n_517),
.B(n_503),
.C(n_505),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_500),
.Y(n_523)
);

AOI322xp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_500),
.A3(n_515),
.B1(n_514),
.B2(n_510),
.C1(n_8),
.C2(n_10),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_522),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_523),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_518),
.C(n_519),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_524),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_9),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_10),
.B(n_385),
.Y(n_529)
);


endmodule