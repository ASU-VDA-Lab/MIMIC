module fake_netlist_1_9414_n_580 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_580);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_580;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_472;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g72 ( .A(n_55), .Y(n_72) );
CKINVDCx20_ASAP7_75t_R g73 ( .A(n_24), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_18), .Y(n_74) );
BUFx2_ASAP7_75t_L g75 ( .A(n_63), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_68), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_34), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_44), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_64), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_6), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_22), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_49), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_69), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_12), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_0), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_43), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_10), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_54), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_60), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_62), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_17), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_67), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_17), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_51), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_25), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_12), .B(n_5), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_15), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_1), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_114), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_73), .Y(n_118) );
NOR2xp33_ASAP7_75t_R g119 ( .A(n_73), .B(n_32), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_78), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_83), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_78), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_75), .B(n_0), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_107), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_107), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_114), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_108), .B(n_1), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_93), .B(n_3), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_91), .Y(n_132) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_83), .A2(n_36), .B(n_66), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_76), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_98), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_92), .B(n_74), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_77), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_112), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_79), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_72), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_90), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_94), .B(n_4), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_86), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_88), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_92), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g149 ( .A1(n_106), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_90), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_121), .B(n_104), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
OR2x2_ASAP7_75t_SL g161 ( .A(n_130), .B(n_74), .Y(n_161) );
NAND2x1p5_ASAP7_75t_L g162 ( .A(n_116), .B(n_101), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_129), .A2(n_115), .B1(n_113), .B2(n_95), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_121), .B(n_102), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_151), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_138), .B(n_80), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_116), .B(n_80), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_122), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_123), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_132), .B(n_109), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_136), .B(n_105), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_122), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_122), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_122), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_135), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_122), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_139), .B(n_103), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_150), .B(n_111), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_126), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_137), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_124), .B(n_82), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_124), .B(n_82), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_150), .B(n_111), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_134), .B(n_110), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_140), .A2(n_100), .B1(n_96), .B2(n_90), .Y(n_194) );
NAND3x1_ASAP7_75t_L g195 ( .A(n_131), .B(n_7), .C(n_8), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
BUFx4f_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_118), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_143), .B(n_153), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_152), .B(n_85), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_153), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_201), .B(n_141), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_179), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_160), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_200), .B(n_146), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_201), .B(n_147), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_187), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
INVx3_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_203), .B(n_145), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_197), .B(n_119), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_203), .B(n_148), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_185), .B(n_125), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_155), .B(n_90), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_199), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_155), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_165), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_200), .B(n_127), .Y(n_221) );
OR2x6_ASAP7_75t_L g222 ( .A(n_195), .B(n_149), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_197), .B(n_133), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_167), .B(n_120), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_168), .B(n_128), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_168), .B(n_90), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_172), .A2(n_87), .B(n_72), .C(n_142), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_167), .B(n_7), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_187), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_179), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_189), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_158), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_189), .B(n_133), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_167), .B(n_8), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_159), .Y(n_238) );
AND3x1_ASAP7_75t_SL g239 ( .A(n_161), .B(n_149), .C(n_11), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_180), .Y(n_240) );
OR2x6_ASAP7_75t_L g241 ( .A(n_195), .B(n_87), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_189), .B(n_87), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_180), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_157), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_197), .B(n_87), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_162), .B(n_87), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_162), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_186), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_193), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_158), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_183), .B(n_72), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_173), .B(n_72), .Y(n_254) );
AO22x1_ASAP7_75t_L g255 ( .A1(n_158), .A2(n_142), .B1(n_11), .B2(n_14), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_161), .A2(n_142), .B1(n_14), .B2(n_15), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_192), .B(n_9), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_229), .A2(n_158), .B1(n_164), .B2(n_162), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_236), .A2(n_193), .B(n_196), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_208), .B(n_192), .Y(n_261) );
INVx2_ASAP7_75t_R g262 ( .A(n_210), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_247), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_204), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_208), .B(n_202), .Y(n_265) );
BUFx3_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
NOR2xp67_ASAP7_75t_L g267 ( .A(n_225), .B(n_193), .Y(n_267) );
OA22x2_ASAP7_75t_L g268 ( .A1(n_222), .A2(n_163), .B1(n_190), .B2(n_191), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_230), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_257), .B(n_191), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g272 ( .A1(n_246), .A2(n_174), .B(n_175), .C(n_184), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_247), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_231), .B(n_164), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_244), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_247), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_234), .B(n_213), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_248), .B(n_164), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_249), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_220), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_252), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_229), .B(n_164), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_205), .B(n_164), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_209), .B(n_164), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_SL g289 ( .A1(n_243), .A2(n_194), .B(n_166), .C(n_154), .Y(n_289) );
NOR2xp33_ASAP7_75t_SL g290 ( .A(n_245), .B(n_159), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_215), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_227), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_229), .B(n_159), .Y(n_293) );
NAND2x1_ASAP7_75t_L g294 ( .A(n_206), .B(n_154), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_242), .B(n_166), .Y(n_295) );
BUFx10_ASAP7_75t_L g296 ( .A(n_237), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_245), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_237), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_237), .B(n_9), .Y(n_300) );
INVx6_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_268), .A2(n_222), .B1(n_207), .B2(n_257), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_291), .B(n_207), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_261), .B(n_226), .Y(n_306) );
NAND3xp33_ASAP7_75t_SL g307 ( .A(n_283), .B(n_218), .C(n_256), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_263), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_268), .A2(n_222), .B1(n_241), .B2(n_221), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_259), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_291), .B(n_224), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_270), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_300), .A2(n_284), .B(n_282), .C(n_292), .Y(n_313) );
CKINVDCx6p67_ASAP7_75t_R g314 ( .A(n_266), .Y(n_314) );
BUFx8_ASAP7_75t_SL g315 ( .A(n_297), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_268), .A2(n_222), .B1(n_241), .B2(n_217), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_269), .B(n_251), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_300), .A2(n_241), .B1(n_219), .B2(n_223), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_288), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_269), .B(n_251), .Y(n_322) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_299), .A2(n_241), .B1(n_239), .B2(n_211), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_260), .A2(n_223), .B(n_250), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_261), .B(n_282), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_297), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_265), .B(n_224), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_300), .Y(n_328) );
OAI211xp5_ASAP7_75t_L g329 ( .A1(n_309), .A2(n_216), .B(n_265), .C(n_218), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_328), .A2(n_299), .B1(n_290), .B2(n_296), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_323), .A2(n_285), .B1(n_293), .B2(n_296), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
OAI21x1_ASAP7_75t_SL g333 ( .A1(n_319), .A2(n_258), .B(n_277), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_323), .A2(n_285), .B1(n_293), .B2(n_271), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_328), .B(n_270), .Y(n_335) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_319), .A2(n_286), .B(n_287), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_306), .A2(n_285), .B1(n_293), .B2(n_271), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_311), .A2(n_278), .B1(n_263), .B2(n_266), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_306), .A2(n_284), .B1(n_292), .B2(n_280), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_327), .A2(n_272), .B1(n_289), .B2(n_275), .C(n_277), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_311), .B(n_275), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_305), .B(n_262), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_327), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_273), .B1(n_253), .B2(n_263), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_326), .Y(n_350) );
OAI221xp5_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_274), .B1(n_281), .B2(n_254), .C(n_238), .Y(n_351) );
OAI221xp5_ASAP7_75t_L g352 ( .A1(n_304), .A2(n_238), .B1(n_273), .B2(n_267), .C(n_214), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_348), .B(n_346), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_329), .B(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_338), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_334), .A2(n_309), .B1(n_317), .B2(n_325), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_333), .B(n_313), .Y(n_358) );
NOR3xp33_ASAP7_75t_SL g359 ( .A(n_352), .B(n_307), .C(n_315), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_338), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_350), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_346), .B(n_312), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_341), .A2(n_317), .B(n_228), .C(n_308), .Y(n_363) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_337), .B(n_307), .C(n_217), .D(n_267), .Y(n_364) );
AOI33xp33_ASAP7_75t_L g365 ( .A1(n_340), .A2(n_217), .A3(n_170), .B1(n_169), .B2(n_19), .B3(n_16), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_343), .B(n_301), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_343), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_345), .B(n_301), .Y(n_369) );
NAND3xp33_ASAP7_75t_SL g370 ( .A(n_330), .B(n_211), .C(n_235), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
NOR4xp25_ASAP7_75t_SL g372 ( .A(n_352), .B(n_255), .C(n_235), .D(n_314), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_347), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_347), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_331), .A2(n_314), .B1(n_301), .B2(n_278), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_333), .A2(n_314), .B1(n_301), .B2(n_278), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_332), .A2(n_324), .B(n_321), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_335), .B(n_308), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_332), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_351), .A2(n_301), .B1(n_322), .B2(n_318), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_335), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_308), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_373), .B(n_351), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_367), .Y(n_388) );
NAND3xp33_ASAP7_75t_L g389 ( .A(n_359), .B(n_342), .C(n_349), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_367), .Y(n_390) );
OAI33xp33_ASAP7_75t_L g391 ( .A1(n_356), .A2(n_339), .A3(n_19), .B1(n_16), .B2(n_170), .B3(n_169), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_354), .B(n_342), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_383), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_383), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_384), .B(n_308), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_376), .B(n_302), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_381), .B(n_302), .Y(n_398) );
AOI31xp33_ASAP7_75t_L g399 ( .A1(n_355), .A2(n_223), .A3(n_336), .B(n_322), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_374), .B(n_316), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_379), .B(n_320), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_355), .A2(n_357), .B1(n_382), .B2(n_375), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_360), .B(n_321), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_368), .B(n_321), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_371), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_365), .B(n_336), .C(n_324), .D(n_238), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_378), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_362), .B(n_320), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_358), .B(n_320), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_385), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_365), .B(n_316), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_369), .B(n_316), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_358), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_358), .B(n_262), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
OAI33xp33_ASAP7_75t_L g419 ( .A1(n_363), .A2(n_176), .A3(n_171), .B1(n_177), .B2(n_178), .B3(n_182), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_361), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_366), .B(n_262), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_369), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_364), .Y(n_424) );
AND2x4_ASAP7_75t_SL g425 ( .A(n_370), .B(n_263), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_372), .B(n_255), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_373), .B(n_276), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_424), .A2(n_278), .B1(n_322), .B2(n_318), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_424), .A2(n_278), .B1(n_318), .B2(n_322), .Y(n_432) );
NOR4xp25_ASAP7_75t_SL g433 ( .A(n_390), .B(n_295), .C(n_23), .D(n_26), .Y(n_433) );
NAND2xp33_ASAP7_75t_SL g434 ( .A(n_390), .B(n_322), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_388), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_412), .B(n_318), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_407), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_420), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_412), .B(n_318), .Y(n_441) );
OAI33xp33_ASAP7_75t_L g442 ( .A1(n_402), .A2(n_177), .A3(n_188), .B1(n_182), .B2(n_178), .B3(n_171), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_393), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_388), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_393), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_389), .A2(n_294), .B(n_264), .C(n_298), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_394), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_409), .B(n_233), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_413), .B(n_21), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_409), .B(n_279), .Y(n_452) );
NOR3xp33_ASAP7_75t_SL g453 ( .A(n_389), .B(n_27), .C(n_29), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_427), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_392), .B(n_233), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_388), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_416), .B(n_30), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_403), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_33), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g464 ( .A1(n_399), .A2(n_298), .B(n_279), .Y(n_464) );
OAI322xp33_ASAP7_75t_L g465 ( .A1(n_386), .A2(n_294), .A3(n_176), .B1(n_188), .B2(n_232), .C1(n_250), .C2(n_233), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_422), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_411), .B(n_37), .Y(n_467) );
BUFx12f_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_386), .B(n_276), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_417), .A2(n_288), .B(n_298), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g473 ( .A(n_417), .B(n_288), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_404), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_418), .B(n_219), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_40), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_464), .B(n_425), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_459), .B(n_408), .Y(n_479) );
AOI222xp33_ASAP7_75t_L g480 ( .A1(n_470), .A2(n_423), .B1(n_391), .B2(n_418), .C1(n_425), .C2(n_395), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_444), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_460), .B(n_410), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g483 ( .A(n_453), .B(n_426), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_468), .A2(n_406), .B1(n_419), .B2(n_425), .Y(n_486) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_435), .A2(n_414), .B(n_426), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_443), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_435), .B(n_400), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_440), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_461), .B(n_428), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_474), .B(n_408), .Y(n_495) );
NAND3xp33_ASAP7_75t_SL g496 ( .A(n_440), .B(n_415), .C(n_421), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_466), .B(n_400), .Y(n_497) );
NOR2xp33_ASAP7_75t_SL g498 ( .A(n_468), .B(n_398), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_466), .B(n_398), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_462), .B(n_396), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_434), .A2(n_396), .B1(n_401), .B2(n_264), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_432), .A2(n_401), .B1(n_264), .B2(n_250), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_434), .B(n_401), .Y(n_503) );
OAI211xp5_ASAP7_75t_L g504 ( .A1(n_472), .A2(n_250), .B(n_233), .C(n_232), .Y(n_504) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_450), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_447), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_452), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_446), .A2(n_401), .B(n_212), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_448), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_449), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_442), .A2(n_232), .B1(n_206), .B2(n_233), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_436), .A2(n_41), .B(n_42), .C(n_45), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g515 ( .A(n_433), .B(n_46), .C(n_47), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_469), .B(n_232), .Y(n_516) );
XNOR2xp5_ASAP7_75t_L g517 ( .A(n_492), .B(n_476), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_484), .Y(n_518) );
INVxp33_ASAP7_75t_L g519 ( .A(n_478), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_481), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_512), .B(n_471), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_507), .B(n_471), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_490), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_478), .A2(n_473), .B(n_465), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_485), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_489), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_498), .A2(n_467), .B1(n_441), .B2(n_430), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_479), .B(n_495), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_494), .B(n_451), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_506), .Y(n_532) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_496), .B(n_454), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_479), .B(n_455), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_495), .B(n_451), .Y(n_535) );
AOI31xp33_ASAP7_75t_L g536 ( .A1(n_503), .A2(n_463), .A3(n_458), .B(n_475), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_505), .B(n_463), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_509), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_510), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_482), .B(n_475), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_500), .B(n_232), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_493), .B(n_50), .Y(n_543) );
AOI222xp33_ASAP7_75t_L g544 ( .A1(n_519), .A2(n_483), .B1(n_486), .B2(n_499), .C1(n_515), .C2(n_516), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_527), .Y(n_545) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_517), .B(n_497), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_520), .B(n_490), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_524), .A2(n_504), .B(n_483), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_519), .A2(n_486), .B1(n_480), .B2(n_487), .C(n_501), .Y(n_549) );
OAI21xp5_ASAP7_75t_SL g550 ( .A1(n_517), .A2(n_502), .B(n_508), .Y(n_550) );
INVxp33_ASAP7_75t_L g551 ( .A(n_530), .Y(n_551) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_523), .Y(n_552) );
XOR2x2_ASAP7_75t_L g553 ( .A(n_528), .B(n_513), .Y(n_553) );
OAI211xp5_ASAP7_75t_SL g554 ( .A1(n_541), .A2(n_513), .B(n_514), .C(n_511), .Y(n_554) );
OAI222xp33_ASAP7_75t_L g555 ( .A1(n_530), .A2(n_514), .B1(n_53), .B2(n_56), .C1(n_57), .C2(n_59), .Y(n_555) );
OAI31xp33_ASAP7_75t_SL g556 ( .A1(n_552), .A2(n_536), .A3(n_533), .B(n_518), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_553), .A2(n_534), .B1(n_537), .B2(n_540), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_548), .B(n_540), .C(n_527), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_549), .A2(n_535), .B1(n_542), .B2(n_538), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_545), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_550), .A2(n_525), .B1(n_532), .B2(n_531), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_546), .A2(n_529), .B1(n_522), .B2(n_526), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_548), .B(n_543), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_544), .B(n_521), .C(n_539), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_551), .B(n_61), .Y(n_565) );
OAI321xp33_ASAP7_75t_L g566 ( .A1(n_549), .A2(n_156), .A3(n_198), .B1(n_65), .B2(n_70), .C(n_204), .Y(n_566) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_554), .A2(n_156), .B(n_198), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_554), .B(n_555), .C(n_547), .Y(n_568) );
OAI311xp33_ASAP7_75t_L g569 ( .A1(n_555), .A2(n_544), .A3(n_550), .B1(n_549), .C1(n_480), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_564), .A2(n_568), .B1(n_563), .B2(n_559), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_560), .Y(n_571) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_561), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_562), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_573), .B(n_564), .C(n_566), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_570), .A2(n_556), .B1(n_558), .B2(n_557), .C(n_569), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_575), .B(n_572), .Y(n_576) );
NOR3xp33_ASAP7_75t_L g577 ( .A(n_574), .B(n_567), .C(n_565), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_578), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_579), .A2(n_577), .B(n_571), .Y(n_580) );
endmodule