module fake_aes_7062_n_15 (n_3, n_1, n_2, n_0, n_15);
input n_3;
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_3), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
CKINVDCx5p33_ASAP7_75t_R g6 ( .A(n_2), .Y(n_6) );
BUFx6f_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_4), .B(n_0), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_8), .B(n_6), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_12), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_13), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
endmodule