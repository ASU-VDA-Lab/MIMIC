module fake_jpeg_20635_n_289 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_13),
.B(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_44),
.B1(n_21),
.B2(n_34),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_28),
.C(n_26),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_21),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_21),
.B(n_17),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_59),
.C(n_27),
.Y(n_86)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_62),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_46),
.B(n_37),
.C(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_12),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_55),
.B1(n_63),
.B2(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_13),
.Y(n_88)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_20),
.B1(n_23),
.B2(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_15),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_18),
.B(n_15),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_29),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_31),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_16),
.B(n_18),
.C(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_24),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_84),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_85),
.B(n_60),
.C(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_51),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_55),
.B1(n_49),
.B2(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_59),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_102),
.B1(n_105),
.B2(n_104),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_22),
.B1(n_14),
.B2(n_2),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_58),
.B(n_49),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_107),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_62),
.B1(n_65),
.B2(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_77),
.B1(n_76),
.B2(n_62),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_59),
.B1(n_57),
.B2(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_76),
.B1(n_68),
.B2(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_35),
.B1(n_38),
.B2(n_59),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_38),
.B1(n_66),
.B2(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_12),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_25),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_116),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_81),
.B1(n_82),
.B2(n_74),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_120),
.B1(n_90),
.B2(n_100),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_70),
.B(n_78),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_130),
.B(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_70),
.B(n_88),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_96),
.B(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_80),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_72),
.B1(n_38),
.B2(n_69),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_72),
.B1(n_77),
.B2(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_68),
.B1(n_18),
.B2(n_16),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_16),
.B1(n_13),
.B2(n_29),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_12),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_135),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_22),
.B1(n_14),
.B2(n_7),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_22),
.B1(n_14),
.B2(n_7),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_22),
.C(n_14),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_102),
.C(n_105),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_92),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_153),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_150),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_135),
.B(n_6),
.Y(n_180)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_96),
.B(n_92),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_124),
.B(n_127),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_131),
.B1(n_130),
.B2(n_135),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_5),
.B(n_10),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_135),
.C(n_14),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_158),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_93),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_109),
.B1(n_106),
.B2(n_91),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_157),
.B1(n_4),
.B2(n_9),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_99),
.B1(n_90),
.B2(n_108),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_22),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_121),
.B1(n_123),
.B2(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_133),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_110),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_178),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_185),
.B1(n_190),
.B2(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_188),
.B1(n_165),
.B2(n_142),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_181),
.B(n_186),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_126),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_191),
.C(n_186),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_163),
.B1(n_162),
.B2(n_159),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_6),
.B(n_10),
.Y(n_181)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_5),
.B1(n_10),
.B2(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_164),
.B1(n_155),
.B2(n_154),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_7),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_201),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_154),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_206),
.B(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_140),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_146),
.B1(n_149),
.B2(n_136),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_204),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_166),
.B1(n_180),
.B2(n_191),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_187),
.B(n_157),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_160),
.B1(n_139),
.B2(n_2),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_139),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_176),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_0),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_0),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_179),
.C(n_173),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_215),
.C(n_226),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_178),
.C(n_168),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_221),
.B(n_206),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_227),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_228),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_181),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_203),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_170),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_177),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_229),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_199),
.B(n_198),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_224),
.B(n_198),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_196),
.B1(n_193),
.B2(n_200),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_195),
.B1(n_202),
.B2(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_212),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_172),
.B1(n_208),
.B2(n_171),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_215),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_213),
.C(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_251),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_234),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_238),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_227),
.C(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_174),
.C(n_205),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_255),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_205),
.B(n_183),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_231),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_263),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_263),
.B(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_264),
.B(n_265),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_7),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_0),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_248),
.B1(n_253),
.B2(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.Y(n_279)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_1),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_275),
.B(n_8),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_277),
.B(n_278),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_8),
.B(n_9),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_8),
.B(n_11),
.C(n_1),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_275),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_279),
.A2(n_274),
.B(n_272),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_269),
.B(n_270),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_267),
.C(n_283),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_285),
.C(n_11),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_2),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_288),
.Y(n_289)
);


endmodule