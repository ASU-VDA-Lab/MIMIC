module fake_jpeg_22944_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_5),
.B(n_2),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx12_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_6),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_18),
.B(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_27),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_19),
.B1(n_7),
.B2(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_23),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B(n_6),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_24),
.C(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_12),
.B(n_3),
.Y(n_36)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_34),
.C2(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_1),
.C(n_3),
.Y(n_40)
);


endmodule