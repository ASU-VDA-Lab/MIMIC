module fake_aes_2034_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_74), .Y(n_77) );
INVxp67_ASAP7_75t_L g78 ( .A(n_46), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_40), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_39), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_9), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
CKINVDCx14_ASAP7_75t_R g83 ( .A(n_55), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_5), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_8), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_51), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_41), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_28), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_37), .Y(n_90) );
NOR2xp67_ASAP7_75t_L g91 ( .A(n_13), .B(n_50), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_10), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_0), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_3), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_38), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_17), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_0), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_33), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_56), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_15), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_17), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_14), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_23), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_76), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_58), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_70), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_27), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_26), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_53), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_45), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_35), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_3), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_30), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_18), .B(n_6), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_85), .B(n_1), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_85), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_112), .B(n_2), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_112), .B(n_2), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_102), .Y(n_136) );
INVx5_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_94), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_102), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_92), .A2(n_34), .B(n_71), .Y(n_142) );
XNOR2xp5_ASAP7_75t_L g143 ( .A(n_105), .B(n_4), .Y(n_143) );
INVx5_ASAP7_75t_L g144 ( .A(n_94), .Y(n_144) );
INVxp67_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_110), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_83), .B(n_7), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_110), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_82), .B(n_8), .Y(n_149) );
INVx5_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
NAND2xp33_ASAP7_75t_SL g153 ( .A(n_80), .B(n_9), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_99), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_116), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_100), .Y(n_161) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_103), .A2(n_42), .B(n_69), .Y(n_162) );
INVxp67_ASAP7_75t_L g163 ( .A(n_98), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_84), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_107), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_106), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_136), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_143), .A2(n_81), .B1(n_117), .B2(n_121), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_145), .B(n_95), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_127), .A2(n_97), .B1(n_121), .B2(n_84), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_127), .B(n_118), .Y(n_171) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_147), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_137), .B(n_90), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_132), .B(n_111), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
OAI21xp33_ASAP7_75t_L g178 ( .A1(n_132), .A2(n_95), .B(n_86), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_131), .B(n_97), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
AO22x2_ASAP7_75t_L g181 ( .A1(n_131), .A2(n_86), .B1(n_93), .B2(n_123), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_160), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_161), .B(n_78), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_125), .B(n_93), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_160), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_137), .B(n_90), .Y(n_191) );
INVx6_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_161), .B(n_89), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_137), .B(n_114), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_137), .B(n_114), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_137), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_137), .B(n_119), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_137), .B(n_115), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_130), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_141), .B(n_91), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_147), .B(n_108), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
AND2x6_ASAP7_75t_L g204 ( .A(n_141), .B(n_101), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_146), .B(n_96), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_130), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_146), .B(n_12), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_150), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_130), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_163), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_211) );
NAND3x1_ASAP7_75t_L g212 ( .A(n_165), .B(n_140), .C(n_125), .Y(n_212) );
BUFx4_ASAP7_75t_L g213 ( .A(n_129), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_164), .B(n_16), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_130), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
INVx3_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_133), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_166), .B(n_18), .Y(n_223) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_151), .B(n_47), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_151), .B(n_19), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_158), .B(n_20), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_150), .B(n_21), .Y(n_227) );
OAI22xp33_ASAP7_75t_SL g228 ( .A1(n_165), .A2(n_22), .B1(n_24), .B2(n_25), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_183), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_204), .A2(n_202), .B1(n_189), .B2(n_181), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_215), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_190), .Y(n_233) );
AND2x4_ASAP7_75t_SL g234 ( .A(n_189), .B(n_140), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_192), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_185), .A2(n_142), .B(n_162), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_187), .Y(n_238) );
AND2x6_ASAP7_75t_L g239 ( .A(n_180), .B(n_154), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_190), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_204), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_189), .A2(n_126), .B1(n_153), .B2(n_158), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_167), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_189), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_201), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_216), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_181), .B(n_142), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_204), .A2(n_158), .B1(n_155), .B2(n_157), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_179), .B(n_138), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_179), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_229), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_179), .B(n_150), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_193), .B(n_150), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_193), .B(n_152), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_188), .B(n_154), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_222), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_226), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_188), .B(n_154), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_205), .B(n_152), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_202), .B(n_223), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_208), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_204), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_226), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_168), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_202), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_169), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_226), .Y(n_273) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_175), .B(n_162), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_222), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_199), .Y(n_276) );
OAI22xp5_ASAP7_75t_SL g277 ( .A1(n_212), .A2(n_162), .B1(n_138), .B2(n_156), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_202), .B(n_138), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_199), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_180), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_204), .A2(n_134), .B1(n_157), .B2(n_156), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_203), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_204), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_202), .B(n_138), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_225), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_192), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_195), .B(n_157), .Y(n_288) );
AOI22xp5_ASAP7_75t_SL g289 ( .A1(n_228), .A2(n_162), .B1(n_156), .B2(n_155), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_176), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_177), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_196), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_197), .B(n_155), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_198), .B(n_152), .Y(n_294) );
AOI22xp5_ASAP7_75t_SL g295 ( .A1(n_211), .A2(n_139), .B1(n_134), .B2(n_148), .Y(n_295) );
OAI22x1_ASAP7_75t_L g296 ( .A1(n_241), .A2(n_212), .B1(n_200), .B2(n_181), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_278), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_239), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_239), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_239), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_239), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_235), .B(n_170), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_272), .B(n_253), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_234), .B(n_170), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_239), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_231), .A2(n_171), .B1(n_174), .B2(n_178), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_242), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_230), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_234), .A2(n_171), .B1(n_174), .B2(n_191), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_245), .A2(n_191), .B1(n_200), .B2(n_194), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_232), .A2(n_173), .B1(n_139), .B2(n_196), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_238), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
OR2x6_ASAP7_75t_L g318 ( .A(n_268), .B(n_213), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_284), .B(n_224), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_239), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_244), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_233), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_253), .B(n_139), .Y(n_326) );
BUFx10_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_230), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_266), .B(n_128), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_266), .B(n_128), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_238), .Y(n_331) );
BUFx3_ASAP7_75t_L g332 ( .A(n_284), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_271), .Y(n_333) );
HAxp5_ASAP7_75t_L g334 ( .A(n_270), .B(n_144), .CON(n_334), .SN(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_248), .B(n_182), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_244), .A2(n_224), .B1(n_144), .B2(n_135), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_263), .Y(n_337) );
BUFx5_ASAP7_75t_L g338 ( .A(n_240), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_252), .B(n_144), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_252), .B(n_144), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_246), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g342 ( .A1(n_241), .A2(n_144), .B1(n_128), .B2(n_148), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_246), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_252), .B(n_144), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_254), .B(n_133), .Y(n_345) );
CKINVDCx11_ASAP7_75t_R g346 ( .A(n_325), .Y(n_346) );
AOI222xp33_ASAP7_75t_L g347 ( .A1(n_307), .A2(n_233), .B1(n_270), .B2(n_254), .C1(n_285), .C2(n_279), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_322), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_304), .B(n_266), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_316), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_322), .B(n_265), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_304), .B(n_243), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_318), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_341), .A2(n_257), .B1(n_273), .B2(n_290), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
NAND3x1_ASAP7_75t_L g357 ( .A(n_307), .B(n_251), .C(n_237), .Y(n_357) );
BUFx12f_ASAP7_75t_L g358 ( .A(n_318), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_311), .B(n_267), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_328), .B(n_286), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_296), .A2(n_279), .B1(n_285), .B2(n_271), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_345), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_305), .B(n_285), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_341), .A2(n_273), .B1(n_290), .B2(n_269), .Y(n_364) );
OR2x6_ASAP7_75t_L g365 ( .A(n_318), .B(n_263), .Y(n_365) );
INVx8_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_312), .A2(n_282), .B1(n_264), .B2(n_260), .C(n_295), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_318), .B(n_259), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_296), .B(n_291), .Y(n_369) );
INVx4_ASAP7_75t_L g370 ( .A(n_319), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_319), .B(n_273), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_332), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
CKINVDCx14_ASAP7_75t_R g375 ( .A(n_345), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_329), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_352), .A2(n_277), .B1(n_329), .B2(n_330), .C1(n_293), .C2(n_309), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_375), .A2(n_353), .B1(n_374), .B2(n_365), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_347), .A2(n_335), .B1(n_329), .B2(n_330), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_369), .A2(n_289), .B(n_250), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_359), .B(n_329), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_343), .B(n_316), .C(n_320), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_367), .A2(n_320), .B(n_314), .Y(n_384) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_365), .B(n_343), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_360), .A2(n_330), .B1(n_342), .B2(n_294), .C(n_326), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_348), .B(n_330), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_363), .B(n_343), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_349), .A2(n_262), .B1(n_288), .B2(n_148), .C(n_135), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_350), .A2(n_337), .B(n_331), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_358), .A2(n_250), .B1(n_338), .B2(n_332), .Y(n_395) );
OR2x6_ASAP7_75t_L g396 ( .A(n_366), .B(n_332), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_366), .A2(n_250), .B1(n_338), .B2(n_269), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_346), .B(n_327), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_362), .B(n_331), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_370), .B(n_365), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_366), .A2(n_250), .B1(n_263), .B2(n_269), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_376), .B(n_339), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_353), .A2(n_269), .B1(n_333), .B2(n_334), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_390), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_388), .B(n_368), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_366), .B1(n_361), .B2(n_365), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_381), .A2(n_372), .B(n_355), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_382), .B(n_374), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_400), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_382), .B(n_355), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_378), .A2(n_387), .B1(n_400), .B2(n_396), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_389), .A2(n_372), .B1(n_274), .B2(n_334), .C1(n_297), .C2(n_299), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_399), .B(n_334), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_385), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_378), .B(n_356), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_396), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g420 ( .A1(n_380), .A2(n_336), .B(n_356), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_384), .A2(n_357), .B(n_354), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_391), .B(n_297), .Y(n_423) );
OAI21x1_ASAP7_75t_L g424 ( .A1(n_397), .A2(n_357), .B(n_364), .Y(n_424) );
OR2x2_ASAP7_75t_SL g425 ( .A(n_401), .B(n_133), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_396), .A2(n_370), .B1(n_373), .B2(n_371), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_395), .B(n_370), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_402), .B(n_371), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_386), .B(n_371), .Y(n_429) );
AO22x1_ASAP7_75t_L g430 ( .A1(n_398), .A2(n_371), .B1(n_300), .B2(n_308), .Y(n_430) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_386), .A2(n_256), .B1(n_340), .B2(n_344), .C(n_255), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_403), .A2(n_338), .B1(n_269), .B2(n_299), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_381), .A2(n_338), .B1(n_337), .B2(n_300), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_393), .A2(n_333), .B1(n_300), .B2(n_308), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_401), .A2(n_338), .B1(n_337), .B2(n_300), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
OAI22xp5_ASAP7_75t_SL g437 ( .A1(n_378), .A2(n_274), .B1(n_298), .B2(n_301), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_390), .B(n_337), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_377), .A2(n_338), .B1(n_321), .B2(n_308), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_420), .A2(n_135), .B1(n_133), .B2(n_148), .C(n_302), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_404), .B(n_133), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g443 ( .A1(n_420), .A2(n_315), .B(n_302), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_411), .B(n_135), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_135), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_414), .B(n_135), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_425), .A2(n_301), .B1(n_298), .B2(n_321), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_413), .B(n_148), .C(n_217), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_406), .B(n_405), .C(n_426), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_408), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_429), .A2(n_148), .B1(n_317), .B2(n_323), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_323), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_417), .B(n_317), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_429), .B(n_323), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_439), .A2(n_321), .B(n_308), .C(n_333), .Y(n_457) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_430), .A2(n_321), .B(n_333), .C(n_227), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_417), .B(n_323), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_419), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_408), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_407), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_410), .B(n_323), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_407), .Y(n_467) );
AOI211xp5_ASAP7_75t_SL g468 ( .A1(n_437), .A2(n_306), .B(n_313), .C(n_324), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_410), .B(n_323), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_425), .A2(n_303), .B1(n_310), .B2(n_317), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_317), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_409), .B(n_317), .Y(n_472) );
OAI33xp33_ASAP7_75t_L g473 ( .A1(n_416), .A2(n_214), .A3(n_207), .B1(n_210), .B2(n_203), .B3(n_324), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_438), .B(n_338), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_438), .B(n_338), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_419), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_437), .A2(n_317), .B1(n_338), .B2(n_306), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_423), .B(n_313), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_428), .B(n_327), .Y(n_479) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_427), .B(n_327), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_407), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_436), .A2(n_310), .A3(n_303), .B(n_249), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
NOR3xp33_ASAP7_75t_SL g486 ( .A(n_431), .B(n_327), .C(n_292), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g487 ( .A1(n_421), .A2(n_258), .B1(n_249), .B2(n_247), .C1(n_303), .C2(n_310), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
AOI33xp33_ASAP7_75t_L g489 ( .A1(n_422), .A2(n_214), .A3(n_207), .B1(n_210), .B2(n_258), .B3(n_247), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_409), .B(n_29), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_451), .B(n_409), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_456), .B(n_415), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_440), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_440), .B(n_422), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_464), .B(n_424), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_455), .B(n_424), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_480), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_484), .B(n_453), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_453), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_454), .B(n_427), .Y(n_501) );
INVxp67_ASAP7_75t_L g502 ( .A(n_463), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_447), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_463), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_455), .B(n_415), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_442), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_470), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_450), .A2(n_427), .B1(n_436), .B2(n_434), .Y(n_508) );
OAI211xp5_ASAP7_75t_L g509 ( .A1(n_449), .A2(n_435), .B(n_432), .C(n_433), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_479), .B(n_430), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_447), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_476), .B(n_436), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_462), .B(n_217), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_471), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_217), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_471), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_462), .B(n_217), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_447), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_446), .B(n_32), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_446), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_481), .B(n_36), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_460), .Y(n_522) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_441), .B(n_220), .C(n_287), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_476), .Y(n_524) );
AND2x4_ASAP7_75t_SL g525 ( .A(n_491), .B(n_220), .Y(n_525) );
NAND5xp2_ASAP7_75t_L g526 ( .A(n_468), .B(n_43), .C(n_44), .D(n_48), .E(n_54), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_488), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_444), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_480), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_481), .B(n_57), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_460), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_480), .Y(n_532) );
BUFx2_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_444), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_445), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_466), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_465), .B(n_59), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_466), .B(n_60), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_465), .B(n_62), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_63), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_469), .B(n_64), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_459), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_459), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_467), .B(n_220), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_469), .B(n_67), .Y(n_546) );
XNOR2x1_ASAP7_75t_L g547 ( .A(n_449), .B(n_68), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_467), .B(n_72), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_499), .B(n_461), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_536), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_527), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_502), .B(n_486), .C(n_490), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_495), .B(n_467), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_537), .B(n_490), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_500), .B(n_461), .Y(n_557) );
BUFx3_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_514), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_547), .B(n_485), .C(n_482), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_496), .Y(n_561) );
XNOR2xp5_ASAP7_75t_L g562 ( .A(n_547), .B(n_470), .Y(n_562) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_526), .A2(n_443), .B(n_448), .C(n_487), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_511), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_505), .B(n_485), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_510), .B(n_491), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_495), .B(n_461), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_504), .B(n_456), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_543), .A2(n_473), .B1(n_478), .B2(n_477), .C(n_475), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_524), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_524), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_544), .B(n_482), .Y(n_572) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_498), .B(n_491), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_529), .A2(n_474), .B1(n_491), .B2(n_456), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_516), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_520), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_506), .B(n_489), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_505), .B(n_472), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_501), .B(n_472), .Y(n_579) );
AOI32xp33_ASAP7_75t_L g580 ( .A1(n_532), .A2(n_452), .A3(n_472), .B1(n_483), .B2(n_458), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_501), .B(n_472), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_496), .B(n_483), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_492), .B(n_457), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_529), .B(n_287), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_528), .B(n_275), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_497), .B(n_275), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_535), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_508), .B(n_236), .C(n_261), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_497), .B(n_261), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_512), .B(n_236), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_533), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_503), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_533), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_523), .B(n_236), .C(n_280), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_507), .A2(n_236), .B1(n_192), .B2(n_209), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_551), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_560), .B(n_525), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_551), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_565), .B(n_531), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_570), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_558), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_554), .B(n_509), .C(n_546), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g603 ( .A1(n_562), .A2(n_493), .B(n_542), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_571), .Y(n_604) );
AOI32xp33_ASAP7_75t_L g605 ( .A1(n_573), .A2(n_525), .A3(n_521), .B1(n_530), .B2(n_548), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_559), .B(n_518), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_568), .Y(n_607) );
XNOR2x2_ASAP7_75t_L g608 ( .A(n_588), .B(n_530), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_553), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_564), .Y(n_610) );
NOR2xp33_ASAP7_75t_R g611 ( .A(n_583), .B(n_521), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_582), .A2(n_539), .B1(n_519), .B2(n_515), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_575), .B(n_534), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_594), .B(n_548), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_549), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_580), .B(n_493), .C(n_541), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_563), .A2(n_541), .B(n_540), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_577), .A2(n_493), .B(n_515), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_578), .B(n_522), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_587), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_561), .B(n_522), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_564), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_578), .B(n_518), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_572), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_572), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_579), .B(n_540), .Y(n_627) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_563), .B(n_538), .C(n_517), .D(n_513), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_566), .A2(n_538), .B1(n_513), .B2(n_545), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
OAI211xp5_ASAP7_75t_SL g631 ( .A1(n_561), .A2(n_545), .B(n_283), .C(n_280), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_592), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_574), .A2(n_236), .B1(n_276), .B2(n_283), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_550), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_555), .A2(n_276), .B(n_209), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_555), .B(n_219), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_567), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_577), .A2(n_182), .B1(n_184), .B2(n_219), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
NAND4xp25_ASAP7_75t_L g640 ( .A(n_569), .B(n_182), .C(n_184), .D(n_590), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_556), .B(n_184), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_586), .B(n_568), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_591), .B(n_593), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_557), .B(n_592), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_589), .A2(n_569), .B(n_581), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
AOI22x1_ASAP7_75t_L g647 ( .A1(n_585), .A2(n_584), .B1(n_595), .B2(n_562), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_561), .A2(n_296), .B1(n_551), .B2(n_553), .C(n_228), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_602), .A2(n_645), .B1(n_628), .B2(n_616), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_597), .A2(n_617), .B(n_632), .Y(n_650) );
XNOR2xp5_ASAP7_75t_L g651 ( .A(n_601), .B(n_647), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_611), .B(n_605), .Y(n_652) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_632), .Y(n_653) );
OAI21xp33_ASAP7_75t_SL g654 ( .A1(n_597), .A2(n_643), .B(n_604), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g655 ( .A1(n_612), .A2(n_600), .B(n_648), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_SL g656 ( .A1(n_638), .A2(n_643), .B(n_641), .C(n_618), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_596), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
AOI22x1_ASAP7_75t_L g659 ( .A1(n_608), .A2(n_607), .B1(n_627), .B2(n_598), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_640), .B(n_631), .C(n_603), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_607), .A2(n_614), .B1(n_629), .B2(n_634), .Y(n_661) );
NAND4xp75_ASAP7_75t_L g662 ( .A(n_654), .B(n_636), .C(n_608), .D(n_642), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_652), .B(n_635), .C(n_633), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_658), .B(n_609), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_650), .A2(n_644), .B(n_623), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_660), .B(n_607), .C(n_626), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_649), .A2(n_625), .B(n_639), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_659), .A2(n_646), .B1(n_637), .B2(n_624), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_655), .A2(n_621), .B1(n_630), .B2(n_599), .C(n_610), .Y(n_669) );
OAI311xp33_ASAP7_75t_L g670 ( .A1(n_667), .A2(n_656), .A3(n_651), .B1(n_657), .C1(n_661), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_664), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_663), .A2(n_653), .B1(n_620), .B2(n_624), .Y(n_672) );
NAND3xp33_ASAP7_75t_SL g673 ( .A(n_668), .B(n_653), .C(n_623), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g674 ( .A1(n_671), .A2(n_666), .B(n_669), .C(n_664), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g675 ( .A1(n_670), .A2(n_665), .B(n_662), .C(n_622), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_673), .A2(n_620), .B1(n_610), .B2(n_599), .Y(n_676) );
XNOR2xp5_ASAP7_75t_L g677 ( .A(n_676), .B(n_672), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_675), .B(n_619), .C(n_615), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_678), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g680 ( .A(n_679), .B(n_677), .Y(n_680) );
XNOR2xp5_ASAP7_75t_L g681 ( .A(n_680), .B(n_674), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_606), .B(n_613), .Y(n_682) );
endmodule