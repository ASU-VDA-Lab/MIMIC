module fake_jpeg_14915_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_3),
.B(n_0),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_18),
.B(n_21),
.Y(n_23)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_19),
.B(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_11),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_25),
.C(n_26),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_10),
.C(n_9),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_12),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g28 ( 
.A1(n_19),
.A2(n_6),
.A3(n_17),
.B1(n_15),
.B2(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_1),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_26),
.B1(n_16),
.B2(n_24),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_8),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_8),
.C(n_6),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_31),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_1),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.C(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_35),
.B2(n_37),
.Y(n_45)
);


endmodule