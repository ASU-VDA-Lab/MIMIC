module fake_aes_12137_n_486 (n_117, n_44, n_133, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_139, n_16, n_13, n_113, n_95, n_124, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_136, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_134, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_132, n_51, n_96, n_39, n_486);
input n_117;
input n_44;
input n_133;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_139;
input n_16;
input n_13;
input n_113;
input n_95;
input n_124;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_51;
input n_96;
input n_39;
output n_486;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_479;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_475;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_5), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_47), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g143 ( .A(n_12), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_68), .Y(n_144) );
INVx2_ASAP7_75t_SL g145 ( .A(n_89), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_100), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_52), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_124), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_24), .Y(n_149) );
INVxp67_ASAP7_75t_SL g150 ( .A(n_122), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_50), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_66), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_3), .Y(n_154) );
BUFx10_ASAP7_75t_L g155 ( .A(n_51), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_106), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_19), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_49), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_43), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
INVx4_ASAP7_75t_R g161 ( .A(n_128), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_67), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_94), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_20), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_86), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_28), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_71), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_31), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_115), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_53), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_30), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_48), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_81), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_69), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_54), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_60), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
INVxp67_ASAP7_75t_L g179 ( .A(n_80), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_64), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_105), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_85), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_39), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_127), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_117), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_73), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_93), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_91), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_103), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_9), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_116), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_6), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_82), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_18), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_102), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_10), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_15), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_61), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_57), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_76), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_45), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_101), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_65), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_139), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_131), .Y(n_209) );
BUFx5_ASAP7_75t_L g210 ( .A(n_113), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_210), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_210), .Y(n_212) );
INVx6_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_153), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_174), .B(n_0), .Y(n_215) );
INVx5_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_142), .A2(n_21), .B(n_17), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_193), .B(n_1), .Y(n_218) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_148), .A2(n_23), .B(n_22), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_143), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_195), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_154), .Y(n_224) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_172), .A2(n_26), .B(n_25), .Y(n_225) );
INVx6_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_210), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_151), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_145), .B(n_2), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_157), .Y(n_230) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_144), .A2(n_29), .B(n_27), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_229), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx6_ASAP7_75t_L g234 ( .A(n_229), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_213), .Y(n_236) );
INVx5_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
INVx3_ASAP7_75t_L g238 ( .A(n_229), .Y(n_238) );
INVx4_ASAP7_75t_L g239 ( .A(n_215), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_228), .B(n_140), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_212), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_213), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_212), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_227), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_227), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_228), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_230), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_214), .Y(n_252) );
OR2x6_ASAP7_75t_L g253 ( .A(n_218), .B(n_200), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_220), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_234), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_235), .Y(n_257) );
CKINVDCx11_ASAP7_75t_R g258 ( .A(n_253), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_234), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_235), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_250), .A2(n_225), .B(n_217), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_239), .B(n_223), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_239), .B(n_149), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_253), .B(n_213), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_238), .B(n_156), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_238), .B(n_160), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_242), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_232), .B(n_241), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_232), .B(n_226), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_247), .B(n_226), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_247), .B(n_230), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_249), .B(n_224), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
NOR2xp33_ASAP7_75t_SL g274 ( .A(n_252), .B(n_147), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_234), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_251), .B(n_162), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_233), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_236), .B(n_201), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_242), .Y(n_279) );
NOR2xp33_ASAP7_75t_SL g280 ( .A(n_251), .B(n_159), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_243), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_243), .B(n_222), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_257), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_273), .A2(n_245), .B(n_246), .C(n_244), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_246), .B(n_244), .C(n_152), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_264), .A2(n_179), .B(n_182), .C(n_150), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
AO31x2_ASAP7_75t_L g288 ( .A1(n_277), .A2(n_260), .A3(n_267), .B(n_257), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_280), .B(n_141), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_258), .Y(n_290) );
O2A1O1Ixp5_ASAP7_75t_L g291 ( .A1(n_261), .A2(n_194), .B(n_208), .C(n_196), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_278), .B(n_146), .Y(n_292) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_265), .A2(n_163), .B(n_168), .C(n_167), .Y(n_293) );
AO32x1_ASAP7_75t_L g294 ( .A1(n_281), .A2(n_189), .A3(n_169), .B1(n_170), .B2(n_177), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_276), .A2(n_231), .B(n_217), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_263), .A2(n_231), .B(n_217), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_263), .A2(n_231), .B(n_175), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_265), .A2(n_181), .B(n_180), .Y(n_299) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_282), .B(n_2), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_258), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_268), .A2(n_184), .B1(n_186), .B2(n_183), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_188), .B(n_191), .C(n_187), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_274), .A2(n_266), .B1(n_259), .B2(n_256), .Y(n_306) );
AND2x6_ASAP7_75t_L g307 ( .A(n_270), .B(n_197), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_267), .A2(n_203), .B(n_198), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_295), .A2(n_279), .B(n_271), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_296), .A2(n_209), .B(n_207), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_302), .Y(n_311) );
BUFx8_ASAP7_75t_L g312 ( .A(n_290), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_287), .B(n_275), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_308), .A2(n_254), .B(n_248), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_298), .A2(n_255), .B(n_254), .Y(n_316) );
AOI21x1_ASAP7_75t_L g317 ( .A1(n_300), .A2(n_299), .B(n_305), .Y(n_317) );
AOI21xp5_ASAP7_75t_SL g318 ( .A1(n_285), .A2(n_176), .B(n_178), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_291), .A2(n_255), .B(n_210), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_297), .A2(n_210), .B(n_185), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g322 ( .A1(n_284), .A2(n_165), .B(n_164), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_293), .A2(n_210), .B(n_185), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_288), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_292), .A2(n_171), .B(n_166), .Y(n_325) );
OAI21x1_ASAP7_75t_L g326 ( .A1(n_304), .A2(n_185), .B(n_178), .Y(n_326) );
AOI21x1_ASAP7_75t_L g327 ( .A1(n_289), .A2(n_161), .B(n_178), .Y(n_327) );
AO31x2_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_220), .A3(n_221), .B(n_190), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_286), .B(n_173), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_306), .Y(n_330) );
AO21x1_ASAP7_75t_L g331 ( .A1(n_294), .A2(n_221), .B(n_33), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_307), .A2(n_199), .B1(n_192), .B2(n_206), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_288), .B(n_4), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_309), .A2(n_216), .B(n_34), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_332), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_330), .A2(n_202), .B1(n_205), .B2(n_204), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_324), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_316), .A2(n_35), .B(n_32), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_310), .A2(n_37), .B(n_36), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_334), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_312), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_321), .A2(n_40), .B(n_38), .Y(n_345) );
BUFx12f_ASAP7_75t_L g346 ( .A(n_314), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_315), .A2(n_42), .B(n_41), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_320), .A2(n_240), .B(n_237), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_331), .A2(n_46), .B(n_44), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_323), .A2(n_92), .B(n_138), .Y(n_351) );
AO21x2_ASAP7_75t_L g352 ( .A1(n_317), .A2(n_90), .B(n_137), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVx4_ASAP7_75t_SL g354 ( .A(n_328), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_326), .A2(n_88), .B(n_134), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_327), .A2(n_87), .B(n_133), .Y(n_356) );
NOR2x1_ASAP7_75t_SL g357 ( .A(n_335), .B(n_7), .Y(n_357) );
NOR2xp33_ASAP7_75t_SL g358 ( .A(n_322), .B(n_8), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_333), .B(n_11), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_318), .A2(n_97), .B(n_130), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_325), .B(n_13), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_328), .A2(n_98), .B(n_129), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
AO21x1_ASAP7_75t_L g365 ( .A1(n_329), .A2(n_14), .B(n_16), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_364), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_342), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_358), .Y(n_372) );
OAI21x1_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_55), .B(n_56), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_340), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_353), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_340), .B(n_58), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_339), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_359), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_343), .A2(n_62), .B(n_63), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_344), .B(n_72), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_362), .B(n_74), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_357), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_349), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
OA21x2_ASAP7_75t_L g390 ( .A1(n_347), .A2(n_75), .B(n_77), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
AO21x2_ASAP7_75t_L g392 ( .A1(n_352), .A2(n_78), .B(n_79), .Y(n_392) );
BUFx2_ASAP7_75t_L g393 ( .A(n_361), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_352), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_348), .A2(n_83), .B(n_84), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_360), .B(n_99), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_393), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_398), .B(n_104), .Y(n_404) );
OAI321xp33_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_107), .A3(n_108), .B1(n_109), .B2(n_111), .C(n_112), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_386), .B(n_114), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_396), .B(n_375), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_391), .A2(n_125), .B(n_118), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_369), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_367), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_372), .A2(n_119), .B1(n_120), .B2(n_121), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_387), .B(n_123), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_377), .B(n_384), .Y(n_419) );
BUFx3_ASAP7_75t_L g420 ( .A(n_402), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_369), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_381), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_380), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_373), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_373), .Y(n_431) );
INVx2_ASAP7_75t_R g432 ( .A(n_400), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_394), .B(n_401), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_388), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_388), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_382), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_409), .B(n_403), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_403), .B(n_416), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_407), .B(n_370), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_371), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_410), .B(n_382), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_415), .B(n_395), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_433), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_368), .Y(n_448) );
BUFx2_ASAP7_75t_SL g449 ( .A(n_420), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_388), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_421), .B(n_423), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_424), .B(n_419), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_425), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_425), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_437), .B(n_439), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_438), .B(n_440), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_436), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_427), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_441), .B(n_422), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_454), .B(n_432), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_442), .B(n_432), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g465 ( .A(n_459), .B(n_408), .Y(n_465) );
OR2x6_ASAP7_75t_L g466 ( .A(n_449), .B(n_430), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_447), .B(n_426), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_467), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_466), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_462), .B(n_452), .Y(n_471) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_470), .A2(n_466), .B(n_465), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_469), .Y(n_473) );
OAI211xp5_ASAP7_75t_L g474 ( .A1(n_472), .A2(n_464), .B(n_463), .C(n_471), .Y(n_474) );
NAND3xp33_ASAP7_75t_SL g475 ( .A(n_474), .B(n_414), .C(n_473), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g476 ( .A(n_475), .B(n_405), .C(n_411), .D(n_417), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_476), .B(n_468), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_477), .B(n_460), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_478), .Y(n_479) );
AOI22x1_ASAP7_75t_L g480 ( .A1(n_479), .A2(n_434), .B1(n_412), .B2(n_431), .Y(n_480) );
AOI22xp5_ASAP7_75t_SL g481 ( .A1(n_480), .A2(n_428), .B1(n_429), .B2(n_412), .Y(n_481) );
OAI222xp33_ASAP7_75t_L g482 ( .A1(n_481), .A2(n_443), .B1(n_435), .B2(n_450), .C1(n_444), .C2(n_445), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_482), .A2(n_457), .B1(n_412), .B2(n_458), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_483), .A2(n_458), .B1(n_446), .B2(n_448), .Y(n_484) );
AND2x2_ASAP7_75t_SL g485 ( .A(n_484), .B(n_456), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_485), .A2(n_451), .B1(n_453), .B2(n_455), .Y(n_486) );
endmodule