module real_aes_9033_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g234 ( .A1(n_0), .A2(n_235), .B(n_238), .C(n_242), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_1), .B(n_226), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_2), .B(n_236), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g152 ( .A1(n_3), .A2(n_40), .B1(n_153), .B2(n_155), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_4), .A2(n_9), .B1(n_166), .B2(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g167 ( .A(n_4), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_4), .A2(n_196), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_5), .A2(n_228), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g183 ( .A(n_6), .Y(n_183) );
AND2x6_ASAP7_75t_L g201 ( .A(n_6), .B(n_181), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_6), .B(n_507), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_7), .A2(n_201), .B(n_203), .C(n_292), .Y(n_291) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_8), .A2(n_21), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g166 ( .A(n_9), .Y(n_166) );
INVx1_ASAP7_75t_L g221 ( .A(n_10), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_11), .B(n_236), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_12), .Y(n_100) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_13), .A2(n_23), .B1(n_90), .B2(n_94), .Y(n_93) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_14), .A2(n_203), .B(n_206), .C(n_214), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_15), .B(n_113), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_16), .A2(n_203), .B(n_214), .C(n_306), .Y(n_305) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_17), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g101 ( .A1(n_18), .A2(n_34), .B1(n_102), .B2(n_107), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_19), .A2(n_196), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g199 ( .A(n_20), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_22), .A2(n_254), .B(n_255), .C(n_259), .Y(n_253) );
OAI221xp5_ASAP7_75t_L g174 ( .A1(n_23), .A2(n_37), .B1(n_51), .B2(n_175), .C(n_176), .Y(n_174) );
INVxp67_ASAP7_75t_L g177 ( .A(n_23), .Y(n_177) );
AOI22xp33_ASAP7_75t_SL g134 ( .A1(n_24), .A2(n_56), .B1(n_135), .B2(n_138), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_25), .B(n_308), .Y(n_307) );
AOI22xp33_ASAP7_75t_SL g157 ( .A1(n_26), .A2(n_47), .B1(n_158), .B2(n_160), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_27), .B(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g299 ( .A(n_28), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_29), .B(n_236), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_30), .B(n_196), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_31), .A2(n_254), .B(n_259), .C(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g239 ( .A(n_32), .Y(n_239) );
INVx1_ASAP7_75t_L g282 ( .A(n_33), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_35), .B(n_196), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_36), .Y(n_223) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_37), .A2(n_63), .B1(n_90), .B2(n_94), .Y(n_97) );
INVxp67_ASAP7_75t_L g178 ( .A(n_37), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_38), .A2(n_82), .B1(n_83), .B2(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_38), .Y(n_514) );
INVx1_ASAP7_75t_L g181 ( .A(n_39), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_41), .B(n_196), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_42), .B(n_226), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_43), .A2(n_213), .B(n_269), .C(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g220 ( .A(n_44), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_45), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_46), .B(n_236), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_48), .B(n_237), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g142 ( .A1(n_49), .A2(n_59), .B1(n_143), .B2(n_147), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_50), .B(n_121), .Y(n_120) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_68), .B1(n_90), .B2(n_91), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_52), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_53), .B(n_208), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_54), .A2(n_203), .B(n_259), .C(n_322), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g267 ( .A(n_55), .Y(n_267) );
AOI22xp33_ASAP7_75t_SL g124 ( .A1(n_57), .A2(n_75), .B1(n_125), .B2(n_129), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_58), .B(n_211), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_60), .A2(n_163), .B1(n_169), .B2(n_170), .Y(n_162) );
INVx1_ASAP7_75t_L g169 ( .A(n_60), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_61), .Y(n_261) );
INVx1_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
INVx2_ASAP7_75t_L g218 ( .A(n_64), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_65), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_66), .B(n_241), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_67), .B(n_196), .Y(n_252) );
INVx1_ASAP7_75t_L g256 ( .A(n_69), .Y(n_256) );
INVxp67_ASAP7_75t_L g272 ( .A(n_70), .Y(n_272) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_72), .A2(n_164), .B1(n_165), .B2(n_168), .Y(n_163) );
INVx1_ASAP7_75t_L g168 ( .A(n_72), .Y(n_168) );
INVx1_ASAP7_75t_L g289 ( .A(n_73), .Y(n_289) );
AOI22xp5_ASAP7_75t_SL g503 ( .A1(n_73), .A2(n_82), .B1(n_83), .B2(n_289), .Y(n_503) );
INVx1_ASAP7_75t_L g323 ( .A(n_74), .Y(n_323) );
AND2x2_ASAP7_75t_L g284 ( .A(n_76), .B(n_217), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_171), .B1(n_184), .B2(n_499), .C(n_502), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_162), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND2x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_132), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_111), .Y(n_84) );
OAI21xp5_ASAP7_75t_SL g85 ( .A1(n_86), .A2(n_100), .B(n_101), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x6_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x4_ASAP7_75t_L g108 ( .A(n_88), .B(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_93), .Y(n_88) );
AND2x2_ASAP7_75t_L g106 ( .A(n_89), .B(n_97), .Y(n_106) );
INVx2_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
OR2x2_ASAP7_75t_L g118 ( .A(n_93), .B(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g123 ( .A(n_93), .B(n_119), .Y(n_123) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
AND2x6_ASAP7_75t_L g137 ( .A(n_95), .B(n_117), .Y(n_137) );
AND2x2_ASAP7_75t_L g154 ( .A(n_95), .B(n_146), .Y(n_154) );
AND2x4_ASAP7_75t_L g159 ( .A(n_95), .B(n_123), .Y(n_159) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g116 ( .A(n_96), .B(n_99), .Y(n_116) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g141 ( .A(n_97), .B(n_110), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_97), .B(n_99), .Y(n_150) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_99), .Y(n_110) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g127 ( .A(n_105), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g126 ( .A(n_106), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g129 ( .A(n_106), .B(n_130), .Y(n_129) );
BUFx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_120), .C(n_124), .Y(n_111) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx4_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x6_ASAP7_75t_L g122 ( .A(n_116), .B(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g145 ( .A(n_116), .B(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g146 ( .A(n_119), .B(n_128), .Y(n_146) );
BUFx4f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g140 ( .A(n_123), .B(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g148 ( .A(n_128), .Y(n_148) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_151), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_142), .Y(n_133) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx11_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx8_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g156 ( .A(n_141), .B(n_146), .Y(n_156) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g161 ( .A(n_146), .B(n_149), .Y(n_161) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_157), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_163), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
AND3x1_ASAP7_75t_SL g173 ( .A(n_174), .B(n_179), .C(n_182), .Y(n_173) );
INVxp67_ASAP7_75t_L g507 ( .A(n_174), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_179), .A2(n_197), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_179), .Y(n_518) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_180), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_180), .B(n_183), .Y(n_512) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OR2x2_ASAP7_75t_SL g517 ( .A(n_182), .B(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_188), .B(n_435), .Y(n_187) );
NOR5xp2_ASAP7_75t_L g188 ( .A(n_189), .B(n_366), .C(n_395), .D(n_415), .E(n_422), .Y(n_188) );
OAI211xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_246), .B(n_310), .C(n_353), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_191), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_437) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_225), .Y(n_191) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_192), .Y(n_313) );
AND2x4_ASAP7_75t_L g346 ( .A(n_192), .B(n_347), .Y(n_346) );
INVx5_ASAP7_75t_L g364 ( .A(n_192), .Y(n_364) );
AND2x2_ASAP7_75t_L g373 ( .A(n_192), .B(n_365), .Y(n_373) );
AND2x2_ASAP7_75t_L g385 ( .A(n_192), .B(n_250), .Y(n_385) );
AND2x2_ASAP7_75t_L g481 ( .A(n_192), .B(n_349), .Y(n_481) );
OR2x6_ASAP7_75t_L g192 ( .A(n_193), .B(n_222), .Y(n_192) );
AOI21xp5_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_202), .B(n_215), .Y(n_193) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_195), .Y(n_501) );
BUFx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_201), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_197), .B(n_201), .Y(n_290) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
INVx1_ASAP7_75t_L g213 ( .A(n_198), .Y(n_213) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g204 ( .A(n_199), .Y(n_204) );
INVx1_ASAP7_75t_L g297 ( .A(n_199), .Y(n_297) );
INVx1_ASAP7_75t_L g205 ( .A(n_200), .Y(n_205) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_200), .Y(n_209) );
INVx3_ASAP7_75t_L g237 ( .A(n_200), .Y(n_237) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_200), .Y(n_241) );
INVx1_ASAP7_75t_L g308 ( .A(n_200), .Y(n_308) );
BUFx3_ASAP7_75t_L g214 ( .A(n_201), .Y(n_214) );
INVx4_ASAP7_75t_SL g244 ( .A(n_201), .Y(n_244) );
INVx5_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
AND2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
BUFx3_ASAP7_75t_L g243 ( .A(n_204), .Y(n_243) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_204), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_210), .B(n_212), .Y(n_206) );
INVx2_ASAP7_75t_L g211 ( .A(n_208), .Y(n_211) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx4_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_211), .A2(n_256), .B(n_257), .C(n_258), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_211), .A2(n_258), .B(n_282), .C(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g224 ( .A(n_217), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_217), .A2(n_252), .B(n_253), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_217), .A2(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x2_ASAP7_75t_L g229 ( .A(n_218), .B(n_219), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g347 ( .A(n_225), .Y(n_347) );
AND2x2_ASAP7_75t_L g365 ( .A(n_225), .B(n_319), .Y(n_365) );
AND2x2_ASAP7_75t_L g384 ( .A(n_225), .B(n_318), .Y(n_384) );
AND2x2_ASAP7_75t_L g424 ( .A(n_225), .B(n_364), .Y(n_424) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_230), .B(n_245), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_227), .A2(n_288), .B(n_298), .Y(n_287) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_227), .A2(n_320), .B(n_328), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_227), .B(n_329), .Y(n_328) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_228), .A2(n_304), .B(n_305), .Y(n_303) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g300 ( .A(n_229), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_232), .A2(n_233), .B(n_234), .C(n_244), .Y(n_231) );
INVx2_ASAP7_75t_L g254 ( .A(n_233), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g266 ( .A1(n_233), .A2(n_244), .B(n_267), .C(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_236), .B(n_272), .Y(n_271) );
INVx5_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx4_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_243), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_244), .Y(n_259) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_274), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI322xp5_ASAP7_75t_L g483 ( .A1(n_249), .A2(n_285), .A3(n_338), .B1(n_346), .B2(n_400), .C1(n_484), .C2(n_487), .Y(n_483) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_262), .Y(n_249) );
INVx5_ASAP7_75t_L g315 ( .A(n_250), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_250), .B(n_317), .Y(n_332) );
BUFx2_ASAP7_75t_L g410 ( .A(n_250), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_250), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g487 ( .A(n_250), .B(n_394), .Y(n_487) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_260), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_262), .B(n_276), .Y(n_341) );
INVx1_ASAP7_75t_L g368 ( .A(n_262), .Y(n_368) );
AND2x2_ASAP7_75t_L g381 ( .A(n_262), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g482 ( .A(n_262), .B(n_400), .Y(n_482) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g336 ( .A(n_263), .B(n_276), .Y(n_336) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_263), .Y(n_344) );
OR2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g361 ( .A(n_263), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_263), .B(n_287), .Y(n_390) );
INVxp67_ASAP7_75t_L g414 ( .A(n_263), .Y(n_414) );
AND2x2_ASAP7_75t_L g421 ( .A(n_263), .B(n_285), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_263), .B(n_301), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_263), .B(n_286), .Y(n_447) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_273), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_269), .A2(n_323), .B(n_324), .C(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_285), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_276), .B(n_302), .Y(n_391) );
OR2x2_ASAP7_75t_L g413 ( .A(n_276), .B(n_286), .Y(n_413) );
AND2x2_ASAP7_75t_L g426 ( .A(n_276), .B(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_276), .B(n_381), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_276), .A2(n_437), .B(n_442), .C(n_451), .Y(n_436) );
AND2x2_ASAP7_75t_L g497 ( .A(n_276), .B(n_301), .Y(n_497) );
INVx5_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g350 ( .A(n_277), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_277), .B(n_345), .Y(n_357) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_277), .Y(n_359) );
OR2x2_ASAP7_75t_L g370 ( .A(n_277), .B(n_286), .Y(n_370) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_277), .B(n_361), .Y(n_375) );
AND2x2_ASAP7_75t_L g400 ( .A(n_277), .B(n_286), .Y(n_400) );
AND2x2_ASAP7_75t_L g420 ( .A(n_277), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g458 ( .A(n_277), .B(n_285), .Y(n_458) );
OR2x2_ASAP7_75t_L g461 ( .A(n_277), .B(n_447), .Y(n_461) );
OR2x6_ASAP7_75t_L g277 ( .A(n_278), .B(n_284), .Y(n_277) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_301), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_286), .A2(n_405), .B(n_408), .C(n_414), .Y(n_404) );
INVx5_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_287), .B(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g339 ( .A(n_287), .B(n_302), .Y(n_339) );
OR2x2_ASAP7_75t_L g345 ( .A(n_287), .B(n_301), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_291), .Y(n_288) );
OAI322xp33_ASAP7_75t_L g502 ( .A1(n_289), .A2(n_503), .A3(n_504), .B1(n_508), .B2(n_509), .C1(n_513), .C2(n_515), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_295), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_295), .A2(n_307), .B(n_309), .Y(n_306) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_SL g362 ( .A(n_301), .Y(n_362) );
OR2x2_ASAP7_75t_L g490 ( .A(n_301), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_330), .B(n_333), .C(n_342), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI31xp33_ASAP7_75t_L g415 ( .A1(n_312), .A2(n_416), .A3(n_418), .B(n_419), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_313), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_314), .B(n_346), .Y(n_352) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_315), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g372 ( .A(n_315), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g377 ( .A(n_315), .B(n_347), .Y(n_377) );
AND2x2_ASAP7_75t_L g387 ( .A(n_315), .B(n_346), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_315), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g407 ( .A(n_315), .B(n_364), .Y(n_407) );
AND2x2_ASAP7_75t_L g412 ( .A(n_315), .B(n_384), .Y(n_412) );
OR2x2_ASAP7_75t_L g431 ( .A(n_315), .B(n_317), .Y(n_431) );
OR2x2_ASAP7_75t_L g433 ( .A(n_315), .B(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_315), .Y(n_480) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g380 ( .A(n_317), .B(n_347), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_317), .B(n_364), .Y(n_403) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_327), .Y(n_320) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g440 ( .A(n_332), .B(n_364), .Y(n_440) );
AOI322xp5_ASAP7_75t_L g442 ( .A1(n_332), .A2(n_346), .A3(n_384), .B1(n_443), .B2(n_444), .C1(n_445), .C2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g450 ( .A(n_332), .Y(n_450) );
NAND2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
INVx1_ASAP7_75t_SL g444 ( .A(n_334), .Y(n_444) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
OR2x2_ASAP7_75t_L g396 ( .A(n_335), .B(n_341), .Y(n_396) );
INVx1_ASAP7_75t_L g427 ( .A(n_335), .Y(n_427) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI32xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .A3(n_348), .B1(n_350), .B2(n_352), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AOI21xp33_ASAP7_75t_SL g382 ( .A1(n_345), .A2(n_360), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g397 ( .A(n_346), .Y(n_397) );
AND2x4_ASAP7_75t_L g394 ( .A(n_347), .B(n_364), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_347), .B(n_430), .Y(n_429) );
AOI322xp5_ASAP7_75t_L g459 ( .A1(n_348), .A2(n_375), .A3(n_394), .B1(n_427), .B2(n_460), .C1(n_462), .C2(n_463), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_348), .A2(n_425), .B1(n_489), .B2(n_490), .C(n_492), .Y(n_488) );
AND2x2_ASAP7_75t_L g376 ( .A(n_349), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g356 ( .A(n_351), .Y(n_356) );
OR2x2_ASAP7_75t_L g428 ( .A(n_351), .B(n_413), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .A3(n_358), .B(n_363), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_387), .B1(n_388), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g399 ( .A(n_356), .B(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_358), .A2(n_399), .B1(n_452), .B2(n_455), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g441 ( .A(n_361), .B(n_410), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_361), .B(n_400), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_362), .B(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g475 ( .A(n_362), .B(n_413), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_363), .A2(n_458), .B1(n_471), .B2(n_474), .Y(n_470) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx2_ASAP7_75t_L g379 ( .A(n_364), .Y(n_379) );
AND2x2_ASAP7_75t_L g462 ( .A(n_364), .B(n_384), .Y(n_462) );
OR2x2_ASAP7_75t_L g464 ( .A(n_364), .B(n_431), .Y(n_464) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_364), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_365), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_365), .B(n_410), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B(n_374), .C(n_386), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_378), .B2(n_381), .C(n_382), .Y(n_374) );
INVxp67_ASAP7_75t_L g486 ( .A(n_377), .Y(n_486) );
INVx1_ASAP7_75t_L g453 ( .A(n_378), .Y(n_453) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
AND2x2_ASAP7_75t_L g417 ( .A(n_379), .B(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_380), .B(n_407), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g449 ( .A(n_384), .Y(n_449) );
AND2x2_ASAP7_75t_L g455 ( .A(n_384), .B(n_410), .Y(n_455) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_SL g443 ( .A(n_391), .Y(n_443) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_394), .B(n_430), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_398), .B2(n_401), .C(n_404), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g491 ( .A(n_400), .Y(n_491) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g409 ( .A(n_403), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_407), .B(n_466), .Y(n_465) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_413), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_411), .A2(n_457), .B(n_459), .C(n_465), .Y(n_456) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g468 ( .A(n_413), .Y(n_468) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI222xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_428), .B2(n_429), .C1(n_432), .C2(n_433), .Y(n_422) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g498 ( .A(n_429), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_430), .B(n_473), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_430), .A2(n_477), .B1(n_479), .B2(n_482), .Y(n_476) );
INVx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
NOR4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_456), .C(n_469), .D(n_488), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_438), .B(n_468), .Y(n_478) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g445 ( .A(n_443), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_446), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .C(n_483), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx2_ASAP7_75t_L g485 ( .A(n_481), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
OAI21xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_495), .B(n_498), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_517), .Y(n_516) );
endmodule