module real_jpeg_16729_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_564),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_1),
.B(n_565),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_103),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_2),
.A2(n_103),
.B1(n_210),
.B2(n_215),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_2),
.A2(n_103),
.B1(n_285),
.B2(n_288),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_3),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g439 ( 
.A(n_4),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_5),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_6),
.A2(n_264),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_6),
.A2(n_264),
.B1(n_457),
.B2(n_459),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_6),
.A2(n_264),
.B1(n_514),
.B2(n_519),
.Y(n_513)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_7),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_7),
.Y(n_404)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_8),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_8),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_8),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_8),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_9),
.A2(n_91),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_91),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_9),
.A2(n_91),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_10),
.A2(n_42),
.B1(n_325),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_10),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_10),
.A2(n_355),
.B1(n_383),
.B2(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_10),
.A2(n_355),
.B1(n_447),
.B2(n_452),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_10),
.A2(n_355),
.B1(n_489),
.B2(n_490),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_12),
.A2(n_320),
.A3(n_324),
.B1(n_326),
.B2(n_331),
.Y(n_319)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_12),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_12),
.A2(n_216),
.B1(n_330),
.B2(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_12),
.B(n_27),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_12),
.B(n_125),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_12),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_12),
.B(n_66),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_12),
.A2(n_99),
.B1(n_330),
.B2(n_522),
.Y(n_521)
);

OAI32xp33_ASAP7_75t_L g525 ( 
.A1(n_12),
.A2(n_526),
.A3(n_528),
.B1(n_529),
.B2(n_533),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_14),
.A2(n_50),
.B1(n_151),
.B2(n_155),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_14),
.A2(n_50),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_14),
.A2(n_50),
.B1(n_338),
.B2(n_344),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_15),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_16),
.A2(n_54),
.B1(n_138),
.B2(n_143),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_16),
.A2(n_54),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_16),
.A2(n_54),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_17),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_232),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_230),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_204),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_22),
.B(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_146),
.C(n_165),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_23),
.A2(n_146),
.B1(n_147),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_64),
.B2(n_145),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_24),
.A2(n_25),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_25),
.B(n_65),
.C(n_95),
.Y(n_229)
);

OAI21x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_41),
.B(n_51),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_26),
.A2(n_41),
.B1(n_56),
.B2(n_209),
.Y(n_208)
);

OAI22x1_ASAP7_75t_SL g298 ( 
.A1(n_26),
.A2(n_56),
.B1(n_261),
.B2(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_26),
.A2(n_56),
.B1(n_354),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_27),
.B(n_52),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_27),
.B(n_199),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_27),
.A2(n_55),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_33),
.Y(n_396)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_36),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_37),
.Y(n_142)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_37),
.Y(n_317)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_44),
.Y(n_333)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_45),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_56),
.A2(n_198),
.B(n_203),
.Y(n_197)
);

OAI21x1_ASAP7_75t_SL g260 ( 
.A1(n_56),
.A2(n_261),
.B(n_266),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_60),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_60),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_60),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_62),
.Y(n_214)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_62),
.Y(n_263)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_63),
.Y(n_335)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_95),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_65),
.A2(n_219),
.B1(n_220),
.B2(n_228),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_65),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_75),
.B(n_85),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_66),
.B(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_66),
.B(n_255),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_66),
.A2(n_75),
.B1(n_444),
.B2(n_446),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_66),
.A2(n_75),
.B1(n_446),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_67),
.B(n_86),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_67),
.A2(n_187),
.B1(n_194),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_67),
.A2(n_194),
.B1(n_512),
.B2(n_513),
.Y(n_511)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_67)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_68),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_68),
.Y(n_252)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_68),
.Y(n_287)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_68),
.Y(n_458)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_68),
.Y(n_496)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_69),
.Y(n_433)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_72),
.Y(n_290)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_72),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_75),
.A2(n_164),
.B(n_549),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_79),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_83),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_84),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_86),
.A2(n_194),
.B(n_195),
.Y(n_373)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI21x1_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_108),
.B(n_135),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_108),
.B1(n_125),
.B2(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_104),
.Y(n_383)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_107),
.Y(n_527)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_108),
.A2(n_137),
.B(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_108),
.A2(n_221),
.B(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_109),
.A2(n_150),
.B1(n_222),
.B2(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_109),
.A2(n_136),
.B(n_223),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_109),
.A2(n_222),
.B1(n_311),
.B2(n_379),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g392 ( 
.A1(n_109),
.A2(n_222),
.B1(n_379),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_109),
.A2(n_222),
.B1(n_393),
.B2(n_521),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_125),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_116),
.B1(n_119),
.B2(n_122),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_116),
.Y(n_312)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_125),
.Y(n_222)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_131),
.Y(n_125)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_127),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_128),
.Y(n_466)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_133),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_147),
.A2(n_148),
.B(n_156),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

INVxp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_164),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_158),
.B(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_163),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_165),
.A2(n_166),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_184),
.B(n_196),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_168),
.B1(n_196),
.B2(n_197),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_167),
.A2(n_168),
.B1(n_186),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_181),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_172),
.Y(n_294)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_173),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_174),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_174),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_174),
.A2(n_456),
.B(n_462),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_174),
.A2(n_330),
.B1(n_487),
.B2(n_488),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_174),
.A2(n_475),
.B1(n_488),
.B2(n_502),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_176),
.Y(n_490)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_177),
.Y(n_461)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_178),
.Y(n_431)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_181),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_194),
.B(n_195),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_193),
.Y(n_453)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_229),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_225),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_274),
.B(n_563),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_270),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_234),
.B(n_270),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_235),
.A2(n_237),
.B1(n_238),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_235),
.Y(n_413)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_239),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_260),
.C(n_267),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g361 ( 
.A(n_240),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_253),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_241),
.B(n_253),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_242),
.Y(n_462)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_245),
.A2(n_337),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_260),
.B(n_268),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_262),
.A2(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_299)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_263),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_415),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_366),
.B(n_407),
.C(n_408),
.D(n_414),
.Y(n_276)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_277),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_357),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_278),
.B(n_357),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_305),
.C(n_307),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_279),
.A2(n_280),
.B1(n_305),
.B2(n_306),
.Y(n_368)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_297),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_298),
.C(n_304),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_295),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g384 ( 
.A(n_282),
.B(n_295),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B(n_291),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_283),
.A2(n_284),
.B1(n_337),
.B2(n_348),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_283),
.A2(n_474),
.B1(n_479),
.B2(n_480),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_283),
.A2(n_291),
.B(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_300),
.A2(n_303),
.B1(n_380),
.B2(n_383),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_300),
.A2(n_303),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_300),
.A2(n_303),
.B1(n_440),
.B2(n_476),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_318),
.C(n_352),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_309),
.B(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_315),
.Y(n_523)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_336),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_319),
.B(n_336),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_330),
.B(n_435),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_SL g444 ( 
.A1(n_330),
.A2(n_434),
.B(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g529 ( 
.A(n_330),
.B(n_530),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_343),
.Y(n_347)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_351),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_358),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_359),
.B(n_361),
.C(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.C(n_385),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_369),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_384),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_384),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.C(n_378),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_378),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_405),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_405),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.C(n_391),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_387),
.B(n_560),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_389),
.A2(n_390),
.B1(n_391),
.B2(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_391),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_397),
.C(n_399),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_392),
.B(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_397),
.A2(n_398),
.B1(n_400),
.B2(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_400),
.Y(n_553)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR3xp33_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_417),
.C(n_420),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_411),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_421),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_556),
.B(n_562),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_543),
.B(n_555),
.Y(n_422)
);

OAI21x1_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_507),
.B(n_542),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_471),
.B(n_506),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_454),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_454),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_442),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_427),
.A2(n_442),
.B1(n_443),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_427),
.Y(n_483)
);

OAI32xp33_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_429),
.A3(n_432),
.B1(n_434),
.B2(n_437),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_463),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_455),
.B(n_464),
.C(n_470),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_470),
.Y(n_463)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_465),
.Y(n_512)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_472),
.A2(n_484),
.B(n_505),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_482),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_482),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_500),
.B(n_504),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_491),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_497),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_501),
.B(n_503),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_508),
.B(n_509),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_524),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_520),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_511),
.B(n_520),
.C(n_524),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_513),
.Y(n_549)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_540),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_525),
.B(n_540),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_537),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_545),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_544),
.B(n_545),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_546),
.A2(n_550),
.B1(n_551),
.B2(n_554),
.Y(n_545)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_546),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_548),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_547),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_548),
.B(n_550),
.C(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_559),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_559),
.Y(n_562)
);


endmodule