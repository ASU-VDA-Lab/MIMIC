module fake_jpeg_28578_n_58 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_24),
.B1(n_25),
.B2(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_3),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_24),
.B1(n_5),
.B2(n_6),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_14),
.B1(n_19),
.B2(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_4),
.Y(n_48)
);

BUFx12f_ASAP7_75t_SL g52 ( 
.A(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_44),
.Y(n_54)
);

OAI321xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_40),
.A3(n_42),
.B1(n_12),
.B2(n_8),
.C(n_16),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_49),
.B1(n_45),
.B2(n_47),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_55),
.C(n_47),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.A3(n_51),
.B1(n_52),
.B2(n_21),
.C(n_4),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_5),
.B(n_7),
.C(n_51),
.Y(n_58)
);


endmodule