module fake_jpeg_29433_n_401 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_401);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_401;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_49),
.B(n_81),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_16),
.A2(n_9),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_50),
.B(n_23),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_9),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_70),
.Y(n_92)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_8),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_77),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_0),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_20),
.B1(n_39),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_86),
.A2(n_96),
.B1(n_38),
.B2(n_52),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_25),
.C(n_20),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_77),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_44),
.A2(n_16),
.B1(n_37),
.B2(n_36),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_0),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_20),
.B1(n_21),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_127),
.B1(n_133),
.B2(n_89),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_27),
.B1(n_39),
.B2(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_26),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_116),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_45),
.B(n_29),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_59),
.B(n_29),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_51),
.B(n_38),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_22),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_55),
.B(n_38),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_42),
.B1(n_32),
.B2(n_24),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_60),
.A2(n_42),
.B1(n_32),
.B2(n_24),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_137),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_138),
.A2(n_161),
.B(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_148),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_125),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_149),
.B1(n_156),
.B2(n_163),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_169),
.B(n_115),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_76),
.B1(n_71),
.B2(n_67),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_119),
.Y(n_151)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_87),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_170),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_99),
.A2(n_38),
.B1(n_52),
.B2(n_4),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_174),
.B1(n_176),
.B2(n_181),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_106),
.B(n_38),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_168),
.C(n_131),
.Y(n_184)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

OR2x2_ASAP7_75t_SL g168 ( 
.A(n_105),
.B(n_92),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_106),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_102),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_3),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_88),
.A2(n_6),
.B1(n_7),
.B2(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_180),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_148),
.Y(n_222)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_6),
.B1(n_7),
.B2(n_111),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_151),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_128),
.B1(n_110),
.B2(n_115),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_144),
.B(n_152),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_186),
.A2(n_214),
.B(n_206),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_118),
.C(n_102),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_187),
.B(n_160),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_179),
.A2(n_150),
.B(n_163),
.C(n_156),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_139),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_93),
.B(n_120),
.C(n_110),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_201),
.A2(n_202),
.B(n_172),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_99),
.B1(n_109),
.B2(n_111),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_219),
.B1(n_145),
.B2(n_178),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_109),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_138),
.A2(n_93),
.B(n_103),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_129),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_129),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_174),
.B1(n_169),
.B2(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_154),
.A2(n_108),
.B1(n_166),
.B2(n_136),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_146),
.B1(n_147),
.B2(n_155),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_166),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_223),
.A2(n_215),
.B(n_210),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_237),
.Y(n_264)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_227),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_228),
.A2(n_238),
.B1(n_242),
.B2(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_246),
.C(n_208),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_141),
.B(n_180),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_236),
.B(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_233),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_224),
.B1(n_218),
.B2(n_225),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_175),
.B(n_177),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_188),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_183),
.A2(n_158),
.B1(n_167),
.B2(n_159),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_257),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_183),
.A2(n_140),
.B1(n_151),
.B2(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_198),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_215),
.B(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_190),
.B(n_191),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_184),
.A2(n_212),
.B1(n_193),
.B2(n_187),
.C(n_221),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_216),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_211),
.Y(n_266)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_255),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_192),
.A2(n_201),
.B1(n_219),
.B2(n_196),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_260),
.A2(n_287),
.B1(n_255),
.B2(n_250),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_285),
.Y(n_303)
);

AO21x2_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_196),
.B(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_224),
.B1(n_236),
.B2(n_244),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_235),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_265),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_233),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_246),
.C(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_270),
.C(n_279),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_204),
.C(n_205),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_271),
.A2(n_275),
.B(n_268),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_237),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_280),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_205),
.C(n_211),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_213),
.C(n_195),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_232),
.A2(n_210),
.B1(n_207),
.B2(n_197),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_271),
.B(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_294),
.B1(n_299),
.B2(n_301),
.Y(n_329)
);

OAI22x1_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_242),
.B1(n_228),
.B2(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_295),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

INVx3_ASAP7_75t_SL g297 ( 
.A(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_251),
.C(n_239),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_306),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_244),
.B1(n_239),
.B2(n_231),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_284),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_305),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_252),
.B1(n_243),
.B2(n_240),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_261),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_245),
.C(n_249),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_308),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_267),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_272),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_310),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_227),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_254),
.Y(n_311)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_318),
.Y(n_341)
);

OAI321xp33_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_294),
.A3(n_266),
.B1(n_296),
.B2(n_302),
.C(n_268),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_269),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_328),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_262),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_326),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_285),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_270),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_279),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_292),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_282),
.C(n_277),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_287),
.C(n_263),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_329),
.A2(n_304),
.B1(n_306),
.B2(n_263),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_338),
.A2(n_322),
.B1(n_319),
.B2(n_317),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_327),
.A2(n_309),
.B1(n_312),
.B2(n_308),
.Y(n_340)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_305),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_347),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_291),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_344),
.B(n_345),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_263),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_349),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_315),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_352),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_295),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_353),
.C(n_326),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_247),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_288),
.C(n_281),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_341),
.A2(n_333),
.B(n_318),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_344),
.B(n_349),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_364),
.C(n_366),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_345),
.B(n_329),
.CI(n_323),
.CON(n_357),
.SN(n_357)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_358),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_348),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_297),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_331),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_361),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_276),
.C(n_288),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_276),
.C(n_281),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_300),
.C(n_272),
.Y(n_367)
);

AOI31xp33_ASAP7_75t_L g374 ( 
.A1(n_367),
.A2(n_207),
.A3(n_197),
.B(n_198),
.Y(n_374)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_368),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_361),
.A2(n_339),
.B1(n_338),
.B2(n_353),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_375),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_370),
.A2(n_374),
.B(n_377),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_SL g373 ( 
.A1(n_357),
.A2(n_297),
.B(n_351),
.C(n_336),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_336),
.Y(n_375)
);

HAxp5_ASAP7_75t_SL g376 ( 
.A(n_354),
.B(n_365),
.CON(n_376),
.SN(n_376)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_355),
.C(n_362),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_SL g377 ( 
.A(n_362),
.B(n_363),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_381),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_356),
.C(n_364),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_357),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_385),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_366),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_386),
.B(n_355),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_388),
.A2(n_373),
.B(n_383),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_390),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_376),
.B(n_372),
.Y(n_391)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_373),
.B(n_392),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_386),
.C(n_384),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_373),
.C(n_388),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_394),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_395),
.B(n_396),
.CI(n_397),
.CON(n_398),
.SN(n_398)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_389),
.C(n_399),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_398),
.Y(n_401)
);


endmodule