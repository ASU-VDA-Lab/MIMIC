module fake_aes_2155_n_19 (n_1, n_2, n_0, n_19);
input n_1;
input n_2;
input n_0;
output n_19;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_3;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_6;
wire n_4;
wire n_7;
AND2x4_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
BUFx6f_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_SL g5 ( .A(n_1), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
OAI22xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_7) );
OAI21x1_ASAP7_75t_L g8 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_10), .B(n_6), .Y(n_11) );
BUFx2_ASAP7_75t_SL g12 ( .A(n_9), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_3), .B1(n_5), .B2(n_4), .C(n_9), .Y(n_13) );
O2A1O1Ixp33_ASAP7_75t_L g14 ( .A1(n_12), .A2(n_3), .B(n_4), .C(n_10), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_14), .B(n_3), .Y(n_15) );
NOR3x2_ASAP7_75t_L g16 ( .A(n_13), .B(n_3), .C(n_4), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_4), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
AOI21x1_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_4), .B(n_18), .Y(n_19) );
endmodule