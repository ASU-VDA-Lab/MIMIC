module fake_jpeg_25809_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_33;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_36),
.B1(n_29),
.B2(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_29),
.B1(n_30),
.B2(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_76)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_57),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_17),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_32),
.B(n_1),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_86),
.B(n_87),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_45),
.B1(n_57),
.B2(n_66),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_79),
.B1(n_19),
.B2(n_31),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_20),
.CON(n_81),
.SN(n_81)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_24),
.C(n_20),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_92),
.B1(n_58),
.B2(n_65),
.Y(n_96)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_43),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_32),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_66),
.B1(n_54),
.B2(n_58),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_99),
.B1(n_92),
.B2(n_82),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_106),
.B1(n_110),
.B2(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_22),
.B1(n_25),
.B2(n_48),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_107),
.Y(n_126)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_20),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_22),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_71),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_63),
.B1(n_56),
.B2(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_26),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_63),
.B1(n_56),
.B2(n_28),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_119),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_28),
.B1(n_33),
.B2(n_27),
.Y(n_113)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_43),
.A3(n_39),
.B1(n_37),
.B2(n_24),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_77),
.C(n_20),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_39),
.C(n_37),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.C(n_86),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_24),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_132),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_136),
.B(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_130),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_125),
.B1(n_131),
.B2(n_141),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_90),
.B1(n_73),
.B2(n_83),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_117),
.A2(n_73),
.B1(n_78),
.B2(n_85),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_128),
.A2(n_88),
.B1(n_31),
.B2(n_69),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_94),
.B1(n_109),
.B2(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_86),
.B1(n_91),
.B2(n_77),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_133),
.A2(n_144),
.B1(n_97),
.B2(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_21),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_80),
.A3(n_86),
.B1(n_19),
.B2(n_16),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_77),
.B(n_1),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_20),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_119),
.B1(n_112),
.B2(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_111),
.B1(n_107),
.B2(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_159),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_112),
.B1(n_108),
.B2(n_16),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_158),
.B1(n_143),
.B2(n_121),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_135),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_118),
.B1(n_108),
.B2(n_78),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_121),
.B1(n_127),
.B2(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_16),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_156),
.B(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_118),
.C(n_74),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_163),
.C(n_169),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_125),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_70),
.B1(n_31),
.B2(n_33),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_164),
.B1(n_141),
.B2(n_69),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_70),
.C(n_55),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_33),
.B1(n_27),
.B2(n_21),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_21),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_161),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_20),
.C(n_21),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_171),
.B1(n_161),
.B2(n_156),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_173),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_120),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_180),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_142),
.B(n_131),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_148),
.B(n_163),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_144),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_153),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_191),
.B1(n_149),
.B2(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_164),
.B1(n_154),
.B2(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_194),
.B1(n_146),
.B2(n_147),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_138),
.B1(n_33),
.B2(n_27),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_188),
.B1(n_190),
.B2(n_176),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_204),
.B(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_202),
.A2(n_209),
.B1(n_210),
.B2(n_191),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_148),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_217),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_157),
.B(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_169),
.B(n_1),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_21),
.B1(n_27),
.B2(n_24),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_24),
.B1(n_69),
.B2(n_3),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_216),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_215),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_14),
.C(n_13),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_214),
.C(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_13),
.C(n_12),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_11),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_221),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_211),
.C(n_184),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_230),
.C(n_206),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_177),
.C(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_180),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_181),
.B(n_172),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_236),
.B(n_199),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_234),
.B1(n_202),
.B2(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_185),
.B1(n_194),
.B2(n_176),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_175),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_175),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_216),
.C(n_203),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_226),
.B(n_214),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_247),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_230),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_235),
.B1(n_219),
.B2(n_225),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_217),
.CI(n_197),
.CON(n_246),
.SN(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_227),
.B1(n_236),
.B2(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_210),
.Y(n_250)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_198),
.C(n_12),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_224),
.C(n_10),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_198),
.B1(n_222),
.B2(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_255),
.B1(n_0),
.B2(n_2),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_0),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_218),
.B1(n_224),
.B2(n_3),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_252),
.B1(n_246),
.B2(n_243),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_10),
.C(n_9),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_251),
.C(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_0),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_0),
.B(n_2),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_237),
.B(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_268),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_271),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_240),
.B1(n_246),
.B2(n_4),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_254),
.C(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_275),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_264),
.B(n_257),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_259),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_258),
.B(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_4),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_271),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_288),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.C(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_7),
.C(n_5),
.Y(n_290)
);

AOI31xp33_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_5),
.A3(n_6),
.B(n_282),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_292),
.B(n_287),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_299),
.B(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_293),
.B(n_298),
.C(n_294),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_297),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_6),
.B(n_302),
.Y(n_304)
);


endmodule