module fake_jpeg_28164_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_67),
.Y(n_68)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_46),
.B1(n_59),
.B2(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_3),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_80),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_54),
.B1(n_59),
.B2(n_44),
.Y(n_74)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_75),
.B1(n_0),
.B2(n_1),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_56),
.B1(n_43),
.B2(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_58),
.B1(n_60),
.B2(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_0),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_1),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_19),
.B(n_38),
.C(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_90),
.Y(n_101)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_14),
.A3(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_12),
.B1(n_31),
.B2(n_30),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_88),
.B(n_91),
.Y(n_103)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_11),
.B1(n_29),
.B2(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_2),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_82),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_100),
.A2(n_81),
.B(n_90),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_113),
.B(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_3),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_98),
.C(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_117),
.C(n_13),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_109),
.A2(n_72),
.B1(n_105),
.B2(n_6),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_21),
.B(n_24),
.Y(n_123)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_115),
.B(n_116),
.C(n_120),
.D(n_121),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_114),
.B1(n_125),
.B2(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_9),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_22),
.B(n_39),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_4),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_130),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_4),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_5),
.Y(n_134)
);


endmodule