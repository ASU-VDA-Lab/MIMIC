module fake_jpeg_1738_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_49),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_10),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_71),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_0),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_63),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_70),
.B1(n_74),
.B2(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_67),
.B1(n_59),
.B2(n_58),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_80),
.A2(n_75),
.B1(n_61),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_98),
.B1(n_68),
.B2(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_1),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_70),
.B1(n_60),
.B2(n_74),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_69),
.B1(n_57),
.B2(n_3),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_75),
.B1(n_61),
.B2(n_76),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_62),
.B1(n_65),
.B2(n_73),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_77),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_55),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_68),
.B1(n_72),
.B2(n_63),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_114),
.Y(n_128)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_101),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_62),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_111),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_91),
.B(n_5),
.Y(n_123)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_1),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_67),
.B1(n_69),
.B2(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_113),
.B1(n_45),
.B2(n_44),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_57),
.B1(n_2),
.B2(n_3),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_8),
.Y(n_136)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_91),
.B1(n_89),
.B2(n_6),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_132),
.B1(n_130),
.B2(n_127),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_101),
.B(n_10),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_134),
.B1(n_109),
.B2(n_110),
.Y(n_152)
);

AO21x2_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_42),
.B(n_41),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_37),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_36),
.C(n_35),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_123),
.C(n_122),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_139),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_32),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_156),
.B(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_162),
.B1(n_16),
.B2(n_17),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_31),
.C(n_30),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_163),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_127),
.B1(n_131),
.B2(n_13),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_11),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_29),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_169),
.B1(n_175),
.B2(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_169)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_162),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_146),
.B(n_149),
.C(n_21),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_23),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_158),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_15),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_143),
.C(n_141),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_159),
.B1(n_161),
.B2(n_163),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_175),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_153),
.B(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_186),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_172),
.B(n_176),
.C(n_181),
.D(n_167),
.Y(n_187)
);

FAx1_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_191),
.CI(n_20),
.CON(n_198),
.SN(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_170),
.C(n_22),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_174),
.A3(n_178),
.B1(n_177),
.B2(n_171),
.C1(n_169),
.C2(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_170),
.Y(n_196)
);

HAxp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_19),
.CON(n_191),
.SN(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_197),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_184),
.C(n_182),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_183),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_23),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_22),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_203),
.A2(n_198),
.B1(n_191),
.B2(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_206),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_194),
.B(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_208),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_209),
.A2(n_205),
.B(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_206),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_187),
.B(n_189),
.C(n_202),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_192),
.Y(n_213)
);


endmodule