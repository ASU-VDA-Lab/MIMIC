module fake_jpeg_6953_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_17),
.B1(n_28),
.B2(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx2_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_51),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_41),
.B1(n_39),
.B2(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_60),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_24),
.B1(n_22),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_18),
.B1(n_20),
.B2(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_37),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_70),
.B1(n_44),
.B2(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_74),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_40),
.B1(n_34),
.B2(n_24),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_71),
.B1(n_19),
.B2(n_17),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_49),
.B(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_22),
.B1(n_56),
.B2(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_58),
.B1(n_57),
.B2(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_22),
.B1(n_59),
.B2(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_69),
.B1(n_76),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_53),
.B1(n_50),
.B2(n_43),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_67),
.C(n_68),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_94),
.Y(n_112)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_58),
.B1(n_57),
.B2(n_42),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_81),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_70),
.B(n_74),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_103),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_75),
.B(n_67),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_72),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_114),
.B1(n_103),
.B2(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_79),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_21),
.B(n_36),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_93),
.B1(n_85),
.B2(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_108),
.C(n_106),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_14),
.B(n_23),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_97),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_143),
.C(n_26),
.Y(n_156)
);

OAI322xp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_98),
.A3(n_99),
.B1(n_92),
.B2(n_105),
.C1(n_48),
.C2(n_61),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_149),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_99),
.B1(n_23),
.B2(n_16),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_130),
.B1(n_124),
.B2(n_131),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_37),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_148),
.B(n_132),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_36),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_119),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_23),
.B(n_16),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_21),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_116),
.B1(n_126),
.B2(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_155),
.B(n_146),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_159),
.B(n_160),
.Y(n_165)
);

OAI22x1_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_120),
.B1(n_121),
.B2(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_158),
.C(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_157),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_42),
.C(n_23),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_16),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_14),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_169),
.B1(n_150),
.B2(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_136),
.B(n_139),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_156),
.B(n_152),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_166),
.B(n_6),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_6),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_152),
.B1(n_141),
.B2(n_2),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_166),
.B(n_165),
.C(n_7),
.D(n_8),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_172),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_174),
.B1(n_176),
.B2(n_173),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_179),
.B1(n_183),
.B2(n_180),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_13),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_185),
.B(n_184),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_181),
.Y(n_188)
);


endmodule