module real_jpeg_4873_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_44),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_44),
.B1(n_94),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_44),
.B1(n_87),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_64),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_2),
.A2(n_64),
.B1(n_145),
.B2(n_379),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_5),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_87),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_6),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_101),
.B1(n_215),
.B2(n_219),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_6),
.A2(n_101),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_6),
.A2(n_101),
.B1(n_288),
.B2(n_290),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_7),
.Y(n_98)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_7),
.Y(n_114)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_9),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_9),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_10),
.A2(n_27),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_10),
.A2(n_27),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_10),
.B(n_92),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_10),
.A2(n_254),
.B(n_255),
.C(n_261),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_10),
.B(n_279),
.C(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_124),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_10),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_10),
.B(n_49),
.Y(n_320)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_359),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_221),
.B(n_357),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_187),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_187),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_15),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_149),
.CI(n_158),
.CON(n_15),
.SN(n_15)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_16),
.B(n_149),
.C(n_158),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_83),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_17),
.B(n_84),
.C(n_117),
.Y(n_386)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_19),
.B(n_47),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_20),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_23),
.A2(n_34),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_23),
.B(n_34),
.Y(n_232)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AO22x1_ASAP7_75t_SL g49 ( 
.A1(n_25),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_26),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_27),
.A2(n_87),
.B(n_89),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_27),
.B(n_90),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_27),
.A2(n_256),
.B(n_258),
.Y(n_255)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_32),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_33),
.A2(n_161),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_34),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_34),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_37),
.Y(n_166)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_40),
.B(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_43),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_58),
.B(n_68),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_48),
.A2(n_155),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_48),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_49),
.B(n_69),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_49),
.B(n_267),
.Y(n_282)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_57),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_58),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_62),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_62),
.Y(n_270)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_68),
.B(n_282),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_68),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_75),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_75),
.B(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_117),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_99),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_86),
.B(n_104),
.Y(n_237)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_86),
.Y(n_374)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_92),
.B(n_100),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_92),
.B(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_92),
.Y(n_373)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_92)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_94),
.Y(n_218)
);

INVx6_ASAP7_75t_L g382 ( 
.A(n_94),
.Y(n_382)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_95),
.Y(n_200)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_95),
.Y(n_208)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_99),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_104),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_104),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_112),
.B2(n_115),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_109),
.B(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_135),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_118),
.B(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_119),
.Y(n_242)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_124),
.A2(n_136),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_124),
.B(n_214),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_124),
.A2(n_241),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_135),
.B(n_243),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_146),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_136),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_137),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_144),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_142),
.Y(n_254)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_149)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_150),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_150),
.A2(n_157),
.B1(n_253),
.B2(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_150),
.B(n_154),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_150),
.A2(n_157),
.B1(n_370),
.B2(n_371),
.Y(n_369)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_156),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_156),
.B(n_266),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_179),
.C(n_181),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_172),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_160),
.B(n_172),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_167),
.B(n_168),
.Y(n_160)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_168),
.B(n_286),
.Y(n_319)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_171),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_173),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_220),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_188),
.B(n_220),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_191),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_209),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_192),
.B(n_209),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_194),
.B(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_197),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.A3(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_341),
.B(n_354),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_271),
.B(n_340),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_248),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_224),
.B(n_248),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_227),
.B(n_233),
.C(n_235),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_232),
.B(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_236),
.B(n_239),
.C(n_245),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_262),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_249),
.B(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_252),
.A2(n_262),
.B1(n_263),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_265),
.B(n_384),
.Y(n_383)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_334),
.B(n_339),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_324),
.B(n_333),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_296),
.B(n_323),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_283),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_283),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_291),
.Y(n_283)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_303),
.Y(n_302)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_294),
.C(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_306),
.B(n_322),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_300),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx8_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_318),
.B(n_321),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_315),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_330),
.C(n_331),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_338),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_350),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_344),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_347),
.C(n_348),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_350),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_353),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_387),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_362),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_386),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_375),
.B2(n_376),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B(n_374),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_383),
.B(n_385),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_377),
.B(n_383),
.Y(n_385)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);


endmodule