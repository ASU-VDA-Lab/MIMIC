module real_jpeg_26386_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

INVx6_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_0),
.Y(n_97)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_29),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_4),
.B(n_33),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_110),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_4),
.B(n_68),
.C(n_82),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_57),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_4),
.A2(n_65),
.B1(n_243),
.B2(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_34),
.B1(n_37),
.B2(n_43),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_6),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_6),
.A2(n_43),
.B1(n_67),
.B2(n_68),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_7),
.A2(n_27),
.B1(n_40),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_7),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_34),
.B1(n_37),
.B2(n_122),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_122),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_7),
.A2(n_67),
.B1(n_68),
.B2(n_122),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_9),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_9),
.A2(n_34),
.B1(n_37),
.B2(n_86),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_11),
.A2(n_34),
.B1(n_37),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_91)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_14),
.A2(n_34),
.B1(n_37),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_51),
.B1(n_67),
.B2(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_51),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_15),
.A2(n_26),
.B1(n_34),
.B2(n_37),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_15),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_15),
.A2(n_26),
.B1(n_67),
.B2(n_68),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_149),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_20),
.B(n_123),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.C(n_105),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_21),
.B(n_92),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_24),
.B(n_47),
.C(n_63),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_42),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_25),
.A2(n_31),
.B1(n_33),
.B2(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_31),
.A2(n_42),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_31),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_32),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_32),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_34),
.A2(n_38),
.B(n_109),
.C(n_111),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_34),
.B(n_110),
.CON(n_193),
.SN(n_193)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_36),
.B(n_37),
.C(n_46),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_37),
.A2(n_56),
.A3(n_59),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_60),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_50),
.B(n_57),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_52),
.A2(n_118),
.B1(n_143),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_52),
.A2(n_143),
.B1(n_160),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_53),
.B(n_61),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_57),
.B1(n_184),
.B2(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AO22x1_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_55),
.B(n_58),
.Y(n_194)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_59),
.B1(n_82),
.B2(n_84),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_59),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_80),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_64),
.B(n_80),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_74),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_65),
.A2(n_131),
.B(n_133),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_65),
.A2(n_74),
.B(n_133),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_65),
.A2(n_95),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_65),
.A2(n_131),
.B1(n_234),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_66),
.B(n_75),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_72),
.B1(n_78),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_66),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_68),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_67),
.B(n_248),
.Y(n_247)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_79),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_85),
.B(n_87),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_91),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_81),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_81),
.B(n_110),
.Y(n_241)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_103),
.B(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_88),
.A2(n_128),
.B(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_88),
.A2(n_102),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_88),
.A2(n_199),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_88),
.A2(n_102),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_88),
.A2(n_102),
.B1(n_198),
.B2(n_219),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_100),
.B2(n_104),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_99),
.A2(n_115),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_105),
.A2(n_106),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.C(n_120),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_110),
.B(n_249),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_148),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_134),
.B1(n_146),
.B2(n_147),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_185),
.B(n_265),
.C(n_270),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_171),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_171),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_168),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_166),
.B2(n_167),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_154),
.B(n_167),
.C(n_168),
.Y(n_266)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_172),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_177),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_204),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_260),
.B(n_264),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_213),
.B(n_259),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_190),
.B(n_200),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_191),
.B(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_195),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_197),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_201),
.B(n_208),
.C(n_212),
.Y(n_261)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_212),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_254),
.B(n_258),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_230),
.B(n_253),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_222),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_216),
.B(n_222),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_220),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_227),
.C(n_228),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_239),
.B(n_252),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_244),
.B(n_251),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_262),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);


endmodule