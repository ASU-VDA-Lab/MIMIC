module fake_aes_9378_n_689 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_689);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_689;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_617;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_69), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_71), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_26), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_28), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_60), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_50), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_9), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_7), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_54), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_35), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_19), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_48), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_37), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_2), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_1), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_20), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_39), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_55), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_65), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_21), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_76), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_22), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_51), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_31), .Y(n_109) );
INVxp33_ASAP7_75t_L g110 ( .A(n_33), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_30), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_23), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_5), .Y(n_114) );
BUFx10_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_24), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_15), .Y(n_117) );
OR2x2_ASAP7_75t_L g118 ( .A(n_47), .B(n_68), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_34), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_17), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_49), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_11), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_64), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_111), .B(n_0), .Y(n_124) );
BUFx8_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_117), .B(n_0), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
CKINVDCx11_ASAP7_75t_R g128 ( .A(n_120), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_117), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_102), .B(n_1), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_84), .B(n_2), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_110), .B(n_3), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_84), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_77), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_87), .B(n_4), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_95), .B(n_7), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_106), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_89), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
BUFx12f_ASAP7_75t_L g146 ( .A(n_115), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_114), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_147) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_88), .B(n_44), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_90), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_122), .B(n_12), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_91), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_120), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_98), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_100), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_103), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_107), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_108), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_113), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_116), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_78), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_79), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_96), .B(n_13), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_152), .B(n_104), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_166), .B(n_104), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
INVx4_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_148), .A2(n_78), .B1(n_119), .B2(n_112), .Y(n_173) );
INVxp33_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_166), .B(n_105), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_141), .A2(n_115), .B1(n_119), .B2(n_105), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
INVxp33_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_152), .B(n_82), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_130), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_164), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_134), .B(n_82), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_146), .B(n_112), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_146), .B(n_101), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_165), .Y(n_188) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
OR2x2_ASAP7_75t_L g190 ( .A(n_131), .B(n_109), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_134), .B(n_109), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_137), .B(n_101), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_137), .B(n_86), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_125), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_141), .A2(n_86), .B1(n_123), .B2(n_97), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_138), .B(n_99), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_130), .B(n_14), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_132), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_151), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_126), .Y(n_206) );
INVx5_ASAP7_75t_L g207 ( .A(n_126), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_126), .B(n_75), .Y(n_208) );
OAI21xp33_ASAP7_75t_SL g209 ( .A1(n_148), .A2(n_16), .B(n_17), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_138), .B(n_16), .Y(n_210) );
BUFx2_ASAP7_75t_L g211 ( .A(n_125), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_126), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_144), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_132), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_127), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_140), .B(n_18), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_140), .B(n_25), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_155), .B(n_27), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_155), .B(n_29), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_160), .B(n_36), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_139), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_179), .B(n_125), .Y(n_226) );
AND2x6_ASAP7_75t_SL g227 ( .A(n_186), .B(n_124), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_216), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_220), .B(n_125), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_170), .B(n_161), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_220), .Y(n_232) );
OR2x6_ASAP7_75t_L g233 ( .A(n_186), .B(n_147), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_179), .B(n_160), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_215), .B(n_161), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_213), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_189), .A2(n_157), .B1(n_159), .B2(n_162), .Y(n_237) );
NAND3xp33_ASAP7_75t_L g238 ( .A(n_176), .B(n_167), .C(n_133), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
BUFx3_ASAP7_75t_L g240 ( .A(n_195), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_190), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_186), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_215), .B(n_163), .Y(n_244) );
INVx8_ASAP7_75t_L g245 ( .A(n_186), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_215), .B(n_163), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_193), .B(n_158), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_178), .B(n_153), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_135), .B(n_143), .C(n_157), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g251 ( .A1(n_173), .A2(n_156), .B1(n_133), .B2(n_129), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_183), .B(n_158), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_189), .A2(n_156), .B1(n_154), .B2(n_142), .Y(n_254) );
NOR2x2_ASAP7_75t_L g255 ( .A(n_174), .B(n_188), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_195), .B(n_154), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_189), .A2(n_159), .B1(n_157), .B2(n_149), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_194), .B(n_149), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_211), .Y(n_259) );
NOR3xp33_ASAP7_75t_L g260 ( .A(n_181), .B(n_142), .C(n_129), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_211), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_175), .B(n_159), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_169), .B(n_150), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_208), .A2(n_150), .B1(n_145), .B2(n_151), .Y(n_264) );
BUFx8_ASAP7_75t_L g265 ( .A(n_201), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_169), .B(n_145), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_187), .B(n_151), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_203), .B(n_145), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_224), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_177), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_169), .B(n_151), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_208), .A2(n_151), .B1(n_41), .B2(n_43), .Y(n_272) );
OAI22xp5_ASAP7_75t_SL g273 ( .A1(n_203), .A2(n_40), .B1(n_45), .B2(n_52), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_172), .B(n_53), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_206), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_208), .Y(n_276) );
NAND3xp33_ASAP7_75t_SL g277 ( .A(n_197), .B(n_56), .C(n_57), .Y(n_277) );
AND2x6_ASAP7_75t_SL g278 ( .A(n_201), .B(n_58), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_168), .B(n_61), .Y(n_279) );
NOR2x1p5_ASAP7_75t_L g280 ( .A(n_190), .B(n_62), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_212), .A2(n_63), .B1(n_67), .B2(n_72), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
AOI22xp33_ASAP7_75t_SL g283 ( .A1(n_187), .A2(n_73), .B1(n_198), .B2(n_208), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_172), .B(n_199), .Y(n_284) );
NOR2x2_ASAP7_75t_L g285 ( .A(n_184), .B(n_208), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_172), .B(n_212), .Y(n_286) );
NOR2xp33_ASAP7_75t_SL g287 ( .A(n_187), .B(n_198), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_212), .B(n_198), .Y(n_288) );
O2A1O1Ixp5_ASAP7_75t_L g289 ( .A1(n_206), .A2(n_219), .B(n_221), .C(n_210), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_246), .Y(n_292) );
BUFx12f_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_249), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_284), .A2(n_206), .B(n_207), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_241), .B(n_207), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_230), .A2(n_221), .B(n_207), .C(n_216), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_230), .B(n_207), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_243), .Y(n_300) );
NOR2xp33_ASAP7_75t_R g301 ( .A(n_245), .B(n_208), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_287), .A2(n_207), .B(n_218), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_289), .A2(n_217), .B(n_180), .Y(n_304) );
INVx5_ASAP7_75t_L g305 ( .A(n_256), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_265), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_232), .A2(n_222), .B1(n_180), .B2(n_182), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_256), .Y(n_308) );
NAND2x1_ASAP7_75t_L g309 ( .A(n_256), .B(n_222), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_276), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_238), .B(n_222), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_234), .B(n_202), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_240), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_259), .B(n_202), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_235), .B(n_182), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_232), .A2(n_205), .B1(n_191), .B2(n_185), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_286), .A2(n_205), .B(n_191), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_260), .B(n_171), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_271), .A2(n_171), .B(n_185), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_254), .B(n_196), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_232), .A2(n_196), .B1(n_214), .B2(n_223), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_233), .B(n_214), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_236), .Y(n_324) );
NOR2xp33_ASAP7_75t_SL g325 ( .A(n_245), .B(n_223), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_276), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_250), .A2(n_225), .B(n_200), .C(n_204), .Y(n_327) );
AOI21x1_ASAP7_75t_L g328 ( .A1(n_267), .A2(n_225), .B(n_200), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_232), .A2(n_200), .B1(n_204), .B2(n_242), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_226), .B(n_200), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_239), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_267), .A2(n_200), .B(n_204), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_288), .A2(n_204), .B(n_263), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_247), .A2(n_204), .B(n_248), .C(n_262), .Y(n_334) );
NOR2xp33_ASAP7_75t_R g335 ( .A(n_245), .B(n_261), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_259), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_229), .A2(n_266), .B(n_274), .Y(n_337) );
INVx11_ASAP7_75t_L g338 ( .A(n_265), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_261), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_269), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_237), .B(n_257), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_335), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_337), .A2(n_242), .B(n_229), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_294), .A2(n_251), .B1(n_233), .B2(n_237), .C(n_257), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_305), .A2(n_242), .B1(n_283), .B2(n_233), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_290), .B(n_258), .Y(n_346) );
OAI21xp5_ASAP7_75t_L g347 ( .A1(n_334), .A2(n_264), .B(n_252), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_292), .B(n_280), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_311), .A2(n_279), .B(n_242), .C(n_253), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_305), .B(n_228), .Y(n_350) );
AO21x2_ASAP7_75t_L g351 ( .A1(n_327), .A2(n_277), .B(n_281), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_305), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_339), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g355 ( .A1(n_334), .A2(n_311), .B(n_297), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_308), .A2(n_279), .B1(n_273), .B2(n_264), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_304), .A2(n_270), .B(n_282), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_341), .A2(n_272), .B1(n_285), .B2(n_278), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_310), .Y(n_359) );
BUFx12f_ASAP7_75t_L g360 ( .A(n_300), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_293), .A2(n_272), .B1(n_270), .B2(n_282), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_340), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_298), .A2(n_255), .B(n_321), .C(n_295), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_312), .B(n_314), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_332), .A2(n_329), .B(n_330), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_302), .B(n_324), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_331), .B(n_305), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_336), .B(n_299), .Y(n_368) );
NOR2xp33_ASAP7_75t_SL g369 ( .A(n_325), .B(n_301), .Y(n_369) );
AO32x2_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_307), .A3(n_317), .B1(n_323), .B2(n_309), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_296), .A2(n_291), .B(n_319), .C(n_333), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_336), .B(n_296), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_342), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_346), .B(n_313), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_344), .A2(n_301), .B1(n_306), .B2(n_315), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
OA21x2_ASAP7_75t_L g379 ( .A1(n_355), .A2(n_318), .B(n_303), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_320), .B(n_310), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_374), .B(n_310), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_374), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_362), .B(n_310), .Y(n_383) );
OR2x6_ASAP7_75t_L g384 ( .A(n_345), .B(n_326), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g385 ( .A1(n_363), .A2(n_326), .B1(n_338), .B2(n_348), .C(n_358), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_362), .B(n_326), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_342), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_352), .A2(n_326), .B(n_351), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_364), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_368), .B(n_366), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_358), .A2(n_343), .B(n_372), .C(n_373), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_368), .B(n_366), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_349), .A2(n_357), .B(n_351), .Y(n_393) );
BUFx4f_ASAP7_75t_L g394 ( .A(n_369), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_356), .A2(n_347), .B(n_361), .C(n_365), .Y(n_395) );
CKINVDCx6p67_ASAP7_75t_R g396 ( .A(n_360), .Y(n_396) );
AO31x2_ASAP7_75t_L g397 ( .A1(n_370), .A2(n_351), .A3(n_365), .B(n_359), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_354), .B(n_371), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_359), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_370), .B(n_364), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_382), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_381), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_382), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_394), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_402), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_399), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_376), .A2(n_369), .B1(n_353), .B2(n_350), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_390), .B(n_353), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_392), .B(n_350), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_400), .B(n_350), .Y(n_412) );
NAND2x1_ASAP7_75t_L g413 ( .A(n_378), .B(n_359), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_393), .A2(n_370), .B(n_359), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_389), .B(n_350), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_401), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_389), .B(n_370), .Y(n_420) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_391), .A2(n_370), .B(n_360), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_399), .Y(n_422) );
OR2x6_ASAP7_75t_L g423 ( .A(n_384), .B(n_394), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_385), .A2(n_394), .B1(n_377), .B2(n_384), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_381), .B(n_386), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_397), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_384), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_395), .B(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
AOI211xp5_ASAP7_75t_L g433 ( .A1(n_398), .A2(n_387), .B(n_396), .C(n_394), .Y(n_433) );
INVx3_ASAP7_75t_SL g434 ( .A(n_396), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_435), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_428), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_420), .B(n_397), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_420), .B(n_397), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_431), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_428), .B(n_397), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_432), .B(n_388), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_418), .B(n_388), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_432), .B(n_388), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_436), .B(n_380), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_436), .B(n_380), .Y(n_447) );
INVxp67_ASAP7_75t_L g448 ( .A(n_419), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_418), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_407), .B(n_380), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_435), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
NAND2x1_ASAP7_75t_L g455 ( .A(n_423), .B(n_384), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_416), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_425), .B(n_384), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_408), .B(n_378), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_403), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_410), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_427), .B(n_378), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
BUFx2_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_405), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_431), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_425), .B(n_379), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_423), .B(n_379), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_408), .B(n_379), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_434), .B(n_387), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_405), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_421), .B(n_379), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_408), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_417), .Y(n_476) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_421), .A2(n_375), .B(n_414), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_417), .B(n_422), .Y(n_478) );
BUFx12f_ASAP7_75t_L g479 ( .A(n_434), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_427), .B(n_404), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_404), .B(n_426), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_417), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_422), .B(n_414), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_410), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_439), .B(n_429), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_451), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_429), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_449), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_439), .B(n_414), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_466), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_440), .B(n_430), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_440), .B(n_430), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_466), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_484), .B(n_415), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_469), .B(n_423), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_448), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_441), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_448), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_440), .B(n_422), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_480), .B(n_415), .Y(n_503) );
INVx4_ASAP7_75t_L g504 ( .A(n_479), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_460), .B(n_411), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_479), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_463), .B(n_411), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_480), .B(n_404), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_457), .B(n_404), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_457), .B(n_426), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_472), .B(n_426), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_472), .B(n_412), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_479), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
AND2x4_ASAP7_75t_SL g517 ( .A(n_461), .B(n_412), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_471), .B(n_434), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_437), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_478), .B(n_433), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_450), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_442), .B(n_426), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_461), .B(n_409), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_441), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_441), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_437), .B(n_433), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_442), .B(n_406), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_442), .B(n_406), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_437), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_444), .B(n_424), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_443), .B(n_406), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_450), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_478), .B(n_409), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_462), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_462), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_443), .B(n_413), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_443), .B(n_413), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_445), .B(n_446), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g540 ( .A1(n_473), .A2(n_469), .B(n_465), .C(n_464), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_539), .B(n_465), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_499), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_501), .Y(n_543) );
BUFx2_ASAP7_75t_L g544 ( .A(n_504), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_504), .B(n_453), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_486), .B(n_464), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_508), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_539), .B(n_445), .Y(n_549) );
NAND2x1_ASAP7_75t_L g550 ( .A(n_504), .B(n_469), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_535), .B(n_467), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_503), .B(n_467), .Y(n_552) );
INVxp67_ASAP7_75t_SL g553 ( .A(n_536), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_491), .B(n_445), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_495), .B(n_446), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_503), .B(n_467), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_526), .A2(n_455), .B1(n_469), .B2(n_477), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_495), .B(n_446), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_492), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_494), .B(n_462), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_494), .B(n_502), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_491), .B(n_447), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_502), .B(n_447), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_493), .B(n_447), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_496), .B(n_470), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_487), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_505), .B(n_444), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_519), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_497), .B(n_475), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_522), .B(n_469), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_515), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_540), .B(n_473), .C(n_481), .D(n_468), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_475), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_507), .B(n_470), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_485), .B(n_453), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_485), .B(n_453), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_506), .B(n_481), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_488), .B(n_474), .Y(n_583) );
NOR2xp67_ASAP7_75t_SL g584 ( .A(n_514), .B(n_474), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_522), .B(n_483), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_514), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_532), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_509), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_527), .B(n_483), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_527), .B(n_483), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_510), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_528), .B(n_452), .Y(n_592) );
NOR2x1_ASAP7_75t_L g593 ( .A(n_544), .B(n_526), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_545), .B(n_506), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_547), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_564), .B(n_488), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_572), .B(n_498), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_557), .A2(n_538), .B(n_523), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_591), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_588), .B(n_530), .Y(n_600) );
INVxp33_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_542), .Y(n_602) );
INVxp67_ASAP7_75t_SL g603 ( .A(n_553), .Y(n_603) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_553), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_543), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_559), .B(n_518), .C(n_530), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_548), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_560), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_572), .B(n_498), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_554), .B(n_528), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_554), .B(n_520), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_568), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_586), .B(n_529), .C(n_455), .Y(n_614) );
OAI321xp33_ASAP7_75t_L g615 ( .A1(n_575), .A2(n_533), .A3(n_537), .B1(n_510), .B2(n_511), .C(n_513), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_563), .A2(n_517), .B1(n_498), .B2(n_511), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_537), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_592), .B(n_531), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_559), .B(n_517), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_569), .B(n_531), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_576), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_584), .A2(n_512), .B(n_468), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_549), .B(n_500), .Y(n_625) );
OAI32xp33_ASAP7_75t_L g626 ( .A1(n_555), .A2(n_512), .A3(n_474), .B1(n_500), .B2(n_525), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_561), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_570), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_581), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_629), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_615), .A2(n_546), .B1(n_582), .B2(n_558), .C(n_541), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_598), .B(n_592), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_599), .B(n_590), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_607), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_594), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_608), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_601), .A2(n_570), .B1(n_562), .B2(n_578), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_600), .B(n_590), .Y(n_638) );
XOR2xp5_ASAP7_75t_L g639 ( .A(n_606), .B(n_571), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_611), .B(n_582), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_614), .A2(n_561), .B(n_477), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_610), .B(n_546), .Y(n_642) );
AOI32xp33_ASAP7_75t_L g643 ( .A1(n_601), .A2(n_579), .A3(n_580), .B1(n_583), .B2(n_565), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_612), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_618), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_597), .B(n_585), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_594), .A2(n_567), .B(n_566), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_593), .A2(n_556), .B1(n_552), .B2(n_577), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_603), .A2(n_477), .B(n_534), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_603), .B(n_565), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_619), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_604), .B(n_589), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_641), .A2(n_620), .B(n_624), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_635), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_648), .A2(n_604), .B(n_628), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_631), .B(n_596), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_650), .A2(n_628), .B(n_616), .C(n_620), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_630), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_639), .A2(n_632), .B1(n_637), .B2(n_640), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_647), .A2(n_602), .B1(n_605), .B2(n_595), .C(n_622), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_642), .B(n_597), .Y(n_661) );
AOI32xp33_ASAP7_75t_L g662 ( .A1(n_651), .A2(n_609), .A3(n_617), .B1(n_613), .B2(n_589), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_634), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_646), .B(n_609), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_636), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_643), .A2(n_626), .B1(n_623), .B2(n_621), .C(n_613), .Y(n_666) );
AOI221xp5_ASAP7_75t_SL g667 ( .A1(n_666), .A2(n_641), .B1(n_652), .B2(n_649), .C(n_644), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_653), .A2(n_649), .B1(n_645), .B2(n_633), .C(n_638), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_655), .B(n_627), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_658), .Y(n_670) );
OAI21x1_ASAP7_75t_SL g671 ( .A1(n_660), .A2(n_627), .B(n_625), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_659), .B(n_587), .C(n_454), .D(n_456), .Y(n_672) );
NOR4xp25_ASAP7_75t_L g673 ( .A(n_657), .B(n_454), .C(n_456), .D(n_585), .Y(n_673) );
AOI21xp5_ASAP7_75t_SL g674 ( .A1(n_660), .A2(n_477), .B(n_525), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g675 ( .A1(n_673), .A2(n_656), .B(n_654), .C(n_661), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_668), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_664), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_667), .B(n_452), .C(n_470), .Y(n_677) );
NOR2xp33_ASAP7_75t_SL g678 ( .A(n_669), .B(n_458), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_677), .Y(n_679) );
NOR3xp33_ASAP7_75t_SL g680 ( .A(n_676), .B(n_672), .C(n_670), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_675), .A2(n_674), .B(n_671), .C(n_452), .Y(n_681) );
OAI22xp5_ASAP7_75t_SL g682 ( .A1(n_679), .A2(n_678), .B1(n_524), .B2(n_534), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_680), .B(n_524), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_683), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_684), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_681), .B(n_682), .Y(n_686) );
OA21x2_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_482), .B(n_476), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_687), .A2(n_458), .B1(n_476), .B2(n_482), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_458), .B1(n_476), .B2(n_482), .Y(n_689) );
endmodule