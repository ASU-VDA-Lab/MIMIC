module real_jpeg_7073_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_2),
.B(n_157),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_2),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_206),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_52),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_61),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_3),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_3),
.B(n_83),
.Y(n_326)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_5),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_5),
.B(n_134),
.Y(n_133)
);

NAND2x1p5_ASAP7_75t_L g178 ( 
.A(n_5),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_5),
.B(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_7),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_8),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_8),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_8),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_9),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_9),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_9),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_9),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_9),
.B(n_83),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_9),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_10),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_10),
.B(n_328),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_11),
.Y(n_136)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_11),
.Y(n_247)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_13),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_13),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_13),
.B(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_13),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_13),
.B(n_222),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_14),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_14),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_14),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_15),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_16),
.B(n_37),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_16),
.B(n_30),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_17),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_17),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_17),
.B(n_80),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_17),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_17),
.B(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_308),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_258),
.B(n_307),
.Y(n_19)
);

AOI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_215),
.B(n_257),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_164),
.B(n_214),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_128),
.B(n_163),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_91),
.B(n_127),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_69),
.B(n_90),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_46),
.B(n_68),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_42),
.B(n_45),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_38),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_31),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_40),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_41),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_60),
.C(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_54),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_67),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_89),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_89),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_77),
.C(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_75),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_111),
.C(n_112),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_85),
.Y(n_243)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_94),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_110),
.C(n_113),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_98),
.C(n_102),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_122),
.C(n_125),
.Y(n_161)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_120),
.Y(n_300)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_121),
.Y(n_254)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_121),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_122),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_162),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_131),
.B(n_138),
.C(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_188),
.C(n_189),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_152),
.C(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_146),
.C(n_148),
.Y(n_185)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_149),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_160),
.B2(n_161),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_156),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_212),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_212),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_186),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_167),
.B(n_168),
.C(n_186),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_182),
.B2(n_183),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_169),
.B(n_234),
.C(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_171),
.B(n_176),
.C(n_181),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_180),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_191),
.C(n_211),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_199),
.B1(n_210),
.B2(n_211),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.B(n_198),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_195),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_198),
.B(n_219),
.C(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_205),
.C(n_208),
.Y(n_255)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_205),
.Y(n_209)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_256),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_256),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_232),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_231),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_231),
.C(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_228),
.B2(n_230),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_221),
.B(n_225),
.C(n_302),
.Y(n_301)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_237),
.C(n_248),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_242),
.C(n_244),
.Y(n_275)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_251),
.C(n_294),
.Y(n_293)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_255),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_305),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_290),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_262),
.B(n_290),
.C(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_273),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_274),
.C(n_277),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_264),
.B(n_269),
.C(n_270),
.Y(n_343)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_288),
.B2(n_289),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_288),
.C(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_289),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_295),
.B1(n_303),
.B2(n_304),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_304),
.C(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_299),
.C(n_301),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_346),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_344),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_344),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_330),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_321),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);


endmodule