module real_jpeg_3022_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_200;
wire n_48;
wire n_56;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_213;
wire n_244;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_2),
.A2(n_28),
.B1(n_39),
.B2(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_68),
.B1(n_70),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_3),
.A2(n_39),
.B1(n_41),
.B2(n_81),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_5),
.B(n_129),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_39),
.C(n_54),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_5),
.B(n_53),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_5),
.B(n_27),
.C(n_44),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_39),
.B1(n_41),
.B2(n_167),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_32),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_49),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_167),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_10),
.A2(n_48),
.B1(n_57),
.B2(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_48),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_39),
.B1(n_41),
.B2(n_67),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_67),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_14),
.A2(n_61),
.B1(n_68),
.B2(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_14),
.A2(n_39),
.B1(n_41),
.B2(n_61),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_14),
.A2(n_27),
.B1(n_29),
.B2(n_61),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_15),
.A2(n_68),
.B1(n_70),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_15),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_128),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_15),
.A2(n_39),
.B1(n_41),
.B2(n_128),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_128),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_109),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.C(n_64),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_22),
.A2(n_23),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_24),
.A2(n_35),
.B1(n_36),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_24),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_26),
.A2(n_32),
.B1(n_97),
.B2(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_31),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_27),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_30),
.A2(n_31),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_30),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_30),
.A2(n_31),
.B1(n_147),
.B2(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_30),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_30),
.A2(n_31),
.B1(n_192),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_31),
.A2(n_146),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_31),
.B(n_161),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_32),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_32),
.A2(n_160),
.B(n_217),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_39),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_42),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_42),
.B(n_153),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_86),
.B1(n_87),
.B2(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_46),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_46),
.A2(n_174),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_46),
.A2(n_86),
.B1(n_150),
.B2(n_200),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_49),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_50),
.B(n_64),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_62),
.B1(n_63),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_51),
.A2(n_62),
.B1(n_140),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_51),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_51),
.A2(n_171),
.B(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_52),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_53),
.B(n_125),
.Y(n_233)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_58),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_57),
.B(n_157),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_57),
.B(n_75),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_58),
.A2(n_68),
.A3(n_74),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_62),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_62),
.A2(n_124),
.B(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_78),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_72),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_68),
.A2(n_71),
.B(n_167),
.C(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_68),
.B(n_167),
.Y(n_168)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_73),
.A2(n_102),
.B(n_253),
.Y(n_252)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_79),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_92),
.B2(n_93),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_91),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_86),
.A2(n_152),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_105),
.B2(n_108),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_104),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_104),
.B1(n_106),
.B2(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_97),
.A2(n_167),
.B(n_194),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_110),
.B(n_113),
.Y(n_278)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_115),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_116),
.A2(n_117),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_118),
.B(n_120),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_126),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_127),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_275),
.B(n_279),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_244),
.B(n_272),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_186),
.B(n_243),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_162),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_137),
.B(n_162),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.C(n_154),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_138),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_142),
.C(n_145),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_148),
.B(n_154),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_163),
.B(n_177),
.C(n_185),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_175),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_164),
.B(n_170),
.C(n_172),
.Y(n_257)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_183),
.Y(n_248)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_238),
.B(n_242),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_227),
.B(n_237),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_209),
.B(n_226),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_203),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_195),
.B1(n_201),
.B2(n_202),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_198),
.C(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_220),
.B(n_225),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B(n_219),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_223),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_229),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_259),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_258),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_256),
.C(n_257),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.C(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_271),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_271),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_265),
.C(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_277),
.Y(n_279)
);


endmodule