module fake_jpeg_1558_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_58),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_61),
.Y(n_186)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_65),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_18),
.B(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_71),
.Y(n_160)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_78),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_80),
.Y(n_198)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_23),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_32),
.B(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_99),
.B(n_120),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_55),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_106),
.Y(n_139)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_108),
.B(n_111),
.Y(n_193)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_41),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_116),
.Y(n_128)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_18),
.B(n_16),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_44),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_126),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_58),
.B(n_86),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_136),
.B(n_161),
.C(n_122),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_65),
.A2(n_36),
.B1(n_53),
.B2(n_39),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_142),
.A2(n_157),
.B1(n_163),
.B2(n_189),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_39),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_152),
.B(n_155),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_66),
.B(n_36),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_82),
.A2(n_53),
.B1(n_55),
.B2(n_38),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_158),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_38),
.C(n_37),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_96),
.A2(n_108),
.B1(n_21),
.B2(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_50),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_165),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_48),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_48),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_168),
.B(n_176),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_92),
.A2(n_44),
.B1(n_43),
.B2(n_37),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_181),
.B1(n_197),
.B2(n_199),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_179),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_56),
.B(n_0),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_93),
.A2(n_34),
.B1(n_31),
.B2(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_59),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_9),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_119),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_188),
.B(n_162),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_94),
.A2(n_34),
.B1(n_31),
.B2(n_5),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_98),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_60),
.A2(n_34),
.B1(n_4),
.B2(n_5),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_61),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_202),
.B1(n_197),
.B2(n_199),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_70),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_208),
.B(n_211),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_209),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_122),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_139),
.A2(n_73),
.B1(n_80),
.B2(n_78),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_215),
.B(n_225),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_135),
.B(n_76),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_216),
.B(n_261),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_139),
.A2(n_75),
.B1(n_100),
.B2(n_11),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_217),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_239),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_154),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_128),
.B(n_9),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_221),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_154),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_170),
.B(n_137),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_159),
.B1(n_140),
.B2(n_130),
.Y(n_226)
);

OAI22x1_ASAP7_75t_SL g306 ( 
.A1(n_226),
.A2(n_232),
.B1(n_246),
.B2(n_249),
.Y(n_306)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_227),
.Y(n_314)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_136),
.A2(n_12),
.B1(n_15),
.B2(n_167),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_230),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_286)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_126),
.A2(n_145),
.B1(n_143),
.B2(n_189),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_233),
.A2(n_238),
.B1(n_269),
.B2(n_270),
.Y(n_277)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_187),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_235),
.B(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_174),
.A2(n_142),
.B1(n_157),
.B2(n_129),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_245),
.A2(n_207),
.B1(n_206),
.B2(n_251),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_246),
.Y(n_318)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_190),
.A2(n_196),
.B1(n_163),
.B2(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_248),
.A2(n_245),
.B1(n_210),
.B2(n_207),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_123),
.A2(n_171),
.B(n_131),
.C(n_192),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_263),
.Y(n_278)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_251),
.Y(n_293)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_169),
.A2(n_193),
.B1(n_194),
.B2(n_144),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_150),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_253),
.Y(n_300)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_256),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_147),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_289)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_196),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_125),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_149),
.B(n_173),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_133),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_134),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_186),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_185),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_267),
.B(n_271),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_153),
.A2(n_195),
.B1(n_134),
.B2(n_180),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_144),
.A2(n_198),
.B1(n_151),
.B2(n_180),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_233),
.A2(n_162),
.B1(n_186),
.B2(n_191),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_287),
.A2(n_297),
.B1(n_306),
.B2(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_208),
.B(n_191),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_292),
.A2(n_290),
.B(n_276),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_216),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_303),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_226),
.A2(n_268),
.B1(n_229),
.B2(n_221),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_237),
.C(n_240),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_308),
.C(n_321),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_221),
.B(n_218),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_305),
.A2(n_279),
.B1(n_286),
.B2(n_281),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_227),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_282),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_207),
.B(n_255),
.C(n_212),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_207),
.A2(n_228),
.B(n_214),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_290),
.B(n_295),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_313),
.A2(n_260),
.B1(n_234),
.B2(n_241),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_262),
.A2(n_264),
.B1(n_263),
.B2(n_209),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_204),
.B(n_231),
.C(n_258),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_310),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_323),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_335),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_292),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_331),
.C(n_324),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_342),
.B1(n_344),
.B2(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_296),
.B(n_222),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_329),
.B(n_333),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_257),
.C(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_294),
.B(n_222),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_278),
.A2(n_254),
.B(n_244),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_334),
.A2(n_346),
.B(n_357),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_311),
.Y(n_335)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

BUFx24_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_337),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_273),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_339),
.B(n_359),
.Y(n_369)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_305),
.A2(n_256),
.B1(n_205),
.B2(n_242),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_313),
.A2(n_308),
.B1(n_312),
.B2(n_277),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_278),
.A2(n_297),
.B(n_283),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_279),
.A2(n_301),
.B1(n_287),
.B2(n_317),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_307),
.B1(n_303),
.B2(n_309),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_349),
.A2(n_351),
.B1(n_360),
.B2(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_361),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_291),
.A2(n_300),
.B1(n_289),
.B2(n_321),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_314),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_352),
.Y(n_374)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_284),
.Y(n_353)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_288),
.A2(n_322),
.B1(n_293),
.B2(n_275),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_274),
.B1(n_280),
.B2(n_319),
.Y(n_370)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_316),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_322),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_302),
.A2(n_315),
.B1(n_275),
.B2(n_276),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_274),
.A2(n_280),
.B(n_295),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_330),
.B(n_316),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_355),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_366),
.A2(n_342),
.B1(n_327),
.B2(n_354),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_381),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_386),
.B1(n_387),
.B2(n_360),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_325),
.B(n_319),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_372),
.B(n_383),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_326),
.B(n_338),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_373),
.B(n_389),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_352),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_350),
.B(n_338),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_340),
.A2(n_346),
.B1(n_330),
.B2(n_344),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_340),
.A2(n_329),
.B1(n_357),
.B2(n_349),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_324),
.B(n_331),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_352),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_333),
.C(n_351),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_337),
.C(n_386),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_395),
.A2(n_399),
.B1(n_400),
.B2(n_416),
.Y(n_431)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_398),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_364),
.A2(n_332),
.B1(n_341),
.B2(n_335),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_369),
.B(n_356),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_401),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_413),
.C(n_418),
.Y(n_429)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_404),
.B(n_405),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_364),
.A2(n_361),
.B1(n_336),
.B2(n_343),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_406),
.A2(n_408),
.B1(n_419),
.B2(n_363),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_371),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_417),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_366),
.A2(n_353),
.B1(n_328),
.B2(n_323),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_337),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_411),
.Y(n_421)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_376),
.Y(n_410)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_410),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_337),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_392),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_391),
.C(n_367),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_379),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_393),
.B1(n_379),
.B2(n_384),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_363),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_365),
.B(n_393),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_384),
.A2(n_381),
.B1(n_362),
.B2(n_374),
.Y(n_419)
);

OA22x2_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_370),
.B1(n_392),
.B2(n_388),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_416),
.A2(n_365),
.B(n_385),
.Y(n_422)
);

XOR2x1_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_419),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_409),
.C(n_412),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_424),
.B(n_430),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_398),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_375),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_397),
.B(n_382),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_434),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_437),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_441),
.Y(n_454)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_415),
.Y(n_442)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_394),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_443),
.B(n_396),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_446),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_413),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_431),
.A2(n_400),
.B1(n_404),
.B2(n_396),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_447),
.A2(n_439),
.B1(n_431),
.B2(n_422),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_452),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_432),
.B(n_418),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_453),
.B(n_462),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_460),
.Y(n_471)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_440),
.Y(n_457)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_459),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_444),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_433),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_434),
.B(n_429),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_396),
.C(n_399),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_463),
.B(n_462),
.C(n_446),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_474),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_466),
.A2(n_450),
.B1(n_455),
.B2(n_447),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_438),
.C(n_421),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_467),
.B(n_472),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_445),
.B(n_443),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_475),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_463),
.A2(n_439),
.B(n_427),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_476),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_427),
.C(n_426),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_452),
.C(n_420),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_482),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_467),
.C(n_474),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_SL g497 ( 
.A(n_481),
.B(n_484),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_371),
.Y(n_483)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_483),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_449),
.C(n_453),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_471),
.A2(n_452),
.B(n_426),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_488),
.B(n_478),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_375),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_482),
.B(n_464),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_480),
.Y(n_508)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_479),
.A2(n_466),
.B1(n_473),
.B2(n_478),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_496),
.B(n_498),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_465),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_454),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_499),
.B(n_500),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_486),
.A2(n_448),
.B(n_456),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_481),
.C(n_487),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_503),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_487),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_485),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_507),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_484),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_426),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_500),
.C(n_491),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_512),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_464),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_493),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_513),
.A2(n_435),
.B1(n_441),
.B2(n_425),
.Y(n_517)
);

OAI21x1_ASAP7_75t_SL g516 ( 
.A1(n_514),
.A2(n_505),
.B(n_435),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_516),
.A2(n_517),
.B1(n_428),
.B2(n_436),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g518 ( 
.A(n_509),
.B(n_425),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_518),
.A2(n_514),
.B(n_510),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_519),
.A2(n_520),
.B(n_515),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_428),
.C(n_442),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_420),
.C(n_377),
.Y(n_524)
);

FAx1_ASAP7_75t_SL g525 ( 
.A(n_524),
.B(n_420),
.CI(n_511),
.CON(n_525),
.SN(n_525)
);


endmodule