module fake_jpeg_28569_n_26 (n_3, n_2, n_1, n_0, n_4, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

INVx6_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_8),
.B(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_11),
.B(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_13),
.A2(n_9),
.B1(n_6),
.B2(n_4),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_6),
.B1(n_9),
.B2(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_15),
.B(n_13),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_23),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_22),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_16),
.C(n_10),
.Y(n_26)
);


endmodule