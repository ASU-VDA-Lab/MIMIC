module fake_jpeg_4471_n_126 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_27),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_22),
.B(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_29),
.A2(n_17),
.B1(n_19),
.B2(n_38),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_5),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_29),
.A2(n_17),
.B1(n_19),
.B2(n_26),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_20),
.C(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_34),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_24),
.B1(n_4),
.B2(n_7),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_39),
.B1(n_5),
.B2(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_54),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_24),
.C(n_4),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_4),
.B1(n_52),
.B2(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_55),
.B1(n_42),
.B2(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_50),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_53),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_87),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_50),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_68),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_85),
.B(n_90),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_72),
.B1(n_66),
.B2(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_70),
.B(n_65),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_99),
.B(n_101),
.Y(n_105)
);

NAND2x1_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_106),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_79),
.B(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_82),
.C(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_64),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_99),
.C(n_83),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_96),
.B1(n_95),
.B2(n_84),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_109),
.B1(n_74),
.B2(n_107),
.Y(n_117)
);

NAND2x1_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_94),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_86),
.C(n_74),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_118),
.B(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_113),
.A3(n_110),
.B1(n_115),
.B2(n_112),
.C1(n_80),
.C2(n_41),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_51),
.C(n_102),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_122),
.B(n_81),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule