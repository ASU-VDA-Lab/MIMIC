module fake_jpeg_25022_n_222 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_222);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_18),
.B1(n_19),
.B2(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_27),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_47),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_32),
.C(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_53),
.C(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_24),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_58),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_57),
.B1(n_30),
.B2(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_55),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_32),
.C(n_29),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_25),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_37),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_34),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_19),
.B2(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_11),
.B(n_12),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_68),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_12),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_12),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_47),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_73),
.A2(n_46),
.B1(n_53),
.B2(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_79),
.B1(n_86),
.B2(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_46),
.B1(n_43),
.B2(n_49),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_74),
.Y(n_96)
);

OR2x6_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_54),
.B1(n_43),
.B2(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_73),
.C(n_71),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_95),
.C(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_94),
.B1(n_92),
.B2(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_80),
.B1(n_89),
.B2(n_88),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_20),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_45),
.C(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_70),
.B1(n_59),
.B2(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_85),
.B1(n_58),
.B2(n_67),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_81),
.C(n_87),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_44),
.C(n_28),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_11),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_20),
.B1(n_15),
.B2(n_22),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_118),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_14),
.B(n_22),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_120),
.B1(n_127),
.B2(n_33),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_22),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_97),
.B1(n_90),
.B2(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_123),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_14),
.B1(n_40),
.B2(n_11),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_14),
.B1(n_21),
.B2(n_17),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_67),
.B1(n_40),
.B2(n_11),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_44),
.C(n_67),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_44),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_111),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_132),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_144),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_127),
.B1(n_114),
.B2(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_15),
.B(n_20),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_21),
.B(n_1),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_112),
.B1(n_126),
.B2(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_9),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_112),
.C(n_122),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_9),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_155),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_141),
.B(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_28),
.C(n_25),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_17),
.C(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_7),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_133),
.B1(n_145),
.B2(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_130),
.B1(n_142),
.B2(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_175),
.Y(n_182)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_130),
.B(n_142),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_176),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_149),
.B1(n_147),
.B2(n_131),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_17),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_152),
.C(n_156),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_17),
.C(n_21),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_159),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_157),
.B1(n_162),
.B2(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_37),
.B1(n_5),
.B2(n_8),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_190),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_157),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_168),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_7),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_179),
.C(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_195),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_186),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_175),
.B1(n_177),
.B2(n_37),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_7),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_198),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_204),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_193),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_211),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_199),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_180),
.C(n_8),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_212),
.A2(n_8),
.B(n_10),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_215),
.B(n_207),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_10),
.B(n_1),
.C(n_2),
.D(n_4),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_21),
.B(n_2),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_216),
.B(n_2),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_0),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_0),
.Y(n_222)
);


endmodule