module fake_jpeg_7664_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_61),
.B1(n_69),
.B2(n_31),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_66),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_22),
.B(n_24),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_22),
.B(n_31),
.C(n_24),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_17),
.B1(n_32),
.B2(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_25),
.B1(n_32),
.B2(n_18),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_25),
.B1(n_19),
.B2(n_30),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_33),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_71),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_83),
.B1(n_87),
.B2(n_90),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_32),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_98),
.B(n_72),
.C(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_25),
.B1(n_19),
.B2(n_30),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_26),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_23),
.B(n_29),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_19),
.B1(n_26),
.B2(n_20),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_29),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_28),
.C(n_20),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_15),
.B(n_12),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_99),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_47),
.A2(n_0),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_10),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_55),
.B1(n_29),
.B2(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_105),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_52),
.B1(n_55),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_115),
.B1(n_119),
.B2(n_98),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_109),
.B1(n_4),
.B2(n_5),
.Y(n_149)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_55),
.B(n_63),
.C(n_59),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_73),
.B(n_91),
.Y(n_148)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_113),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_29),
.B1(n_8),
.B2(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_125),
.Y(n_151)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_95),
.B1(n_91),
.B2(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_130),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_94),
.B(n_73),
.C(n_77),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_145),
.Y(n_157)
);

CKINVDCx12_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_92),
.C(n_85),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.C(n_103),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_81),
.C(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_122),
.B(n_104),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_149),
.B(n_119),
.Y(n_159)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_121),
.B(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_158),
.C(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_162),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_125),
.C(n_109),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_135),
.B1(n_149),
.B2(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_117),
.C(n_127),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_114),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_139),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_141),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_179),
.C(n_185),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_182),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_148),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_184),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_116),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_184),
.B(n_172),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_136),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_194),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_159),
.B1(n_155),
.B2(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_154),
.C(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_195),
.C(n_181),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_158),
.C(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_143),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_199),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_180),
.B(n_173),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_192),
.B(n_190),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_202),
.C(n_165),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_162),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_210),
.C(n_211),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_195),
.B1(n_191),
.B2(n_131),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_164),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_144),
.Y(n_218)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_204),
.B1(n_205),
.B2(n_150),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_217),
.B(n_205),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.C(n_211),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_216),
.A2(n_214),
.B(n_212),
.C(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_201),
.C(n_161),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_123),
.B(n_105),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_11),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule