module fake_aes_5542_n_30 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_7), .B(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_3), .B(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
OAI22xp33_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_4), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_14), .B(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx2_ASAP7_75t_SL g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OAI21xp33_ASAP7_75t_SL g25 ( .A1(n_23), .A2(n_20), .B(n_16), .Y(n_25) );
NAND2x1p5_ASAP7_75t_L g26 ( .A(n_24), .B(n_16), .Y(n_26) );
NAND4xp75_ASAP7_75t_L g27 ( .A(n_25), .B(n_19), .C(n_0), .D(n_13), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
OAI22xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .B1(n_19), .B2(n_8), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
endmodule