module real_aes_2260_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_0), .B(n_500), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_1), .A2(n_502), .B(n_503), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_2), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_3), .B(n_178), .Y(n_536) );
INVx1_ASAP7_75t_L g133 ( .A(n_4), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_5), .B(n_142), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_6), .B(n_178), .Y(n_524) );
INVx1_ASAP7_75t_L g188 ( .A(n_7), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g827 ( .A(n_8), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_9), .Y(n_204) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_10), .B(n_175), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_11), .A2(n_38), .B1(n_812), .B2(n_813), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_11), .Y(n_813) );
INVx2_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
AOI221x1_ASAP7_75t_L g581 ( .A1(n_13), .A2(n_27), .B1(n_500), .B2(n_502), .C(n_582), .Y(n_581) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_14), .Y(n_112) );
AND3x1_ASAP7_75t_L g824 ( .A(n_14), .B(n_41), .C(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_15), .B(n_500), .Y(n_553) );
INVx1_ASAP7_75t_L g176 ( .A(n_16), .Y(n_176) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_17), .A2(n_164), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_18), .B(n_218), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_19), .B(n_178), .Y(n_513) );
AO21x1_ASAP7_75t_L g531 ( .A1(n_20), .A2(n_500), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g116 ( .A(n_21), .Y(n_116) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_22), .A2(n_59), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_22), .Y(n_793) );
INVx1_ASAP7_75t_L g173 ( .A(n_23), .Y(n_173) );
INVx1_ASAP7_75t_SL g248 ( .A(n_24), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_25), .Y(n_804) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_26), .B(n_153), .Y(n_152) );
AOI33xp33_ASAP7_75t_L g225 ( .A1(n_28), .A2(n_55), .A3(n_130), .B1(n_148), .B2(n_226), .B3(n_227), .Y(n_225) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_29), .B(n_178), .Y(n_574) );
NAND2x1_ASAP7_75t_L g523 ( .A(n_30), .B(n_175), .Y(n_523) );
INVx1_ASAP7_75t_L g197 ( .A(n_31), .Y(n_197) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_32), .A2(n_88), .B(n_141), .Y(n_140) );
OR2x2_ASAP7_75t_L g143 ( .A(n_32), .B(n_88), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_33), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_34), .B(n_186), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_35), .B(n_175), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_36), .B(n_178), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_37), .B(n_175), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_38), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_39), .A2(n_502), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g136 ( .A(n_40), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g147 ( .A(n_40), .Y(n_147) );
AND2x2_ASAP7_75t_L g162 ( .A(n_40), .B(n_133), .Y(n_162) );
OR2x6_ASAP7_75t_L g114 ( .A(n_41), .B(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_42), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_43), .B(n_500), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_44), .B(n_186), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_45), .A2(n_127), .B1(n_139), .B2(n_142), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_46), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_47), .B(n_153), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_48), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_49), .B(n_175), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_50), .B(n_164), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_51), .B(n_153), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_52), .A2(n_502), .B(n_522), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_53), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_54), .B(n_175), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_56), .B(n_153), .Y(n_216) );
INVx1_ASAP7_75t_L g131 ( .A(n_57), .Y(n_131) );
INVx1_ASAP7_75t_L g155 ( .A(n_57), .Y(n_155) );
AND2x2_ASAP7_75t_L g217 ( .A(n_58), .B(n_218), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_59), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g185 ( .A1(n_60), .A2(n_77), .B1(n_145), .B2(n_186), .C(n_187), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_61), .B(n_186), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_62), .B(n_178), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_63), .B(n_139), .Y(n_206) );
AOI21xp5_ASAP7_75t_SL g236 ( .A1(n_64), .A2(n_145), .B(n_237), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_65), .A2(n_502), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g169 ( .A(n_66), .Y(n_169) );
AO21x1_ASAP7_75t_L g533 ( .A1(n_67), .A2(n_502), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_68), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g215 ( .A(n_69), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_70), .B(n_500), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_71), .A2(n_145), .B(n_214), .Y(n_213) );
INVxp33_ASAP7_75t_L g829 ( .A(n_72), .Y(n_829) );
AND2x2_ASAP7_75t_L g547 ( .A(n_73), .B(n_219), .Y(n_547) );
INVx1_ASAP7_75t_L g137 ( .A(n_74), .Y(n_137) );
INVx1_ASAP7_75t_L g157 ( .A(n_74), .Y(n_157) );
AND2x2_ASAP7_75t_L g526 ( .A(n_75), .B(n_193), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_76), .B(n_186), .Y(n_228) );
AND2x2_ASAP7_75t_L g250 ( .A(n_78), .B(n_193), .Y(n_250) );
INVx1_ASAP7_75t_L g170 ( .A(n_79), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_80), .A2(n_145), .B(n_247), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_81), .A2(n_145), .B(n_151), .C(n_163), .Y(n_144) );
INVx1_ASAP7_75t_L g117 ( .A(n_82), .Y(n_117) );
AND2x2_ASAP7_75t_L g497 ( .A(n_83), .B(n_193), .Y(n_497) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_84), .B(n_193), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_85), .B(n_500), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_86), .A2(n_145), .B1(n_223), .B2(n_224), .Y(n_222) );
AND2x2_ASAP7_75t_L g532 ( .A(n_87), .B(n_142), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_89), .B(n_175), .Y(n_514) );
AND2x2_ASAP7_75t_L g577 ( .A(n_90), .B(n_193), .Y(n_577) );
INVx1_ASAP7_75t_L g238 ( .A(n_91), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_92), .B(n_178), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_93), .A2(n_502), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_94), .B(n_175), .Y(n_583) );
AND2x2_ASAP7_75t_L g229 ( .A(n_95), .B(n_193), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_96), .B(n_178), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_97), .A2(n_195), .B(n_196), .C(n_198), .Y(n_194) );
BUFx2_ASAP7_75t_L g105 ( .A(n_98), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_99), .A2(n_502), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_100), .B(n_153), .Y(n_239) );
AOI21xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_818), .B(n_828), .Y(n_101) );
AO21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_106), .B(n_807), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_105), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g106 ( .A(n_107), .B(n_802), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_791), .B(n_794), .Y(n_107) );
OAI22xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_118), .B1(n_490), .B2(n_789), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_110), .A2(n_118), .B1(n_490), .B2(n_796), .Y(n_795) );
CKINVDCx11_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
OR2x6_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x6_ASAP7_75t_SL g790 ( .A(n_112), .B(n_114), .Y(n_790) );
OR2x2_ASAP7_75t_L g800 ( .A(n_112), .B(n_114), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_112), .B(n_113), .Y(n_806) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g823 ( .A(n_115), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_424), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_347), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_294), .C(n_327), .Y(n_120) );
AOI211xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_251), .B(n_260), .C(n_284), .Y(n_121) );
OAI21xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_180), .B(n_230), .Y(n_122) );
OR2x2_ASAP7_75t_L g304 ( .A(n_123), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g459 ( .A(n_123), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI22xp33_ASAP7_75t_SL g349 ( .A1(n_124), .A2(n_350), .B1(n_354), .B2(n_356), .Y(n_349) );
AND2x2_ASAP7_75t_L g386 ( .A(n_124), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_165), .Y(n_124) );
INVx1_ASAP7_75t_L g283 ( .A(n_125), .Y(n_283) );
AND2x4_ASAP7_75t_L g300 ( .A(n_125), .B(n_281), .Y(n_300) );
INVx2_ASAP7_75t_L g322 ( .A(n_125), .Y(n_322) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_125), .Y(n_405) );
AND2x2_ASAP7_75t_L g476 ( .A(n_125), .B(n_233), .Y(n_476) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_144), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_134), .C(n_138), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x4_ASAP7_75t_L g186 ( .A(n_129), .B(n_135), .Y(n_186) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
OR2x6_ASAP7_75t_L g160 ( .A(n_130), .B(n_149), .Y(n_160) );
INVxp33_ASAP7_75t_L g226 ( .A(n_130), .Y(n_226) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g150 ( .A(n_131), .B(n_133), .Y(n_150) );
AND2x4_ASAP7_75t_L g178 ( .A(n_131), .B(n_156), .Y(n_178) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x6_ASAP7_75t_L g502 ( .A(n_136), .B(n_150), .Y(n_502) );
INVx2_ASAP7_75t_L g149 ( .A(n_137), .Y(n_149) );
AND2x6_ASAP7_75t_L g175 ( .A(n_137), .B(n_154), .Y(n_175) );
INVx4_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_139), .B(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
AND2x4_ASAP7_75t_L g142 ( .A(n_141), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_141), .B(n_143), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_142), .B(n_161), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_142), .A2(n_236), .B(n_240), .Y(n_235) );
INVx1_ASAP7_75t_SL g509 ( .A(n_142), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_142), .B(n_538), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_142), .A2(n_553), .B(n_554), .Y(n_552) );
INVxp67_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NOR2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx1_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_158), .B(n_161), .Y(n_151) );
INVx1_ASAP7_75t_L g171 ( .A(n_153), .Y(n_171) );
AND2x4_ASAP7_75t_L g500 ( .A(n_153), .B(n_162), .Y(n_500) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_160), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_SL g187 ( .A1(n_160), .A2(n_161), .B(n_188), .C(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_161), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_160), .A2(n_161), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_SL g247 ( .A1(n_160), .A2(n_161), .B(n_248), .C(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g223 ( .A(n_161), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_161), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_161), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_161), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_161), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_161), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_161), .A2(n_556), .B(n_557), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_161), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_161), .A2(n_583), .B(n_584), .Y(n_582) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_163), .A2(n_221), .B(n_229), .Y(n_220) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_163), .A2(n_221), .B(n_229), .Y(n_265) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_164), .A2(n_185), .B(n_190), .Y(n_184) );
AND2x2_ASAP7_75t_L g241 ( .A(n_165), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
INVx3_ASAP7_75t_L g281 ( .A(n_165), .Y(n_281) );
AND2x4_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_179), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_171), .B(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B1(n_176), .B2(n_177), .Y(n_172) );
INVxp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVxp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_180), .A2(n_471), .B1(n_473), .B2(n_475), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_180), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_208), .Y(n_181) );
INVx3_ASAP7_75t_L g254 ( .A(n_182), .Y(n_254) );
AND2x2_ASAP7_75t_L g262 ( .A(n_182), .B(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_182), .Y(n_292) );
NAND2x1_ASAP7_75t_SL g486 ( .A(n_182), .B(n_253), .Y(n_486) );
AND2x4_ASAP7_75t_L g182 ( .A(n_183), .B(n_191), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_184), .B(n_265), .Y(n_277) );
AND2x2_ASAP7_75t_L g290 ( .A(n_184), .B(n_191), .Y(n_290) );
AND2x4_ASAP7_75t_L g297 ( .A(n_184), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_184), .Y(n_346) );
INVxp67_ASAP7_75t_L g353 ( .A(n_184), .Y(n_353) );
INVx1_ASAP7_75t_L g358 ( .A(n_184), .Y(n_358) );
INVx1_ASAP7_75t_L g207 ( .A(n_186), .Y(n_207) );
INVx1_ASAP7_75t_L g257 ( .A(n_191), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_191), .B(n_267), .Y(n_276) );
INVx2_ASAP7_75t_L g344 ( .A(n_191), .Y(n_344) );
INVx1_ASAP7_75t_L g383 ( .A(n_191), .Y(n_383) );
OR2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_201), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B1(n_199), .B2(n_200), .Y(n_192) );
INVx3_ASAP7_75t_L g200 ( .A(n_193), .Y(n_200) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_200), .A2(n_211), .B(n_217), .Y(n_210) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_200), .A2(n_211), .B(n_217), .Y(n_267) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_200), .A2(n_541), .B(n_547), .Y(n_540) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_200), .A2(n_541), .B(n_547), .Y(n_562) );
AO21x2_ASAP7_75t_L g570 ( .A1(n_200), .A2(n_571), .B(n_577), .Y(n_570) );
AO21x2_ASAP7_75t_L g595 ( .A1(n_200), .A2(n_571), .B(n_577), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B1(n_206), .B2(n_207), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g313 ( .A(n_208), .B(n_290), .Y(n_313) );
AND2x2_ASAP7_75t_L g381 ( .A(n_208), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g395 ( .A(n_208), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_208), .B(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2x1_ASAP7_75t_L g258 ( .A(n_210), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g351 ( .A(n_210), .B(n_344), .Y(n_351) );
AND2x2_ASAP7_75t_L g442 ( .A(n_210), .B(n_264), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_218), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_218), .A2(n_499), .B(n_501), .Y(n_498) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_218), .A2(n_581), .B(n_585), .Y(n_580) );
OA21x2_ASAP7_75t_L g625 ( .A1(n_218), .A2(n_581), .B(n_585), .Y(n_625) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g253 ( .A(n_220), .Y(n_253) );
INVx2_ASAP7_75t_L g298 ( .A(n_220), .Y(n_298) );
AND2x2_ASAP7_75t_L g343 ( .A(n_220), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_222), .B(n_228), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_241), .Y(n_231) );
AND2x2_ASAP7_75t_L g385 ( .A(n_232), .B(n_386), .Y(n_385) );
OR2x6_ASAP7_75t_L g444 ( .A(n_232), .B(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
AND2x4_ASAP7_75t_L g282 ( .A(n_233), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g317 ( .A(n_233), .B(n_242), .Y(n_317) );
INVx2_ASAP7_75t_L g366 ( .A(n_233), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_233), .B(n_340), .Y(n_415) );
AND2x2_ASAP7_75t_L g452 ( .A(n_233), .B(n_270), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_233), .B(n_335), .Y(n_460) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x2_ASAP7_75t_L g293 ( .A(n_241), .B(n_282), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_241), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_241), .B(n_320), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_241), .B(n_333), .Y(n_454) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_242), .Y(n_272) );
AND2x2_ASAP7_75t_L g280 ( .A(n_242), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_242), .Y(n_303) );
INVx2_ASAP7_75t_L g306 ( .A(n_242), .Y(n_306) );
INVx1_ASAP7_75t_L g339 ( .A(n_242), .Y(n_339) );
INVx1_ASAP7_75t_L g387 ( .A(n_242), .Y(n_387) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_250), .Y(n_242) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_243), .A2(n_520), .B(n_526), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_253), .B(n_256), .Y(n_329) );
OR2x2_ASAP7_75t_L g401 ( .A(n_253), .B(n_402), .Y(n_401) );
AND4x1_ASAP7_75t_SL g447 ( .A(n_253), .B(n_429), .C(n_448), .D(n_449), .Y(n_447) );
OR2x2_ASAP7_75t_L g471 ( .A(n_254), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g308 ( .A(n_257), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_257), .B(n_266), .Y(n_458) );
AND2x2_ASAP7_75t_L g483 ( .A(n_258), .B(n_343), .Y(n_483) );
OAI32xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_268), .A3(n_273), .B1(n_275), .B2(n_278), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g356 ( .A(n_263), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g456 ( .A(n_263), .B(n_410), .Y(n_456) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x2_ASAP7_75t_L g352 ( .A(n_264), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g438 ( .A(n_264), .Y(n_438) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_265), .B(n_267), .Y(n_472) );
INVx3_ASAP7_75t_L g289 ( .A(n_266), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g467 ( .A(n_266), .B(n_394), .Y(n_467) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_267), .Y(n_326) );
AND2x2_ASAP7_75t_L g345 ( .A(n_267), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g479 ( .A(n_269), .Y(n_479) );
NAND2x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_270), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_273), .B(n_379), .Y(n_378) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g311 ( .A(n_274), .B(n_279), .Y(n_311) );
AND2x4_ASAP7_75t_L g333 ( .A(n_274), .B(n_283), .Y(n_333) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_274), .B(n_405), .Y(n_404) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_274), .B(n_355), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_275), .A2(n_398), .B1(n_401), .B2(n_403), .Y(n_397) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_SL g417 ( .A(n_276), .Y(n_417) );
INVx2_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_280), .B(n_286), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_280), .A2(n_416), .B1(n_419), .B2(n_422), .Y(n_418) );
INVx1_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
AND2x2_ASAP7_75t_L g363 ( .A(n_281), .B(n_322), .Y(n_363) );
INVx2_ASAP7_75t_L g286 ( .A(n_282), .Y(n_286) );
OAI21xp5_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_287), .B(n_291), .Y(n_284) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g359 ( .A1(n_288), .A2(n_360), .B1(n_364), .B2(n_365), .Y(n_359) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_289), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_289), .B(n_357), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_289), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NOR3xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_310), .C(n_314), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_304), .B2(n_307), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g324 ( .A(n_297), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g364 ( .A(n_297), .B(n_351), .Y(n_364) );
AND2x2_ASAP7_75t_L g416 ( .A(n_297), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g433 ( .A(n_297), .B(n_383), .Y(n_433) );
AND2x2_ASAP7_75t_L g488 ( .A(n_297), .B(n_382), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx4_ASAP7_75t_L g355 ( .A(n_300), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_300), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx2_ASAP7_75t_L g370 ( .A(n_303), .Y(n_370) );
AND2x2_ASAP7_75t_L g379 ( .A(n_303), .B(n_363), .Y(n_379) );
INVx1_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_308), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_309), .B(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B(n_323), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_316), .B(n_355), .Y(n_464) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AOI21xp33_ASAP7_75t_SL g327 ( .A1(n_319), .A2(n_328), .B(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g474 ( .A(n_319), .B(n_333), .Y(n_474) );
AND2x4_ASAP7_75t_L g337 ( .A(n_320), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g371 ( .A(n_320), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_320), .B(n_387), .Y(n_453) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B(n_341), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_333), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_333), .B(n_338), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_334), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g396 ( .A(n_334), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_334), .Y(n_400) );
AND2x2_ASAP7_75t_L g484 ( .A(n_334), .B(n_452), .Y(n_484) );
AND2x2_ASAP7_75t_L g487 ( .A(n_334), .B(n_404), .Y(n_487) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_SL g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_339), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g466 ( .A(n_343), .Y(n_466) );
AND2x2_ASAP7_75t_L g357 ( .A(n_344), .B(n_358), .Y(n_357) );
NAND4xp75_ASAP7_75t_L g347 ( .A(n_348), .B(n_367), .C(n_388), .D(n_406), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_359), .Y(n_348) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_351), .B(n_438), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_352), .B(n_417), .Y(n_423) );
NAND2xp5_ASAP7_75t_R g439 ( .A(n_355), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g489 ( .A(n_355), .Y(n_489) );
INVx2_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
BUFx3_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g445 ( .A(n_363), .Y(n_445) );
AND2x2_ASAP7_75t_L g399 ( .A(n_365), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g421 ( .A(n_366), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B(n_374), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_370), .B(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_371), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_373), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_380), .B2(n_384), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OA21x2_ASAP7_75t_L g389 ( .A1(n_382), .A2(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g441 ( .A(n_383), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g449 ( .A(n_383), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_384), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g419 ( .A(n_387), .B(n_420), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_395), .B(n_397), .Y(n_388) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g436 ( .A(n_393), .B(n_437), .Y(n_436) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
INVx2_ASAP7_75t_SL g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_418), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B1(n_413), .B2(n_416), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
NOR2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_461), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_434), .C(n_446), .Y(n_425) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_439), .B1(n_441), .B2(n_443), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_450), .C(n_457), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B(n_455), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_480), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_470), .C(n_477), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_468), .B2(n_469), .Y(n_463) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_471), .B(n_476), .C(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B1(n_485), .B2(n_487), .C1(n_488), .C2(n_489), .Y(n_480) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
XNOR2x1_ASAP7_75t_L g810 ( .A(n_490), .B(n_811), .Y(n_810) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_674), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_629), .C(n_658), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_493), .B(n_602), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_527), .B1(n_548), .B2(n_559), .C(n_563), .Y(n_493) );
INVx3_ASAP7_75t_SL g719 ( .A(n_494), .Y(n_719) );
AND2x2_ASAP7_75t_SL g494 ( .A(n_495), .B(n_506), .Y(n_494) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_495), .B(n_518), .Y(n_565) );
INVx4_ASAP7_75t_L g600 ( .A(n_495), .Y(n_600) );
AND2x2_ASAP7_75t_L g622 ( .A(n_495), .B(n_519), .Y(n_622) );
AND2x2_ASAP7_75t_L g628 ( .A(n_495), .B(n_567), .Y(n_628) );
INVx5_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g597 ( .A(n_496), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_496), .B(n_518), .Y(n_673) );
AND2x2_ASAP7_75t_L g678 ( .A(n_496), .B(n_519), .Y(n_678) );
AND2x2_ASAP7_75t_L g690 ( .A(n_496), .B(n_551), .Y(n_690) );
NOR2x1_ASAP7_75t_SL g729 ( .A(n_496), .B(n_567), .Y(n_729) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
AND2x2_ASAP7_75t_L g662 ( .A(n_506), .B(n_611), .Y(n_662) );
AND2x2_ASAP7_75t_L g759 ( .A(n_506), .B(n_690), .Y(n_759) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g591 ( .A(n_508), .Y(n_591) );
INVx2_ASAP7_75t_L g613 ( .A(n_508), .Y(n_613) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_509), .B(n_517), .Y(n_516) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_509), .A2(n_510), .B(n_516), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
AND2x2_ASAP7_75t_L g588 ( .A(n_518), .B(n_550), .Y(n_588) );
INVx2_ASAP7_75t_L g592 ( .A(n_518), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_518), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g691 ( .A(n_518), .B(n_656), .Y(n_691) );
OR2x2_ASAP7_75t_L g738 ( .A(n_518), .B(n_551), .Y(n_738) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_519), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
AND2x2_ASAP7_75t_L g735 ( .A(n_527), .B(n_616), .Y(n_735) );
AND2x2_ASAP7_75t_L g785 ( .A(n_527), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g661 ( .A(n_528), .B(n_605), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
AND2x2_ASAP7_75t_L g594 ( .A(n_529), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g624 ( .A(n_529), .B(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g645 ( .A(n_529), .B(n_625), .Y(n_645) );
AND2x4_ASAP7_75t_L g680 ( .A(n_529), .B(n_668), .Y(n_680) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g561 ( .A(n_530), .Y(n_561) );
OAI21x1_ASAP7_75t_SL g530 ( .A1(n_531), .A2(n_533), .B(n_537), .Y(n_530) );
INVx1_ASAP7_75t_L g538 ( .A(n_532), .Y(n_538) );
AND2x2_ASAP7_75t_L g607 ( .A(n_539), .B(n_560), .Y(n_607) );
AND2x2_ASAP7_75t_L g693 ( .A(n_539), .B(n_625), .Y(n_693) );
AND2x2_ASAP7_75t_L g704 ( .A(n_539), .B(n_569), .Y(n_704) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g568 ( .A(n_540), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g635 ( .A(n_540), .B(n_570), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_550), .B(n_600), .Y(n_657) );
AND2x2_ASAP7_75t_L g701 ( .A(n_550), .B(n_567), .Y(n_701) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_551), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
BUFx3_ASAP7_75t_L g620 ( .A(n_551), .Y(n_620) );
AND2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_613), .Y(n_643) );
OAI322xp33_ASAP7_75t_L g563 ( .A1(n_558), .A2(n_564), .A3(n_568), .B1(n_578), .B2(n_586), .C1(n_593), .C2(n_598), .Y(n_563) );
INVx1_ASAP7_75t_L g724 ( .A(n_558), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_559), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g637 ( .A(n_559), .B(n_579), .Y(n_637) );
INVx2_ASAP7_75t_L g682 ( .A(n_559), .Y(n_682) );
AND2x2_ASAP7_75t_L g698 ( .A(n_559), .B(n_640), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_559), .B(n_716), .Y(n_746) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_560), .B(n_625), .Y(n_649) );
OR2x2_ASAP7_75t_L g670 ( .A(n_560), .B(n_587), .Y(n_670) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g642 ( .A(n_561), .Y(n_642) );
INVx2_ASAP7_75t_L g587 ( .A(n_562), .Y(n_587) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_562), .Y(n_589) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g632 ( .A(n_565), .Y(n_632) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_566), .Y(n_652) );
INVx1_ASAP7_75t_L g750 ( .A(n_566), .Y(n_750) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_566), .Y(n_765) );
NAND2x1_ASAP7_75t_L g775 ( .A(n_568), .B(n_579), .Y(n_775) );
INVx1_ASAP7_75t_L g782 ( .A(n_568), .Y(n_782) );
BUFx2_ASAP7_75t_L g616 ( .A(n_569), .Y(n_616) );
AND2x2_ASAP7_75t_L g692 ( .A(n_569), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx3_ASAP7_75t_L g601 ( .A(n_570), .Y(n_601) );
INVxp67_ASAP7_75t_L g605 ( .A(n_570), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_578), .B(n_594), .C(n_596), .Y(n_593) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_579), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_579), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g766 ( .A(n_579), .B(n_715), .Y(n_766) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g668 ( .A(n_580), .Y(n_668) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_580), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_586) );
AND2x4_ASAP7_75t_SL g715 ( .A(n_587), .B(n_595), .Y(n_715) );
AND2x2_ASAP7_75t_L g728 ( .A(n_588), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_589), .Y(n_730) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g687 ( .A(n_591), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_591), .B(n_600), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_592), .B(n_610), .Y(n_609) );
AND3x2_ASAP7_75t_L g627 ( .A(n_592), .B(n_620), .C(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g651 ( .A(n_592), .Y(n_651) );
AND2x2_ASAP7_75t_L g764 ( .A(n_592), .B(n_765), .Y(n_764) );
BUFx2_ASAP7_75t_L g640 ( .A(n_595), .Y(n_640) );
INVx1_ASAP7_75t_L g718 ( .A(n_595), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_596), .B(n_619), .Y(n_757) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_597), .B(n_701), .Y(n_706) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g697 ( .A(n_600), .B(n_643), .Y(n_697) );
INVx1_ASAP7_75t_SL g648 ( .A(n_601), .Y(n_648) );
AND2x2_ASAP7_75t_L g756 ( .A(n_601), .B(n_668), .Y(n_756) );
AND2x2_ASAP7_75t_L g777 ( .A(n_601), .B(n_649), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_608), .B1(n_614), .B2(n_617), .C(n_623), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g769 ( .A(n_605), .Y(n_769) );
AOI21xp33_ASAP7_75t_SL g623 ( .A1(n_606), .A2(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_607), .B(n_616), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_607), .A2(n_639), .B1(n_641), .B2(n_646), .C1(n_650), .C2(n_653), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_607), .B(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_608), .A2(n_637), .B1(n_660), .B2(n_662), .Y(n_659) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx1_ASAP7_75t_L g644 ( .A(n_611), .Y(n_644) );
AND2x2_ASAP7_75t_L g763 ( .A(n_611), .B(n_729), .Y(n_763) );
OAI32xp33_ASAP7_75t_L g767 ( .A1(n_611), .A2(n_636), .A3(n_688), .B1(n_696), .B2(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g772 ( .A(n_611), .B(n_622), .Y(n_772) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g656 ( .A(n_613), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g663 ( .A1(n_614), .A2(n_664), .B(n_671), .Y(n_663) );
INVx1_ASAP7_75t_L g727 ( .A(n_616), .Y(n_727) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g631 ( .A(n_619), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g639 ( .A(n_622), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g712 ( .A(n_622), .B(n_643), .Y(n_712) );
INVx1_ASAP7_75t_SL g783 ( .A(n_624), .Y(n_783) );
AND2x2_ASAP7_75t_L g717 ( .A(n_625), .B(n_718), .Y(n_717) );
OAI222xp33_ASAP7_75t_L g770 ( .A1(n_626), .A2(n_679), .B1(n_758), .B2(n_771), .C1(n_773), .C2(n_775), .Y(n_770) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x4_ASAP7_75t_L g743 ( .A(n_628), .B(n_744), .Y(n_743) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_633), .B(n_638), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_632), .B(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g711 ( .A(n_634), .Y(n_711) );
INVx1_ASAP7_75t_L g679 ( .A(n_635), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_635), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g733 ( .A(n_640), .Y(n_733) );
AO22x1_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_645), .Y(n_641) );
OAI322xp33_ASAP7_75t_L g753 ( .A1(n_642), .A2(n_703), .A3(n_706), .B1(n_754), .B2(n_755), .C1(n_757), .C2(n_758), .Y(n_753) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_643), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g672 ( .A(n_644), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_645), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g774 ( .A(n_645), .B(n_704), .Y(n_774) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g754 ( .A(n_648), .Y(n_754) );
INVx1_ASAP7_75t_SL g683 ( .A(n_649), .Y(n_683) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
OR2x2_ASAP7_75t_L g685 ( .A(n_657), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g723 ( .A(n_657), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OR2x2_ASAP7_75t_L g696 ( .A(n_667), .B(n_682), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_667), .B(n_704), .Y(n_703) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g726 ( .A(n_670), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NOR2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_739), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_694), .C(n_707), .D(n_720), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .A3(n_680), .B1(n_681), .B2(n_684), .C1(n_689), .C2(n_692), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g776 ( .A1(n_677), .A2(n_777), .B(n_778), .C(n_781), .Y(n_776) );
AND2x2_ASAP7_75t_L g788 ( .A(n_678), .B(n_765), .Y(n_788) );
INVx1_ASAP7_75t_L g710 ( .A(n_680), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_680), .B(n_715), .Y(n_752) );
NAND2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_688), .B(n_701), .Y(n_768) );
AND2x4_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_698), .B2(n_699), .C1(n_702), .C2(n_705), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_697), .A2(n_708), .B1(n_711), .B2(n_712), .C(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_716), .B(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_725), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g780 ( .A(n_729), .Y(n_780) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B(n_736), .Y(n_731) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx2_ASAP7_75t_L g744 ( .A(n_738), .Y(n_744) );
OR2x2_ASAP7_75t_L g779 ( .A(n_738), .B(n_780), .Y(n_779) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_760), .C(n_776), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_753), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_747), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_766), .B1(n_767), .B2(n_769), .C(n_770), .Y(n_760) );
INVxp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_775), .B(n_779), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B(n_784), .C(n_787), .Y(n_781) );
INVxp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_790), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_791), .A2(n_795), .B1(n_798), .B2(n_801), .Y(n_794) );
INVx3_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVxp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_803), .A2(n_809), .B(n_814), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
BUFx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
BUFx3_ASAP7_75t_L g814 ( .A(n_806), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_815), .Y(n_807) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_821), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
AND2x2_ASAP7_75t_SL g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
endmodule