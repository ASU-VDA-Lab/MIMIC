module fake_jpeg_30666_n_270 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_270);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_45),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_64),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_2),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_39),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_26),
.B1(n_32),
.B2(n_34),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_74),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_24),
.B(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_34),
.B1(n_22),
.B2(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_84),
.B1(n_57),
.B2(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_48),
.B1(n_31),
.B2(n_33),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_37),
.B1(n_32),
.B2(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_31),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_37),
.C(n_43),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_29),
.C(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_91),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_109),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_98),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_60),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_107),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_59),
.B1(n_51),
.B2(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_33),
.B(n_29),
.C(n_25),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_20),
.B1(n_19),
.B2(n_5),
.Y(n_129)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_64),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_52),
.B1(n_31),
.B2(n_37),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_24),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_48),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_122),
.C(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_20),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_3),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_20),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_82),
.C(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_19),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_98),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_162),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_96),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_154),
.C(n_141),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_119),
.C(n_113),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_117),
.B1(n_109),
.B2(n_119),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

OAI22x1_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_103),
.B1(n_109),
.B2(n_126),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_104),
.B1(n_100),
.B2(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_105),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_167),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_126),
.B1(n_82),
.B2(n_81),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_95),
.B1(n_116),
.B2(n_111),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_149),
.B(n_133),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_145),
.B1(n_144),
.B2(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_130),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_177),
.C(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_144),
.B1(n_128),
.B2(n_135),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_144),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_161),
.B(n_134),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_130),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_147),
.B1(n_136),
.B2(n_140),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_182),
.B1(n_176),
.B2(n_180),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_133),
.B(n_138),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_185),
.A2(n_133),
.B(n_165),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_175),
.B1(n_178),
.B2(n_186),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_153),
.C(n_155),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_179),
.C(n_172),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_171),
.B(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_176),
.B1(n_186),
.B2(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_217),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_177),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_210),
.C(n_205),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_195),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_196),
.B1(n_197),
.B2(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_156),
.C(n_146),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_17),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_193),
.B1(n_187),
.B2(n_188),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_124),
.B1(n_127),
.B2(n_121),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_231),
.B1(n_127),
.B2(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_201),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_228),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_192),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_230),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_229),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_146),
.C(n_134),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_138),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_213),
.B(n_215),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_234),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_227),
.A2(n_203),
.B1(n_214),
.B2(n_212),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_231),
.B1(n_225),
.B2(n_219),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_140),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_230),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_16),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_16),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_243),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_248),
.B1(n_14),
.B2(n_10),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_3),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_236),
.C(n_237),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_234),
.B(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_253),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_242),
.C(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_255),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_14),
.C(n_19),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_247),
.C(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_4),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_6),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_255),
.B(n_263),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_260),
.B(n_7),
.Y(n_266)
);

O2A1O1Ixp33_ASAP7_75t_SL g267 ( 
.A1(n_266),
.A2(n_264),
.B(n_7),
.C(n_8),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_6),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_7),
.B(n_9),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_19),
.Y(n_270)
);


endmodule