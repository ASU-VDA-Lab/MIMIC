module real_aes_18336_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_1034;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_1639;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1095;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_1404;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1827;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_1851;
wire n_780;
wire n_931;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1842;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1001 ( .A(n_0), .Y(n_1001) );
INVx1_ASAP7_75t_L g728 ( .A(n_1), .Y(n_728) );
AO22x1_ASAP7_75t_L g754 ( .A1(n_1), .A2(n_236), .B1(n_640), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g373 ( .A(n_2), .Y(n_373) );
AND2x2_ASAP7_75t_L g426 ( .A(n_2), .B(n_263), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_2), .B(n_383), .Y(n_445) );
AND2x2_ASAP7_75t_L g459 ( .A(n_2), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g738 ( .A(n_3), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_3), .A2(n_125), .B1(n_599), .B2(n_635), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g1824 ( .A1(n_4), .A2(n_322), .B1(n_867), .B2(n_1825), .Y(n_1824) );
AOI221xp5_ASAP7_75t_L g1841 ( .A1(n_4), .A2(n_270), .B1(n_644), .B2(n_1019), .C(n_1842), .Y(n_1841) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_5), .A2(n_197), .B1(n_952), .B2(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_5), .A2(n_177), .B1(n_904), .B2(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1351 ( .A(n_6), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_7), .A2(n_219), .B1(n_663), .B2(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1593 ( .A(n_8), .Y(n_1593) );
AOI22xp5_ASAP7_75t_L g1639 ( .A1(n_8), .A2(n_213), .B1(n_1613), .B2(n_1627), .Y(n_1639) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_9), .A2(n_227), .B1(n_877), .B2(n_878), .Y(n_876) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_9), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_10), .A2(n_95), .B1(n_1613), .B2(n_1615), .Y(n_1631) );
AOI22xp33_ASAP7_75t_L g1698 ( .A1(n_11), .A2(n_346), .B1(n_1605), .B2(n_1610), .Y(n_1698) );
INVx2_ASAP7_75t_L g503 ( .A(n_12), .Y(n_503) );
OAI22xp5_ASAP7_75t_SL g1493 ( .A1(n_13), .A2(n_291), .B1(n_1494), .B2(n_1496), .Y(n_1493) );
OAI221xp5_ASAP7_75t_L g1506 ( .A1(n_13), .A2(n_291), .B1(n_914), .B2(n_966), .C(n_1507), .Y(n_1506) );
XNOR2x1_ASAP7_75t_L g1474 ( .A(n_14), .B(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1555 ( .A(n_15), .Y(n_1555) );
OAI222xp33_ASAP7_75t_L g1578 ( .A1(n_15), .A2(n_168), .B1(n_929), .B2(n_965), .C1(n_1579), .C2(n_1583), .Y(n_1578) );
INVx1_ASAP7_75t_L g1397 ( .A(n_16), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_17), .A2(n_315), .B1(n_1196), .B2(n_1197), .Y(n_1201) );
INVx1_ASAP7_75t_L g1225 ( .A(n_17), .Y(n_1225) );
INVx1_ASAP7_75t_L g838 ( .A(n_18), .Y(n_838) );
INVx1_ASAP7_75t_L g1395 ( .A(n_19), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g1411 ( .A1(n_19), .A2(n_69), .B1(n_905), .B2(n_980), .Y(n_1411) );
AOI22xp5_ASAP7_75t_L g1647 ( .A1(n_20), .A2(n_222), .B1(n_1605), .B2(n_1610), .Y(n_1647) );
INVx1_ASAP7_75t_L g1206 ( .A(n_21), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_22), .A2(n_129), .B1(n_950), .B2(n_952), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_22), .A2(n_298), .B1(n_905), .B2(n_980), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_23), .A2(n_316), .B1(n_771), .B2(n_882), .Y(n_1309) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_24), .Y(n_368) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_24), .B(n_366), .Y(n_1606) );
INVx1_ASAP7_75t_L g1505 ( .A(n_25), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1696 ( .A1(n_26), .A2(n_193), .B1(n_1613), .B2(n_1697), .Y(n_1696) );
OAI211xp5_ASAP7_75t_SL g1256 ( .A1(n_27), .A2(n_1257), .B(n_1258), .C(n_1262), .Y(n_1256) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_27), .A2(n_279), .B1(n_663), .B2(n_1066), .Y(n_1267) );
OAI22xp5_ASAP7_75t_SL g796 ( .A1(n_28), .A2(n_299), .B1(n_797), .B2(n_798), .Y(n_796) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_28), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_29), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_30), .A2(n_224), .B1(n_516), .B2(n_1298), .Y(n_1301) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_30), .A2(n_330), .B1(n_975), .B2(n_1325), .C(n_1327), .Y(n_1324) );
INVx1_ASAP7_75t_L g1433 ( .A(n_31), .Y(n_1433) );
OAI211xp5_ASAP7_75t_L g1442 ( .A1(n_31), .A2(n_912), .B(n_1198), .C(n_1443), .Y(n_1442) );
AOI22xp33_ASAP7_75t_L g1636 ( .A1(n_32), .A2(n_210), .B1(n_1613), .B2(n_1615), .Y(n_1636) );
INVxp67_ASAP7_75t_L g1818 ( .A(n_32), .Y(n_1818) );
AOI22xp33_ASAP7_75t_L g1862 ( .A1(n_32), .A2(n_1863), .B1(n_1867), .B2(n_1869), .Y(n_1862) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_33), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_34), .A2(n_53), .B1(n_487), .B2(n_515), .Y(n_594) );
INVx1_ASAP7_75t_L g609 ( .A(n_34), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g1049 ( .A1(n_35), .A2(n_637), .B(n_901), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_35), .A2(n_328), .B1(n_516), .B2(n_693), .Y(n_1073) );
INVx1_ASAP7_75t_L g1294 ( .A(n_36), .Y(n_1294) );
OAI221xp5_ASAP7_75t_L g1318 ( .A1(n_36), .A2(n_255), .B1(n_966), .B2(n_1026), .C(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g464 ( .A(n_37), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_38), .A2(n_51), .B1(n_396), .B2(n_403), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_38), .A2(n_159), .B1(n_514), .B2(n_516), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g1193 ( .A1(n_39), .A2(n_111), .B1(n_902), .B2(n_1054), .C(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1226 ( .A(n_39), .Y(n_1226) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_40), .B(n_853), .Y(n_1244) );
INVx1_ASAP7_75t_L g1576 ( .A(n_41), .Y(n_1576) );
INVx1_ASAP7_75t_L g1064 ( .A(n_42), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1453 ( .A1(n_43), .A2(n_318), .B1(n_635), .B2(n_637), .C(n_971), .Y(n_1453) );
INVxp67_ASAP7_75t_SL g1461 ( .A(n_43), .Y(n_1461) );
INVx1_ASAP7_75t_L g1439 ( .A(n_44), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1454 ( .A1(n_44), .A2(n_214), .B1(n_1257), .B2(n_1455), .Y(n_1454) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_45), .A2(n_353), .B1(n_494), .B2(n_583), .C(n_584), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g607 ( .A1(n_45), .A2(n_118), .B1(n_598), .B2(n_601), .C(n_608), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_46), .Y(n_1093) );
OAI211xp5_ASAP7_75t_SL g1122 ( .A1(n_47), .A2(n_1117), .B(n_1123), .C(n_1126), .Y(n_1122) );
INVx1_ASAP7_75t_L g1172 ( .A(n_47), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_48), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_49), .A2(n_290), .B1(n_672), .B2(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g916 ( .A(n_49), .Y(n_916) );
NAND5xp2_ASAP7_75t_L g625 ( .A(n_50), .B(n_626), .C(n_665), .D(n_689), .E(n_698), .Y(n_625) );
INVx1_ASAP7_75t_L g711 ( .A(n_50), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_51), .A2(n_172), .B1(n_479), .B2(n_486), .Y(n_478) );
INVx1_ASAP7_75t_L g1575 ( .A(n_52), .Y(n_1575) );
INVx1_ASAP7_75t_L g603 ( .A(n_53), .Y(n_603) );
INVxp67_ASAP7_75t_SL g1452 ( .A(n_54), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_54), .A2(n_134), .B1(n_1470), .B2(n_1471), .Y(n_1469) );
AOI22xp5_ASAP7_75t_L g1612 ( .A1(n_55), .A2(n_165), .B1(n_1613), .B2(n_1615), .Y(n_1612) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_56), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_57), .A2(n_58), .B1(n_495), .B2(n_878), .Y(n_1004) );
INVx1_ASAP7_75t_L g1028 ( .A(n_57), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_58), .A2(n_135), .B1(n_902), .B2(n_1017), .C(n_1019), .Y(n_1016) );
INVx1_ASAP7_75t_L g1061 ( .A(n_59), .Y(n_1061) );
OAI22xp33_ASAP7_75t_L g1077 ( .A1(n_59), .A2(n_317), .B1(n_691), .B2(n_957), .Y(n_1077) );
INVx1_ASAP7_75t_L g862 ( .A(n_60), .Y(n_862) );
INVx1_ASAP7_75t_L g1504 ( .A(n_61), .Y(n_1504) );
INVx1_ASAP7_75t_L g1131 ( .A(n_62), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_62), .A2(n_1160), .B(n_1162), .C(n_1164), .Y(n_1159) );
XOR2x2_ASAP7_75t_L g1079 ( .A(n_63), .B(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1211 ( .A(n_64), .Y(n_1211) );
OAI332xp33_ASAP7_75t_SL g1215 ( .A1(n_64), .A2(n_679), .A3(n_840), .B1(n_1216), .B2(n_1222), .B3(n_1223), .C1(n_1229), .C2(n_1233), .Y(n_1215) );
AOI221xp5_ASAP7_75t_L g1259 ( .A1(n_65), .A2(n_113), .B1(n_985), .B2(n_1056), .C(n_1260), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_65), .A2(n_260), .B1(n_880), .B2(n_1012), .Y(n_1275) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_66), .A2(n_169), .B1(n_599), .B2(n_635), .C(n_637), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_66), .A2(n_246), .B1(n_516), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_67), .A2(n_246), .B1(n_633), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_67), .A2(n_169), .B1(n_516), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1828 ( .A1(n_68), .A2(n_156), .B1(n_873), .B2(n_1006), .Y(n_1828) );
AOI21xp33_ASAP7_75t_L g1849 ( .A1(n_68), .A2(n_975), .B(n_1017), .Y(n_1849) );
INVx1_ASAP7_75t_L g1383 ( .A(n_69), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_70), .A2(n_264), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
INVx1_ASAP7_75t_L g1232 ( .A(n_70), .Y(n_1232) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_71), .A2(n_342), .B1(n_407), .B2(n_411), .C(n_415), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_71), .A2(n_302), .B1(n_505), .B2(n_507), .C(n_510), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_72), .A2(n_96), .B1(n_907), .B2(n_980), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_72), .A2(n_244), .B1(n_877), .B2(n_880), .Y(n_1076) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_73), .A2(n_174), .B1(n_505), .B2(n_867), .Y(n_866) );
INVxp67_ASAP7_75t_SL g922 ( .A(n_73), .Y(n_922) );
OAI211xp5_ASAP7_75t_SL g570 ( .A1(n_74), .A2(n_526), .B(n_539), .C(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g614 ( .A(n_74), .Y(n_614) );
INVx1_ASAP7_75t_L g1208 ( .A(n_75), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g1831 ( .A(n_76), .Y(n_1831) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_77), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g1853 ( .A1(n_78), .A2(n_882), .B(n_1854), .Y(n_1853) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_79), .A2(n_241), .B1(n_493), .B2(n_877), .Y(n_1344) );
AOI22xp33_ASAP7_75t_SL g1367 ( .A1(n_79), .A2(n_295), .B1(n_1022), .B2(n_1196), .Y(n_1367) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_80), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_80), .A2(n_349), .B1(n_518), .B2(n_522), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g1302 ( .A1(n_81), .A2(n_356), .B1(n_495), .B2(n_1303), .Y(n_1302) );
AOI221xp5_ASAP7_75t_L g1314 ( .A1(n_81), .A2(n_142), .B1(n_644), .B2(n_804), .C(n_972), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_82), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1827 ( .A1(n_83), .A2(n_270), .B1(n_827), .B2(n_878), .Y(n_1827) );
AOI22xp33_ASAP7_75t_L g1847 ( .A1(n_83), .A2(n_322), .B1(n_1022), .B2(n_1848), .Y(n_1847) );
OR2x2_ASAP7_75t_L g1437 ( .A(n_84), .B(n_853), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_85), .A2(n_211), .B1(n_966), .B2(n_1449), .C(n_1450), .Y(n_1448) );
OAI322xp33_ASAP7_75t_L g1459 ( .A1(n_85), .A2(n_820), .A3(n_958), .B1(n_1399), .B2(n_1460), .C1(n_1462), .C2(n_1466), .Y(n_1459) );
AOI22xp33_ASAP7_75t_SL g1343 ( .A1(n_86), .A2(n_232), .B1(n_486), .B2(n_1341), .Y(n_1343) );
INVx1_ASAP7_75t_L g1364 ( .A(n_86), .Y(n_1364) );
AOI22xp33_ASAP7_75t_SL g1530 ( .A1(n_87), .A2(n_205), .B1(n_516), .B2(n_672), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_87), .A2(n_93), .B1(n_907), .B2(n_1196), .Y(n_1541) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_88), .A2(n_158), .B1(n_755), .B2(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_88), .Y(n_834) );
INVx1_ASAP7_75t_L g1478 ( .A(n_89), .Y(n_1478) );
AOI22xp33_ASAP7_75t_SL g1486 ( .A1(n_90), .A2(n_292), .B1(n_670), .B2(n_836), .Y(n_1486) );
AOI221xp5_ASAP7_75t_L g1500 ( .A1(n_90), .A2(n_94), .B1(n_644), .B2(n_804), .C(n_901), .Y(n_1500) );
INVx1_ASAP7_75t_L g934 ( .A(n_91), .Y(n_934) );
INVx1_ASAP7_75t_L g1480 ( .A(n_92), .Y(n_1480) );
AOI22xp33_ASAP7_75t_SL g1533 ( .A1(n_93), .A2(n_296), .B1(n_516), .B2(n_672), .Y(n_1533) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_94), .A2(n_190), .B1(n_505), .B2(n_1470), .Y(n_1492) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_96), .A2(n_268), .B1(n_688), .B2(n_867), .Y(n_1072) );
AOI22xp33_ASAP7_75t_SL g1565 ( .A1(n_97), .A2(n_335), .B1(n_495), .B2(n_670), .Y(n_1565) );
INVxp67_ASAP7_75t_SL g1570 ( .A(n_97), .Y(n_1570) );
INVx1_ASAP7_75t_L g1394 ( .A(n_98), .Y(n_1394) );
AOI221xp5_ASAP7_75t_L g1405 ( .A1(n_98), .A2(n_234), .B1(n_971), .B2(n_975), .C(n_1019), .Y(n_1405) );
CKINVDCx5p33_ASAP7_75t_R g1526 ( .A(n_99), .Y(n_1526) );
CKINVDCx5p33_ASAP7_75t_R g1839 ( .A(n_100), .Y(n_1839) );
AOI22xp5_ASAP7_75t_L g1621 ( .A1(n_101), .A2(n_220), .B1(n_1605), .B2(n_1610), .Y(n_1621) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_102), .A2(n_647), .B(n_649), .C(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g707 ( .A(n_102), .Y(n_707) );
INVx1_ASAP7_75t_L g999 ( .A(n_103), .Y(n_999) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_103), .A2(n_136), .B1(n_966), .B2(n_1026), .C(n_1027), .Y(n_1025) );
INVx1_ASAP7_75t_L g1451 ( .A(n_104), .Y(n_1451) );
CKINVDCx5p33_ASAP7_75t_R g1834 ( .A(n_105), .Y(n_1834) );
OAI22xp5_ASAP7_75t_L g1850 ( .A1(n_105), .A2(n_122), .B1(n_1851), .B2(n_1852), .Y(n_1850) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_106), .A2(n_243), .B1(n_632), .B2(n_755), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_106), .A2(n_266), .B1(n_493), .B2(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g1250 ( .A(n_107), .Y(n_1250) );
INVx1_ASAP7_75t_L g786 ( .A(n_108), .Y(n_786) );
INVx1_ASAP7_75t_L g1002 ( .A(n_109), .Y(n_1002) );
INVx1_ASAP7_75t_L g366 ( .A(n_110), .Y(n_366) );
INVx1_ASAP7_75t_L g1238 ( .A(n_111), .Y(n_1238) );
INVx1_ASAP7_75t_L g1522 ( .A(n_112), .Y(n_1522) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_113), .A2(n_273), .B1(n_688), .B2(n_1012), .Y(n_1273) );
INVx1_ASAP7_75t_L g1521 ( .A(n_114), .Y(n_1521) );
INVx1_ASAP7_75t_L g1263 ( .A(n_115), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1277 ( .A1(n_115), .A2(n_182), .B1(n_691), .B2(n_840), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1528 ( .A1(n_116), .A2(n_294), .B1(n_880), .B2(n_1470), .C(n_1529), .Y(n_1528) );
AOI221xp5_ASAP7_75t_L g1540 ( .A1(n_116), .A2(n_238), .B1(n_644), .B2(n_1056), .C(n_1514), .Y(n_1540) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_117), .A2(n_183), .B1(n_672), .B2(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g920 ( .A(n_117), .Y(n_920) );
INVx1_ASAP7_75t_L g589 ( .A(n_118), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_119), .A2(n_310), .B1(n_840), .B2(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1413 ( .A(n_119), .Y(n_1413) );
OAI222xp33_ASAP7_75t_L g744 ( .A1(n_120), .A2(n_341), .B1(n_532), .B2(n_536), .C1(n_745), .C2(n_747), .Y(n_744) );
INVx1_ASAP7_75t_L g758 ( .A(n_120), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_121), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g1833 ( .A(n_122), .Y(n_1833) );
INVx1_ASAP7_75t_L g1046 ( .A(n_123), .Y(n_1046) );
OAI211xp5_ASAP7_75t_L g1051 ( .A1(n_124), .A2(n_977), .B(n_1052), .C(n_1060), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_124), .A2(n_276), .B1(n_663), .B2(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g734 ( .A(n_125), .Y(n_734) );
OAI211xp5_ASAP7_75t_L g790 ( .A1(n_126), .A2(n_791), .B(n_792), .C(n_793), .Y(n_790) );
INVxp33_ASAP7_75t_SL g814 ( .A(n_126), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_127), .A2(n_166), .B1(n_545), .B2(n_548), .Y(n_544) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_127), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g1625 ( .A1(n_128), .A2(n_329), .B1(n_1605), .B2(n_1610), .Y(n_1625) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_129), .A2(n_250), .B1(n_971), .B2(n_972), .C(n_975), .Y(n_970) );
INVx1_ASAP7_75t_L g1385 ( .A(n_130), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1408 ( .A1(n_130), .A2(n_288), .B1(n_971), .B2(n_1409), .C(n_1410), .Y(n_1408) );
INVxp67_ASAP7_75t_SL g1048 ( .A(n_131), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g1074 ( .A1(n_131), .A2(n_285), .B1(n_516), .B2(n_888), .Y(n_1074) );
INVx1_ASAP7_75t_L g857 ( .A(n_132), .Y(n_857) );
OAI222xp33_ASAP7_75t_L g911 ( .A1(n_132), .A2(n_209), .B1(n_912), .B2(n_915), .C1(n_921), .C2(n_928), .Y(n_911) );
XOR2x2_ASAP7_75t_L g938 ( .A(n_133), .B(n_939), .Y(n_938) );
AOI22xp5_ASAP7_75t_L g1646 ( .A1(n_133), .A2(n_226), .B1(n_1613), .B2(n_1615), .Y(n_1646) );
AOI221xp5_ASAP7_75t_L g1447 ( .A1(n_134), .A2(n_223), .B1(n_635), .B2(n_804), .C(n_985), .Y(n_1447) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_135), .A2(n_138), .B1(n_880), .B2(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g998 ( .A(n_136), .Y(n_998) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_137), .A2(n_358), .B1(n_545), .B2(n_548), .Y(n_569) );
INVxp33_ASAP7_75t_SL g619 ( .A(n_137), .Y(n_619) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_138), .Y(n_1029) );
INVx1_ASAP7_75t_L g1334 ( .A(n_139), .Y(n_1334) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_139), .A2(n_140), .B1(n_929), .B2(n_965), .C(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1335 ( .A(n_140), .Y(n_1335) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_141), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g1296 ( .A1(n_142), .A2(n_191), .B1(n_493), .B2(n_495), .Y(n_1296) );
AOI22xp5_ASAP7_75t_L g1640 ( .A1(n_143), .A2(n_242), .B1(n_1605), .B2(n_1610), .Y(n_1640) );
OA21x2_ASAP7_75t_L g1476 ( .A1(n_144), .A2(n_853), .B(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g576 ( .A(n_145), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_145), .A2(n_257), .B1(n_598), .B2(n_601), .C(n_602), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g946 ( .A1(n_146), .A2(n_167), .B1(n_880), .B2(n_947), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g981 ( .A1(n_146), .A2(n_192), .B1(n_900), .B2(n_982), .C(n_985), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_147), .A2(n_308), .B1(n_957), .B2(n_958), .Y(n_956) );
INVx1_ASAP7_75t_L g987 ( .A(n_147), .Y(n_987) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_148), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_149), .A2(n_159), .B1(n_403), .B2(n_438), .C(n_440), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_149), .A2(n_342), .B1(n_493), .B2(n_495), .C(n_500), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_150), .A2(n_330), .B1(n_1298), .B2(n_1300), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_150), .A2(n_224), .B1(n_904), .B2(n_1197), .Y(n_1313) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_151), .A2(n_311), .B1(n_1145), .B2(n_1146), .Y(n_1144) );
OAI22xp33_ASAP7_75t_L g1152 ( .A1(n_151), .A2(n_311), .B1(n_1153), .B2(n_1156), .Y(n_1152) );
INVx1_ASAP7_75t_L g886 ( .A(n_152), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g1308 ( .A(n_153), .Y(n_1308) );
AO22x1_ASAP7_75t_L g1822 ( .A1(n_154), .A2(n_199), .B1(n_1006), .B2(n_1007), .Y(n_1822) );
NAND2xp5_ASAP7_75t_L g1846 ( .A(n_154), .B(n_972), .Y(n_1846) );
INVx1_ASAP7_75t_L g697 ( .A(n_155), .Y(n_697) );
AOI22xp33_ASAP7_75t_SL g1843 ( .A1(n_156), .A2(n_199), .B1(n_1197), .B2(n_1844), .Y(n_1843) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_157), .Y(n_961) );
INVx1_ASAP7_75t_L g825 ( .A(n_158), .Y(n_825) );
OA22x2_ASAP7_75t_L g1245 ( .A1(n_160), .A2(n_1246), .B1(n_1278), .B2(n_1279), .Y(n_1245) );
CKINVDCx16_ASAP7_75t_R g1278 ( .A(n_160), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_161), .A2(n_347), .B1(n_771), .B2(n_882), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_162), .A2(n_297), .B1(n_771), .B2(n_882), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_163), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_164), .A2(n_1026), .B(n_1044), .C(n_1047), .Y(n_1043) );
INVx1_ASAP7_75t_L g1070 ( .A(n_164), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_166), .Y(n_455) );
INVxp67_ASAP7_75t_SL g968 ( .A(n_167), .Y(n_968) );
INVx1_ASAP7_75t_L g1554 ( .A(n_168), .Y(n_1554) );
INVx1_ASAP7_75t_L g731 ( .A(n_170), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_170), .A2(n_271), .B1(n_633), .B2(n_640), .Y(n_766) );
INVx1_ASAP7_75t_L g1266 ( .A(n_171), .Y(n_1266) );
INVx1_ASAP7_75t_L g441 ( .A(n_172), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_173), .A2(n_282), .B1(n_1135), .B2(n_1139), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1173 ( .A1(n_173), .A2(n_282), .B1(n_1174), .B2(n_1177), .Y(n_1173) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_174), .A2(n_227), .B1(n_897), .B2(n_900), .C(n_902), .Y(n_896) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_175), .Y(n_794) );
INVx1_ASAP7_75t_L g806 ( .A(n_176), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_177), .A2(n_283), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_SL g1340 ( .A1(n_178), .A2(n_303), .B1(n_486), .B2(n_1341), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_178), .A2(n_232), .B1(n_907), .B2(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1485 ( .A(n_179), .Y(n_1485) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_179), .A2(n_230), .B1(n_982), .B2(n_1205), .C(n_1514), .Y(n_1513) );
OAI211xp5_ASAP7_75t_L g627 ( .A1(n_180), .A2(n_628), .B(n_630), .C(n_645), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_180), .B(n_663), .Y(n_662) );
XNOR2x2_ASAP7_75t_L g1288 ( .A(n_181), .B(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1264 ( .A(n_182), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_183), .A2(n_290), .B1(n_904), .B2(n_905), .Y(n_903) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_184), .A2(n_238), .B1(n_505), .B2(n_1470), .C(n_1532), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_184), .A2(n_294), .B1(n_802), .B2(n_907), .Y(n_1543) );
INVx1_ASAP7_75t_L g944 ( .A(n_185), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_185), .A2(n_325), .B1(n_965), .B2(n_966), .C(n_967), .Y(n_964) );
INVx2_ASAP7_75t_L g1608 ( .A(n_186), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_186), .B(n_1609), .Y(n_1611) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_186), .B(n_307), .Y(n_1616) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_187), .A2(n_352), .B1(n_1300), .B2(n_1562), .Y(n_1561) );
INVx1_ASAP7_75t_L g1581 ( .A(n_187), .Y(n_1581) );
CKINVDCx5p33_ASAP7_75t_R g1458 ( .A(n_188), .Y(n_1458) );
AOI22xp5_ASAP7_75t_L g1604 ( .A1(n_189), .A2(n_281), .B1(n_1605), .B2(n_1610), .Y(n_1604) );
INVx1_ASAP7_75t_L g1512 ( .A(n_190), .Y(n_1512) );
INVxp67_ASAP7_75t_SL g1320 ( .A(n_191), .Y(n_1320) );
AOI22xp33_ASAP7_75t_SL g955 ( .A1(n_192), .A2(n_301), .B1(n_493), .B2(n_827), .Y(n_955) );
XNOR2xp5_ASAP7_75t_L g1040 ( .A(n_193), .B(n_1041), .Y(n_1040) );
XOR2x2_ASAP7_75t_L g1187 ( .A(n_194), .B(n_1188), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g1838 ( .A(n_195), .Y(n_1838) );
OAI22xp33_ASAP7_75t_L g1305 ( .A1(n_196), .A2(n_275), .B1(n_957), .B2(n_958), .Y(n_1305) );
INVx1_ASAP7_75t_L g1316 ( .A(n_196), .Y(n_1316) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_197), .A2(n_283), .B1(n_635), .B2(n_637), .C(n_1031), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1626 ( .A1(n_198), .A2(n_314), .B1(n_1613), .B2(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g774 ( .A(n_200), .Y(n_774) );
INVx1_ASAP7_75t_L g884 ( .A(n_201), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_202), .A2(n_287), .B1(n_632), .B2(n_633), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_202), .A2(n_306), .B1(n_495), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g1592 ( .A(n_203), .Y(n_1592) );
AOI21xp33_ASAP7_75t_L g1253 ( .A1(n_204), .A2(n_1203), .B(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_204), .A2(n_331), .B1(n_516), .B2(n_693), .Y(n_1274) );
AOI221xp5_ASAP7_75t_L g1544 ( .A1(n_205), .A2(n_296), .B1(n_598), .B2(n_975), .C(n_1514), .Y(n_1544) );
INVx1_ASAP7_75t_L g1389 ( .A(n_206), .Y(n_1389) );
OAI211xp5_ASAP7_75t_L g1248 ( .A1(n_207), .A2(n_1026), .B(n_1249), .C(n_1251), .Y(n_1248) );
INVx1_ASAP7_75t_L g1271 ( .A(n_207), .Y(n_1271) );
INVx1_ASAP7_75t_L g1491 ( .A(n_208), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_208), .A2(n_280), .B1(n_633), .B2(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g859 ( .A(n_209), .Y(n_859) );
INVx1_ASAP7_75t_L g1432 ( .A(n_211), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_212), .Y(n_733) );
INVx1_ASAP7_75t_L g1435 ( .A(n_214), .Y(n_1435) );
OAI22xp5_ASAP7_75t_L g1352 ( .A1(n_215), .A2(n_357), .B1(n_957), .B2(n_958), .Y(n_1352) );
INVx1_ASAP7_75t_L g1360 ( .A(n_215), .Y(n_1360) );
INVx1_ASAP7_75t_L g1472 ( .A(n_216), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_217), .Y(n_656) );
INVx1_ASAP7_75t_L g501 ( .A(n_218), .Y(n_501) );
INVx2_ASAP7_75t_L g512 ( .A(n_218), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_218), .B(n_503), .Y(n_521) );
OAI211xp5_ASAP7_75t_L g1406 ( .A1(n_219), .A2(n_977), .B(n_1407), .C(n_1412), .Y(n_1406) );
INVx1_ASAP7_75t_L g742 ( .A(n_221), .Y(n_742) );
NAND2xp33_ASAP7_75t_SL g767 ( .A(n_221), .B(n_599), .Y(n_767) );
INVx1_ASAP7_75t_L g1465 ( .A(n_223), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_225), .A2(n_324), .B1(n_673), .B2(n_870), .Y(n_1564) );
INVx1_ASAP7_75t_L g1580 ( .A(n_225), .Y(n_1580) );
AOI22xp33_ASAP7_75t_SL g1559 ( .A1(n_228), .A2(n_259), .B1(n_495), .B2(n_1560), .Y(n_1559) );
INVxp67_ASAP7_75t_SL g1584 ( .A(n_228), .Y(n_1584) );
XNOR2xp5_ASAP7_75t_L g1868 ( .A(n_229), .B(n_1819), .Y(n_1868) );
INVx1_ASAP7_75t_L g1490 ( .A(n_230), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1630 ( .A1(n_231), .A2(n_321), .B1(n_1605), .B2(n_1610), .Y(n_1630) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_233), .A2(n_312), .B1(n_647), .B2(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g704 ( .A(n_233), .Y(n_704) );
INVx1_ASAP7_75t_L g1391 ( .A(n_234), .Y(n_1391) );
INVx1_ASAP7_75t_L g1446 ( .A(n_235), .Y(n_1446) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_236), .A2(n_500), .B(n_515), .Y(n_743) );
INVx1_ASAP7_75t_L g769 ( .A(n_237), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g1589 ( .A1(n_239), .A2(n_1066), .B(n_1590), .Y(n_1589) );
BUFx3_ASAP7_75t_L g485 ( .A(n_240), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_241), .A2(n_252), .B1(n_601), .B2(n_985), .C(n_1056), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_243), .A2(n_284), .B1(n_493), .B2(n_836), .Y(n_835) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_244), .A2(n_268), .B1(n_902), .B2(n_1054), .C(n_1056), .Y(n_1053) );
INVx1_ASAP7_75t_L g1214 ( .A(n_245), .Y(n_1214) );
INVx1_ASAP7_75t_L g1538 ( .A(n_247), .Y(n_1538) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_248), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_249), .A2(n_253), .B1(n_817), .B2(n_1377), .Y(n_1376) );
OAI221xp5_ASAP7_75t_L g1402 ( .A1(n_249), .A2(n_253), .B1(n_928), .B2(n_1026), .C(n_1403), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_250), .A2(n_298), .B1(n_509), .B2(n_952), .Y(n_953) );
INVx1_ASAP7_75t_L g721 ( .A(n_251), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_251), .B(n_545), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g1339 ( .A1(n_252), .A2(n_295), .B1(n_493), .B2(n_867), .Y(n_1339) );
AOI21xp33_ASAP7_75t_L g809 ( .A1(n_254), .A2(n_601), .B(n_637), .Y(n_809) );
INVx1_ASAP7_75t_L g823 ( .A(n_254), .Y(n_823) );
INVx1_ASAP7_75t_L g1293 ( .A(n_255), .Y(n_1293) );
INVx1_ASAP7_75t_L g1373 ( .A(n_256), .Y(n_1373) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_257), .A2(n_509), .B(n_510), .Y(n_593) );
XOR2x2_ASAP7_75t_L g781 ( .A(n_258), .B(n_782), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g1622 ( .A1(n_258), .A2(n_272), .B1(n_1613), .B2(n_1615), .Y(n_1622) );
AOI21xp33_ASAP7_75t_L g1572 ( .A1(n_259), .A2(n_644), .B(n_901), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_260), .A2(n_273), .B1(n_907), .B2(n_980), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_261), .B(n_1330), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1347 ( .A1(n_261), .A2(n_1348), .B1(n_1349), .B2(n_1368), .Y(n_1347) );
INVx1_ASAP7_75t_L g1370 ( .A(n_261), .Y(n_1370) );
CKINVDCx5p33_ASAP7_75t_R g1086 ( .A(n_262), .Y(n_1086) );
BUFx3_ASAP7_75t_L g383 ( .A(n_263), .Y(n_383) );
INVx1_ASAP7_75t_L g460 ( .A(n_263), .Y(n_460) );
INVx1_ASAP7_75t_L g1219 ( .A(n_264), .Y(n_1219) );
XNOR2x1_ASAP7_75t_L g1518 ( .A(n_265), .B(n_1519), .Y(n_1518) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_266), .B(n_601), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g1261 ( .A1(n_267), .A2(n_331), .B1(n_907), .B2(n_1058), .Y(n_1261) );
AOI22xp33_ASAP7_75t_SL g1276 ( .A1(n_267), .A2(n_340), .B1(n_888), .B2(n_1007), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_269), .Y(n_581) );
INVx1_ASAP7_75t_L g740 ( .A(n_271), .Y(n_740) );
INVx1_ASAP7_75t_L g1537 ( .A(n_274), .Y(n_1537) );
INVx1_ASAP7_75t_L g1317 ( .A(n_275), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g1346 ( .A(n_277), .Y(n_1346) );
INVx1_ASAP7_75t_L g1444 ( .A(n_278), .Y(n_1444) );
NAND2xp33_ASAP7_75t_SL g1487 ( .A(n_280), .B(n_870), .Y(n_1487) );
NAND2xp5_ASAP7_75t_SL g803 ( .A(n_284), .B(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_285), .A2(n_328), .B1(n_907), .B2(n_1058), .Y(n_1057) );
INVx1_ASAP7_75t_L g560 ( .A(n_286), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_287), .A2(n_359), .B1(n_495), .B2(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g1398 ( .A(n_288), .Y(n_1398) );
INVx1_ASAP7_75t_L g483 ( .A(n_289), .Y(n_483) );
INVx1_ASAP7_75t_L g491 ( .A(n_289), .Y(n_491) );
INVx1_ASAP7_75t_L g1509 ( .A(n_292), .Y(n_1509) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_293), .Y(n_994) );
OAI211xp5_ASAP7_75t_L g1014 ( .A1(n_297), .A2(n_977), .B(n_1015), .C(n_1023), .Y(n_1014) );
OAI21xp33_ASAP7_75t_L g812 ( .A1(n_299), .A2(n_691), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g1557 ( .A(n_300), .Y(n_1557) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_301), .Y(n_969) );
INVx1_ASAP7_75t_L g442 ( .A(n_302), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g1365 ( .A1(n_303), .A2(n_975), .B(n_1366), .Y(n_1365) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_304), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g1525 ( .A(n_305), .Y(n_1525) );
AOI221xp5_ASAP7_75t_SL g642 ( .A1(n_306), .A2(n_359), .B1(n_599), .B2(n_643), .C(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g1609 ( .A(n_307), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_307), .B(n_1608), .Y(n_1614) );
INVx1_ASAP7_75t_L g988 ( .A(n_308), .Y(n_988) );
INVx1_ASAP7_75t_L g1209 ( .A(n_309), .Y(n_1209) );
INVx1_ASAP7_75t_L g1414 ( .A(n_310), .Y(n_1414) );
INVx1_ASAP7_75t_L g686 ( .A(n_312), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1637 ( .A1(n_313), .A2(n_350), .B1(n_1605), .B2(n_1610), .Y(n_1637) );
XNOR2xp5_ASAP7_75t_L g561 ( .A(n_314), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1234 ( .A(n_315), .Y(n_1234) );
OAI211xp5_ASAP7_75t_L g1311 ( .A1(n_316), .A2(n_1257), .B(n_1312), .C(n_1315), .Y(n_1311) );
INVx1_ASAP7_75t_L g1062 ( .A(n_317), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g1467 ( .A(n_318), .Y(n_1467) );
INVxp67_ASAP7_75t_SL g1337 ( .A(n_319), .Y(n_1337) );
OAI211xp5_ASAP7_75t_L g1354 ( .A1(n_319), .A2(n_977), .B(n_1355), .C(n_1359), .Y(n_1354) );
CKINVDCx16_ASAP7_75t_R g746 ( .A(n_320), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_323), .Y(n_1103) );
AOI22xp5_ASAP7_75t_L g1573 ( .A1(n_324), .A2(n_352), .B1(n_802), .B2(n_907), .Y(n_1573) );
INVx1_ASAP7_75t_L g943 ( .A(n_325), .Y(n_943) );
OAI21xp33_ASAP7_75t_L g881 ( .A1(n_326), .A2(n_882), .B(n_883), .Y(n_881) );
INVx1_ASAP7_75t_L g564 ( .A(n_327), .Y(n_564) );
OAI21xp5_ASAP7_75t_SL g1545 ( .A1(n_332), .A2(n_1066), .B(n_1546), .Y(n_1545) );
INVx1_ASAP7_75t_L g587 ( .A(n_333), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_334), .Y(n_1088) );
INVxp67_ASAP7_75t_SL g1587 ( .A(n_335), .Y(n_1587) );
CKINVDCx5p33_ASAP7_75t_R g1856 ( .A(n_336), .Y(n_1856) );
OAI211xp5_ASAP7_75t_L g1191 ( .A1(n_337), .A2(n_912), .B(n_1192), .C(n_1198), .Y(n_1191) );
INVx1_ASAP7_75t_L g1241 ( .A(n_337), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_338), .A2(n_355), .B1(n_1056), .B2(n_1203), .C(n_1205), .Y(n_1202) );
INVx1_ASAP7_75t_L g1217 ( .A(n_338), .Y(n_1217) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_339), .Y(n_379) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_340), .Y(n_1252) );
NOR2xp33_ASAP7_75t_R g760 ( .A(n_341), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g716 ( .A(n_343), .Y(n_716) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_344), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_344), .A2(n_345), .B1(n_532), .B2(n_536), .C(n_539), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_345), .A2(n_349), .B1(n_422), .B2(n_430), .C(n_435), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_347), .A2(n_977), .B(n_978), .C(n_986), .Y(n_976) );
XOR2x2_ASAP7_75t_L g991 ( .A(n_348), .B(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g420 ( .A(n_351), .Y(n_420) );
INVx2_ASAP7_75t_L g425 ( .A(n_351), .Y(n_425) );
INVx1_ASAP7_75t_L g450 ( .A(n_351), .Y(n_450) );
INVx1_ASAP7_75t_L g604 ( .A(n_353), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_354), .Y(n_1419) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_355), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g1323 ( .A(n_356), .Y(n_1323) );
INVx1_ASAP7_75t_L g1361 ( .A(n_357), .Y(n_1361) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_358), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_384), .B(n_1596), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_369), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g1861 ( .A(n_363), .B(n_372), .Y(n_1861) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g1866 ( .A(n_365), .B(n_368), .Y(n_1866) );
INVx1_ASAP7_75t_L g1871 ( .A(n_365), .Y(n_1871) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g1873 ( .A(n_368), .B(n_1871), .Y(n_1873) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_372), .B(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g417 ( .A(n_373), .B(n_383), .Y(n_417) );
AND2x4_ASAP7_75t_L g638 ( .A(n_373), .B(n_382), .Y(n_638) );
INVx1_ASAP7_75t_L g1145 ( .A(n_374), .Y(n_1145) );
AND2x4_ASAP7_75t_SL g1860 ( .A(n_374), .B(n_1861), .Y(n_1860) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_376), .B(n_381), .Y(n_375) );
OR2x6_ASAP7_75t_L g1137 ( .A(n_376), .B(n_1138), .Y(n_1137) );
INVxp67_ASAP7_75t_L g1586 ( .A(n_376), .Y(n_1586) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
BUFx4f_ASAP7_75t_L g648 ( .A(n_377), .Y(n_648) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx2_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
INVx2_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
NAND2x1_ASAP7_75t_L g414 ( .A(n_379), .B(n_380), .Y(n_414) );
INVx1_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
AND2x2_ASAP7_75t_L g558 ( .A(n_379), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g600 ( .A(n_379), .B(n_380), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_380), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g409 ( .A(n_380), .B(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g429 ( .A(n_380), .Y(n_429) );
INVx1_ASAP7_75t_L g454 ( .A(n_380), .Y(n_454) );
AND2x2_ASAP7_75t_L g463 ( .A(n_380), .B(n_402), .Y(n_463) );
INVx2_ASAP7_75t_L g559 ( .A(n_380), .Y(n_559) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g1125 ( .A(n_382), .Y(n_1125) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_383), .Y(n_1129) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_383), .B(n_432), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_1035), .B2(n_1595), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AO22x2_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_937), .B1(n_1033), .B2(n_1034), .Y(n_386) );
XOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_621), .Y(n_387) );
XNOR2x1_ASAP7_75t_L g1034 ( .A(n_388), .B(n_621), .Y(n_1034) );
BUFx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
XNOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_561), .Y(n_390) );
XNOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_560), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_476), .Y(n_392) );
NAND3xp33_ASAP7_75t_SL g393 ( .A(n_394), .B(n_446), .C(n_469), .Y(n_393) );
AOI211xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_406), .B(n_421), .C(n_437), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_397), .A2(n_404), .B1(n_1028), .B2(n_1029), .C(n_1030), .Y(n_1027) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_397), .Y(n_1404) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g605 ( .A(n_399), .Y(n_605) );
INVx4_ASAP7_75t_L g798 ( .A(n_399), .Y(n_798) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_399), .Y(n_927) );
INVx2_ASAP7_75t_SL g1322 ( .A(n_399), .Y(n_1322) );
INVx1_ASAP7_75t_L g1511 ( .A(n_399), .Y(n_1511) );
INVx8_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_400), .B(n_1129), .Y(n_1143) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g1319 ( .A1(n_404), .A2(n_1320), .B1(n_1321), .B2(n_1323), .C(n_1324), .Y(n_1319) );
OAI221xp5_ASAP7_75t_SL g1403 ( .A1(n_404), .A2(n_1389), .B1(n_1397), .B2(n_1404), .C(n_1405), .Y(n_1403) );
OAI221xp5_ASAP7_75t_L g1443 ( .A1(n_404), .A2(n_1444), .B1(n_1445), .B2(n_1446), .C(n_1447), .Y(n_1443) );
OAI221xp5_ASAP7_75t_L g1450 ( .A1(n_404), .A2(n_439), .B1(n_1451), .B2(n_1452), .C(n_1453), .Y(n_1450) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_405), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
OAI22x1_ASAP7_75t_SL g608 ( .A1(n_405), .A2(n_581), .B1(n_605), .B2(n_609), .Y(n_608) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_405), .Y(n_1116) );
BUFx3_ASAP7_75t_L g1508 ( .A(n_405), .Y(n_1508) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_408), .A2(n_412), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g1579 ( .A1(n_408), .A2(n_792), .B1(n_1580), .B2(n_1581), .C(n_1582), .Y(n_1579) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g765 ( .A(n_409), .Y(n_765) );
BUFx2_ASAP7_75t_L g797 ( .A(n_409), .Y(n_797) );
BUFx2_ASAP7_75t_L g919 ( .A(n_409), .Y(n_919) );
AND2x2_ASAP7_75t_L g453 ( .A(n_410), .B(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_410), .Y(n_655) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g915 ( .A1(n_412), .A2(n_638), .B1(n_916), .B2(n_917), .C(n_920), .Y(n_915) );
BUFx4f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x6_ASAP7_75t_L g435 ( .A(n_413), .B(n_436), .Y(n_435) );
INVx4_ASAP7_75t_L g650 ( .A(n_413), .Y(n_650) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_413), .Y(n_661) );
BUFx4f_ASAP7_75t_L g1571 ( .A(n_413), .Y(n_1571) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g762 ( .A1(n_415), .A2(n_435), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AND2x4_ASAP7_75t_L g610 ( .A(n_417), .B(n_611), .Y(n_610) );
INVx4_ASAP7_75t_L g644 ( .A(n_417), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g799 ( .A(n_417), .B(n_800), .C(n_801), .D(n_803), .Y(n_799) );
INVx1_ASAP7_75t_SL g902 ( .A(n_417), .Y(n_902) );
INVx4_ASAP7_75t_L g985 ( .A(n_417), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_417), .B(n_611), .Y(n_1120) );
INVx1_ASAP7_75t_L g612 ( .A(n_418), .Y(n_612) );
OR2x2_ASAP7_75t_L g695 ( .A(n_418), .B(n_521), .Y(n_695) );
OR2x2_ASAP7_75t_L g821 ( .A(n_418), .B(n_511), .Y(n_821) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_418), .Y(n_1184) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g434 ( .A(n_419), .Y(n_434) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g615 ( .A(n_422), .Y(n_615) );
INVx2_ASAP7_75t_SL g759 ( .A(n_422), .Y(n_759) );
NAND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_427), .Y(n_422) );
INVx1_ASAP7_75t_L g436 ( .A(n_423), .Y(n_436) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
BUFx2_ASAP7_75t_L g444 ( .A(n_425), .Y(n_444) );
INVx2_ASAP7_75t_L g552 ( .A(n_425), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_426), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_426), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g658 ( .A(n_426), .Y(n_658) );
AND2x6_ASAP7_75t_L g908 ( .A(n_426), .B(n_599), .Y(n_908) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_426), .B(n_652), .Y(n_1045) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g652 ( .A(n_429), .Y(n_652) );
INVx1_ASAP7_75t_L g931 ( .A(n_429), .Y(n_931) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_429), .B(n_1129), .Y(n_1128) );
INVx1_ASAP7_75t_SL g757 ( .A(n_430), .Y(n_757) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
OR2x2_ASAP7_75t_L g617 ( .A(n_431), .B(n_434), .Y(n_617) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g474 ( .A(n_434), .Y(n_474) );
INVxp67_ASAP7_75t_L g664 ( .A(n_434), .Y(n_664) );
INVx1_ASAP7_75t_L g1150 ( .A(n_434), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_435), .Y(n_620) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_443), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_443), .B(n_753), .Y(n_752) );
INVx4_ASAP7_75t_L g1106 ( .A(n_443), .Y(n_1106) );
AND2x4_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OR2x6_ASAP7_75t_L g679 ( .A(n_444), .B(n_500), .Y(n_679) );
INVx1_ASAP7_75t_L g778 ( .A(n_444), .Y(n_778) );
OR2x2_ASAP7_75t_L g1529 ( .A(n_444), .B(n_500), .Y(n_1529) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_455), .B1(n_456), .B2(n_464), .C1(n_465), .C2(n_468), .Y(n_446) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_447), .A2(n_619), .B(n_620), .Y(n_618) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g682 ( .A(n_449), .B(n_529), .Y(n_682) );
OR2x2_ASAP7_75t_L g776 ( .A(n_449), .B(n_452), .Y(n_776) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_450), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g831 ( .A(n_450), .Y(n_831) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g475 ( .A(n_453), .B(n_459), .Y(n_475) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_453), .Y(n_632) );
INVx3_ASAP7_75t_L g641 ( .A(n_453), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_456), .A2(n_572), .B1(n_587), .B2(n_614), .C1(n_615), .C2(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g772 ( .A(n_456), .Y(n_772) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g466 ( .A(n_458), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g761 ( .A(n_458), .B(n_467), .Y(n_761) );
AND2x2_ASAP7_75t_L g556 ( .A(n_459), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g629 ( .A(n_459), .B(n_461), .Y(n_629) );
BUFx2_ASAP7_75t_L g659 ( .A(n_459), .Y(n_659) );
AND2x4_ASAP7_75t_SL g788 ( .A(n_459), .B(n_599), .Y(n_788) );
AND2x4_ASAP7_75t_L g894 ( .A(n_459), .B(n_557), .Y(n_894) );
AND2x4_ASAP7_75t_L g910 ( .A(n_459), .B(n_755), .Y(n_910) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_460), .Y(n_1138) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g1022 ( .A(n_462), .Y(n_1022) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g633 ( .A(n_463), .Y(n_633) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_463), .Y(n_755) );
BUFx3_ASAP7_75t_L g907 ( .A(n_463), .Y(n_907) );
AOI211xp5_ASAP7_75t_L g524 ( .A1(n_464), .A2(n_525), .B(n_531), .C(n_544), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g596 ( .A1(n_465), .A2(n_573), .B1(n_597), .B2(n_606), .C1(n_607), .C2(n_610), .Y(n_596) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g808 ( .A(n_467), .Y(n_808) );
BUFx2_ASAP7_75t_SL g1117 ( .A(n_467), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_472), .B(n_840), .Y(n_839) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_473), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_473), .A2(n_555), .B1(n_720), .B2(n_721), .Y(n_719) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AND2x4_ASAP7_75t_L g555 ( .A(n_474), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g893 ( .A(n_475), .Y(n_893) );
BUFx6f_ASAP7_75t_L g1024 ( .A(n_475), .Y(n_1024) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_524), .B(n_550), .C(n_553), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_492), .B1(n_504), .B2(n_513), .C(n_517), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x6_ASAP7_75t_SL g545 ( .A(n_480), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g693 ( .A(n_480), .Y(n_693) );
BUFx2_ASAP7_75t_L g951 ( .A(n_480), .Y(n_951) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_480), .Y(n_1010) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_481), .Y(n_509) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_481), .Y(n_673) );
BUFx8_ASAP7_75t_L g888 ( .A(n_481), .Y(n_888) );
AND2x4_ASAP7_75t_L g481 ( .A(n_482), .B(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g499 ( .A(n_483), .Y(n_499) );
AND2x4_ASAP7_75t_L g497 ( .A(n_484), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_485), .Y(n_488) );
AND2x4_ASAP7_75t_L g494 ( .A(n_485), .B(n_490), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_485), .B(n_491), .Y(n_580) );
OR2x2_ASAP7_75t_L g727 ( .A(n_485), .B(n_499), .Y(n_727) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx12f_ASAP7_75t_L g516 ( .A(n_487), .Y(n_516) );
AND2x4_ASAP7_75t_L g549 ( .A(n_487), .B(n_547), .Y(n_549) );
INVx5_ASAP7_75t_L g871 ( .A(n_487), .Y(n_871) );
BUFx3_ASAP7_75t_L g952 ( .A(n_487), .Y(n_952) );
BUFx3_ASAP7_75t_L g1007 ( .A(n_487), .Y(n_1007) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g535 ( .A(n_488), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_488), .B(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g1168 ( .A(n_488), .Y(n_1168) );
INVx1_ASAP7_75t_L g538 ( .A(n_489), .Y(n_538) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g506 ( .A(n_494), .Y(n_506) );
AND2x2_ASAP7_75t_L g523 ( .A(n_494), .B(n_520), .Y(n_523) );
BUFx2_ASAP7_75t_L g670 ( .A(n_494), .Y(n_670) );
BUFx2_ASAP7_75t_L g688 ( .A(n_494), .Y(n_688) );
BUFx2_ASAP7_75t_L g880 ( .A(n_494), .Y(n_880) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_494), .B(n_502), .Y(n_1163) );
BUFx2_ASAP7_75t_L g1303 ( .A(n_494), .Y(n_1303) );
INVx8_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_496), .Y(n_583) );
INVx2_ASAP7_75t_L g702 ( .A(n_496), .Y(n_702) );
INVx3_ASAP7_75t_L g877 ( .A(n_496), .Y(n_877) );
INVx2_ASAP7_75t_L g1470 ( .A(n_496), .Y(n_1470) );
INVx8_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx3_ASAP7_75t_L g515 ( .A(n_497), .Y(n_515) );
AND2x2_ASAP7_75t_L g519 ( .A(n_497), .B(n_520), .Y(n_519) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_497), .B(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g827 ( .A(n_497), .Y(n_827) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_497), .Y(n_836) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g585 ( .A(n_500), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
NAND3x1_ASAP7_75t_L g830 ( .A(n_501), .B(n_502), .C(n_831), .Y(n_830) );
AND2x4_ASAP7_75t_L g529 ( .A(n_502), .B(n_530), .Y(n_529) );
OR2x4_ASAP7_75t_L g1155 ( .A(n_502), .B(n_727), .Y(n_1155) );
INVx1_ASAP7_75t_L g1158 ( .A(n_502), .Y(n_1158) );
OR2x6_ASAP7_75t_L g1178 ( .A(n_502), .B(n_1179), .Y(n_1178) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp33_ASAP7_75t_SL g511 ( .A(n_503), .B(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g668 ( .A(n_503), .Y(n_668) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g677 ( .A(n_506), .Y(n_677) );
INVx1_ASAP7_75t_L g1471 ( .A(n_506), .Y(n_1471) );
INVx1_ASAP7_75t_L g1560 ( .A(n_506), .Y(n_1560) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g575 ( .A1(n_508), .A2(n_576), .B1(n_577), .B2(n_581), .C(n_582), .Y(n_575) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_508), .A2(n_540), .B1(n_733), .B2(n_734), .C(n_735), .Y(n_732) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_SL g737 ( .A(n_509), .Y(n_737) );
INVx5_ASAP7_75t_L g833 ( .A(n_509), .Y(n_833) );
INVx2_ASAP7_75t_SL g1342 ( .A(n_509), .Y(n_1342) );
BUFx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g530 ( .A(n_512), .Y(n_530) );
AND3x4_ASAP7_75t_L g667 ( .A(n_512), .B(n_552), .C(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g735 ( .A(n_512), .B(n_668), .Y(n_735) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_512), .Y(n_1182) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g873 ( .A(n_516), .Y(n_873) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_519), .A2(n_523), .B1(n_564), .B2(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g547 ( .A(n_521), .Y(n_547) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x6_ASAP7_75t_L g663 ( .A(n_528), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g771 ( .A(n_528), .B(n_664), .Y(n_771) );
AND2x6_ASAP7_75t_L g533 ( .A(n_529), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g537 ( .A(n_529), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g543 ( .A(n_529), .Y(n_543) );
INVx4_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_533), .A2(n_537), .B1(n_572), .B2(n_573), .Y(n_571) );
AND2x4_ASAP7_75t_SL g681 ( .A(n_534), .B(n_682), .Y(n_681) );
NAND2x1_ASAP7_75t_L g817 ( .A(n_534), .B(n_682), .Y(n_817) );
AND2x2_ASAP7_75t_L g858 ( .A(n_534), .B(n_682), .Y(n_858) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_534), .B(n_682), .Y(n_1495) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g685 ( .A(n_538), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g724 ( .A1(n_539), .A2(n_725), .B1(n_732), .B2(n_736), .C(n_741), .Y(n_724) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
INVx1_ASAP7_75t_L g1237 ( .A(n_540), .Y(n_1237) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
BUFx3_ASAP7_75t_L g1099 ( .A(n_541), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_542), .Y(n_1171) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_547), .Y(n_748) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_549), .B(n_778), .Y(n_777) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_550), .Y(n_811) );
INVx1_ASAP7_75t_L g1417 ( .A(n_550), .Y(n_1417) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI21x1_ASAP7_75t_L g626 ( .A1(n_551), .A2(n_627), .B(n_662), .Y(n_626) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_551), .Y(n_1032) );
BUFx2_ASAP7_75t_L g1588 ( .A(n_551), .Y(n_1588) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI31xp33_ASAP7_75t_SL g568 ( .A1(n_552), .A2(n_569), .A3(n_570), .B(n_574), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_552), .A2(n_723), .A3(n_724), .B(n_744), .Y(n_722) );
INVx2_ASAP7_75t_SL g990 ( .A(n_552), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_555), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g696 ( .A(n_555), .Y(n_696) );
BUFx6f_ASAP7_75t_L g901 ( .A(n_557), .Y(n_901) );
INVx2_ASAP7_75t_L g974 ( .A(n_557), .Y(n_974) );
INVx1_ASAP7_75t_L g1204 ( .A(n_557), .Y(n_1204) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g601 ( .A(n_558), .Y(n_601) );
INVx2_ASAP7_75t_L g636 ( .A(n_558), .Y(n_636) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_558), .B(n_1138), .Y(n_1147) );
AOI211x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_565), .C(n_595), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_586), .C(n_588), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g832 ( .A1(n_577), .A2(n_806), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_577), .A2(n_1230), .B1(n_1231), .B2(n_1232), .Y(n_1229) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_695), .Y(n_706) );
INVx1_ASAP7_75t_L g1221 ( .A(n_578), .Y(n_1221) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_579), .Y(n_730) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
BUFx2_ASAP7_75t_L g1179 ( .A(n_580), .Y(n_1179) );
INVx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_593), .C(n_594), .Y(n_588) );
OAI21xp5_ASAP7_75t_SL g741 ( .A1(n_590), .A2(n_742), .B(n_743), .Y(n_741) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g1089 ( .A(n_591), .Y(n_1089) );
INVx2_ASAP7_75t_L g1384 ( .A(n_591), .Y(n_1384) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g700 ( .A(n_592), .B(n_695), .Y(n_700) );
INVx4_ASAP7_75t_L g1228 ( .A(n_592), .Y(n_1228) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_613), .C(n_618), .Y(n_595) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g804 ( .A(n_599), .Y(n_804) );
BUFx3_ASAP7_75t_L g971 ( .A(n_599), .Y(n_971) );
INVx1_ASAP7_75t_L g1018 ( .A(n_599), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g1056 ( .A(n_599), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_599), .B(n_1125), .Y(n_1124) );
BUFx3_ASAP7_75t_L g1327 ( .A(n_599), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g899 ( .A(n_600), .Y(n_899) );
INVx1_ASAP7_75t_L g1055 ( .A(n_601), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1260 ( .A(n_601), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1583 ( .A1(n_605), .A2(n_1584), .B1(n_1585), .B2(n_1587), .Y(n_1583) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g882 ( .A(n_617), .B(n_700), .Y(n_882) );
AND2x4_ASAP7_75t_L g1066 ( .A(n_617), .B(n_700), .Y(n_1066) );
AO22x2_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_848), .B1(n_935), .B2(n_936), .Y(n_621) );
INVx1_ASAP7_75t_L g935 ( .A(n_622), .Y(n_935) );
XNOR2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_781), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_715), .B1(n_779), .B2(n_780), .Y(n_623) );
INVx1_ASAP7_75t_L g780 ( .A(n_624), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_708), .C(n_712), .Y(n_624) );
INVx1_ASAP7_75t_L g709 ( .A(n_626), .Y(n_709) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_629), .A2(n_894), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_629), .A2(n_908), .B1(n_1480), .B2(n_1500), .C(n_1501), .Y(n_1499) );
AOI221xp5_ASAP7_75t_L g1539 ( .A1(n_629), .A2(n_908), .B1(n_1521), .B2(n_1540), .C(n_1541), .Y(n_1539) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B1(n_639), .B2(n_642), .Y(n_630) );
INVx3_ASAP7_75t_L g1059 ( .A(n_632), .Y(n_1059) );
BUFx6f_ASAP7_75t_L g1358 ( .A(n_632), .Y(n_1358) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g643 ( .A(n_636), .Y(n_643) );
INVx3_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g975 ( .A(n_638), .Y(n_975) );
INVx2_ASAP7_75t_L g1205 ( .A(n_638), .Y(n_1205) );
INVx1_ASAP7_75t_L g1254 ( .A(n_638), .Y(n_1254) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g802 ( .A(n_641), .Y(n_802) );
INVx2_ASAP7_75t_L g904 ( .A(n_641), .Y(n_904) );
INVx1_ASAP7_75t_L g980 ( .A(n_641), .Y(n_980) );
INVx2_ASAP7_75t_L g1196 ( .A(n_641), .Y(n_1196) );
INVx2_ASAP7_75t_SL g1844 ( .A(n_641), .Y(n_1844) );
INVx2_ASAP7_75t_L g1020 ( .A(n_643), .Y(n_1020) );
INVx1_ASAP7_75t_L g1326 ( .A(n_643), .Y(n_1326) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_643), .Y(n_1409) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_645) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_647), .Y(n_1109) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx4_ASAP7_75t_L g791 ( .A(n_648), .Y(n_791) );
BUFx6f_ASAP7_75t_L g924 ( .A(n_648), .Y(n_924) );
OAI211xp5_ASAP7_75t_L g1363 ( .A1(n_649), .A2(n_1364), .B(n_1365), .C(n_1367), .Y(n_1363) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g792 ( .A(n_650), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_656), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_652), .A2(n_654), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_653), .A2(n_681), .B1(n_683), .B2(n_686), .C(n_687), .Y(n_680) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g698 ( .A1(n_656), .A2(n_699), .B1(n_701), .B2(n_704), .C1(n_705), .C2(n_707), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_657), .A2(n_659), .B1(n_790), .B2(n_796), .Y(n_789) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NOR2x1_ASAP7_75t_L g930 ( .A(n_658), .B(n_931), .Y(n_930) );
OAI211xp5_ASAP7_75t_L g1047 ( .A1(n_661), .A2(n_1048), .B(n_1049), .C(n_1050), .Y(n_1047) );
OAI211xp5_ASAP7_75t_L g1251 ( .A1(n_661), .A2(n_1252), .B(n_1253), .C(n_1255), .Y(n_1251) );
INVx5_ASAP7_75t_L g846 ( .A(n_663), .Y(n_846) );
INVx3_ASAP7_75t_L g1436 ( .A(n_663), .Y(n_1436) );
INVx1_ASAP7_75t_L g710 ( .A(n_665), .Y(n_710) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_680), .Y(n_665) );
AOI33xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .A3(n_671), .B1(n_674), .B2(n_676), .B3(n_678), .Y(n_666) );
BUFx3_ASAP7_75t_L g865 ( .A(n_667), .Y(n_865) );
AOI33xp33_ASAP7_75t_L g945 ( .A1(n_667), .A2(n_946), .A3(n_949), .B1(n_953), .B2(n_954), .B3(n_955), .Y(n_945) );
AOI33xp33_ASAP7_75t_L g1071 ( .A1(n_667), .A2(n_1072), .A3(n_1073), .B1(n_1074), .B2(n_1075), .B3(n_1076), .Y(n_1071) );
AOI33xp33_ASAP7_75t_L g1272 ( .A1(n_667), .A2(n_1075), .A3(n_1273), .B1(n_1274), .B2(n_1275), .B3(n_1276), .Y(n_1272) );
AOI33xp33_ASAP7_75t_L g1295 ( .A1(n_667), .A2(n_1296), .A3(n_1297), .B1(n_1301), .B2(n_1302), .B3(n_1304), .Y(n_1295) );
AOI33xp33_ASAP7_75t_L g1338 ( .A1(n_667), .A2(n_954), .A3(n_1339), .B1(n_1340), .B2(n_1343), .B3(n_1344), .Y(n_1338) );
INVx1_ASAP7_75t_L g1532 ( .A(n_667), .Y(n_1532) );
AOI33xp33_ASAP7_75t_L g1558 ( .A1(n_667), .A2(n_1559), .A3(n_1561), .B1(n_1564), .B2(n_1565), .B3(n_1566), .Y(n_1558) );
INVx3_ASAP7_75t_L g1167 ( .A(n_668), .Y(n_1167) );
INVx2_ASAP7_75t_L g1231 ( .A(n_672), .Y(n_1231) );
BUFx6f_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
INVx2_ASAP7_75t_L g1092 ( .A(n_673), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_673), .B(n_1158), .Y(n_1157) );
INVx2_ASAP7_75t_L g1299 ( .A(n_673), .Y(n_1299) );
INVx2_ASAP7_75t_L g1563 ( .A(n_673), .Y(n_1563) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_677), .A2(n_702), .B1(n_720), .B2(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g1075 ( .A(n_679), .Y(n_1075) );
INVx1_ASAP7_75t_L g1566 ( .A(n_679), .Y(n_1566) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_681), .A2(n_683), .B1(n_1046), .B2(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_681), .A2(n_683), .B1(n_1250), .B2(n_1271), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g1524 ( .A1(n_681), .A2(n_683), .B1(n_1525), .B2(n_1526), .Y(n_1524) );
AOI22xp5_ASAP7_75t_L g1553 ( .A1(n_681), .A2(n_683), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
AND2x4_ASAP7_75t_SL g683 ( .A(n_682), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g687 ( .A(n_682), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g818 ( .A(n_682), .B(n_684), .Y(n_818) );
INVx1_ASAP7_75t_L g1496 ( .A(n_683), .Y(n_1496) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g847 ( .A(n_687), .Y(n_847) );
INVx3_ASAP7_75t_L g863 ( .A(n_687), .Y(n_863) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_687), .Y(n_1078) );
NOR3xp33_ASAP7_75t_L g1268 ( .A(n_687), .B(n_1269), .C(n_1277), .Y(n_1268) );
NOR3xp33_ASAP7_75t_SL g1481 ( .A(n_687), .B(n_1482), .C(n_1493), .Y(n_1481) );
BUFx2_ASAP7_75t_L g1825 ( .A(n_688), .Y(n_1825) );
INVx1_ASAP7_75t_L g714 ( .A(n_689), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_697), .Y(n_689) );
NAND2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_696), .Y(n_690) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_692), .A2(n_701), .B1(n_1537), .B2(n_1538), .Y(n_1546) );
AOI22xp33_ASAP7_75t_L g1590 ( .A1(n_692), .A2(n_701), .B1(n_1575), .B2(n_1576), .Y(n_1590) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx2_ASAP7_75t_L g1489 ( .A(n_693), .Y(n_1489) );
INVxp67_ASAP7_75t_L g843 ( .A(n_694), .Y(n_843) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g703 ( .A(n_695), .Y(n_703) );
INVx1_ASAP7_75t_L g713 ( .A(n_698), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_699), .A2(n_705), .B1(n_795), .B2(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_701), .A2(n_887), .B1(n_1001), .B2(n_1002), .Y(n_1000) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AND2x4_ASAP7_75t_L g885 ( .A(n_702), .B(n_703), .Y(n_885) );
AND2x4_ASAP7_75t_L g887 ( .A(n_703), .B(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x4_ASAP7_75t_L g853 ( .A(n_706), .B(n_776), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_711), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g779 ( .A(n_715), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_749), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_722), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_729), .B2(n_731), .Y(n_725) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_726), .Y(n_1087) );
INVx1_ASAP7_75t_L g1464 ( .A(n_726), .Y(n_1464) );
BUFx4f_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g842 ( .A(n_727), .Y(n_842) );
OR2x4_ASAP7_75t_L g1176 ( .A(n_727), .B(n_1158), .Y(n_1176) );
BUFx3_ASAP7_75t_L g1224 ( .A(n_727), .Y(n_1224) );
BUFx3_ASAP7_75t_L g1235 ( .A(n_727), .Y(n_1235) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_729), .A2(n_1087), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx3_ASAP7_75t_L g739 ( .A(n_730), .Y(n_739) );
INVx3_ASAP7_75t_L g824 ( .A(n_730), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g763 ( .A1(n_733), .A2(n_764), .B(n_766), .C(n_767), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g822 ( .A1(n_737), .A2(n_823), .B1(n_824), .B2(n_825), .C(n_826), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g1484 ( .A1(n_737), .A2(n_1485), .B(n_1486), .C(n_1487), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_739), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_739), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
OAI22xp5_ASAP7_75t_L g1392 ( .A1(n_739), .A2(n_1393), .B1(n_1394), .B2(n_1395), .Y(n_1392) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_746), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_756) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_768), .C(n_773), .Y(n_749) );
NOR3xp33_ASAP7_75t_SL g750 ( .A(n_751), .B(n_760), .C(n_762), .Y(n_750) );
OAI21xp5_ASAP7_75t_SL g751 ( .A1(n_752), .A2(n_754), .B(n_756), .Y(n_751) );
BUFx2_ASAP7_75t_L g1197 ( .A(n_755), .Y(n_1197) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
BUFx2_ASAP7_75t_L g933 ( .A(n_778), .Y(n_933) );
INVx1_ASAP7_75t_L g1456 ( .A(n_778), .Y(n_1456) );
AND5x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_815), .C(n_837), .D(n_844), .E(n_847), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_811), .B(n_812), .Y(n_783) );
NAND4xp25_ASAP7_75t_L g784 ( .A(n_785), .B(n_789), .C(n_799), .D(n_805), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
AOI221x1_ASAP7_75t_L g815 ( .A1(n_786), .A2(n_794), .B1(n_816), .B2(n_818), .C(n_819), .Y(n_815) );
AOI222xp33_ASAP7_75t_L g1542 ( .A1(n_787), .A2(n_1045), .B1(n_1525), .B2(n_1526), .C1(n_1543), .C2(n_1544), .Y(n_1542) );
INVx1_ASAP7_75t_L g1851 ( .A(n_787), .Y(n_1851) );
BUFx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g914 ( .A(n_788), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_797), .A2(n_807), .B1(n_1091), .B2(n_1097), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_797), .A2(n_1088), .B1(n_1104), .B2(n_1110), .Y(n_1113) );
INVx2_ASAP7_75t_L g1111 ( .A(n_798), .Y(n_1111) );
OAI211xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .B(n_809), .C(n_810), .Y(n_805) );
INVx5_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_816), .A2(n_818), .B1(n_943), .B2(n_944), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_816), .A2(n_818), .B1(n_998), .B2(n_999), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_816), .A2(n_818), .B1(n_1206), .B2(n_1241), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_816), .A2(n_818), .B1(n_1293), .B2(n_1294), .Y(n_1292) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_816), .A2(n_818), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AO22x1_ASAP7_75t_L g856 ( .A1(n_818), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_818), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_818), .A2(n_858), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
AOI22xp33_ASAP7_75t_L g1832 ( .A1(n_818), .A2(n_858), .B1(n_1833), .B2(n_1834), .Y(n_1832) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_820), .A2(n_822), .B1(n_828), .B2(n_832), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx4f_ASAP7_75t_L g1084 ( .A(n_821), .Y(n_1084) );
BUFx8_ASAP7_75t_L g1222 ( .A(n_821), .Y(n_1222) );
BUFx4f_ASAP7_75t_L g1483 ( .A(n_821), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1460 ( .A1(n_824), .A2(n_1299), .B1(n_1444), .B2(n_1461), .Y(n_1460) );
INVx2_ASAP7_75t_SL g868 ( .A(n_827), .Y(n_868) );
INVx1_ASAP7_75t_L g948 ( .A(n_827), .Y(n_948) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_827), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_828), .A2(n_1483), .B1(n_1484), .B2(n_1488), .Y(n_1482) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx3_ASAP7_75t_L g875 ( .A(n_830), .Y(n_875) );
INVx8_ASAP7_75t_L g1096 ( .A(n_833), .Y(n_1096) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_833), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
OR2x6_ASAP7_75t_L g840 ( .A(n_841), .B(n_843), .Y(n_840) );
OR2x2_ASAP7_75t_L g957 ( .A(n_841), .B(n_843), .Y(n_957) );
INVx2_ASAP7_75t_SL g1388 ( .A(n_841), .Y(n_1388) );
INVx2_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_846), .B(n_862), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_846), .B(n_1209), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_846), .B(n_1337), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1556 ( .A(n_846), .B(n_1557), .Y(n_1556) );
INVx2_ASAP7_75t_SL g959 ( .A(n_847), .Y(n_959) );
NAND4xp75_ASAP7_75t_L g992 ( .A(n_847), .B(n_993), .C(n_996), .D(n_1013), .Y(n_992) );
NAND5xp2_ASAP7_75t_L g1430 ( .A(n_847), .B(n_1431), .C(n_1434), .D(n_1437), .E(n_1438), .Y(n_1430) );
NAND3xp33_ASAP7_75t_SL g1523 ( .A(n_847), .B(n_1524), .C(n_1527), .Y(n_1523) );
INVx2_ASAP7_75t_L g936 ( .A(n_848), .Y(n_936) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_934), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g849 ( .A(n_850), .B(n_889), .Y(n_849) );
AOI211x1_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_852), .B(n_854), .C(n_881), .Y(n_850) );
AOI21xp33_ASAP7_75t_SL g960 ( .A1(n_852), .A2(n_961), .B(n_962), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_852), .A2(n_994), .B(n_995), .Y(n_993) );
AOI21xp33_ASAP7_75t_L g1063 ( .A1(n_852), .A2(n_1064), .B(n_1065), .Y(n_1063) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_852), .A2(n_1266), .B(n_1267), .Y(n_1265) );
AOI21xp33_ASAP7_75t_SL g1307 ( .A1(n_852), .A2(n_1308), .B(n_1309), .Y(n_1307) );
NAND2xp33_ASAP7_75t_L g1345 ( .A(n_852), .B(n_1346), .Y(n_1345) );
AOI21xp33_ASAP7_75t_L g1418 ( .A1(n_852), .A2(n_1419), .B(n_1420), .Y(n_1418) );
AOI221xp5_ASAP7_75t_L g1520 ( .A1(n_852), .A2(n_1436), .B1(n_1521), .B2(n_1522), .C(n_1523), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_852), .B(n_1592), .Y(n_1591) );
NAND2xp5_ASAP7_75t_L g1855 ( .A(n_852), .B(n_1856), .Y(n_1855) );
INVx8_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_864), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_861), .B(n_863), .Y(n_860) );
NAND2xp5_ASAP7_75t_R g909 ( .A(n_862), .B(n_910), .Y(n_909) );
NAND4xp25_ASAP7_75t_L g1239 ( .A(n_863), .B(n_1240), .C(n_1242), .D(n_1243), .Y(n_1239) );
INVx1_ASAP7_75t_L g1306 ( .A(n_863), .Y(n_1306) );
NAND4xp25_ASAP7_75t_SL g1332 ( .A(n_863), .B(n_1333), .C(n_1336), .D(n_1338), .Y(n_1332) );
AND4x1_ASAP7_75t_L g1552 ( .A(n_863), .B(n_1553), .C(n_1556), .D(n_1558), .Y(n_1552) );
NAND3xp33_ASAP7_75t_L g1829 ( .A(n_863), .B(n_1830), .C(n_1832), .Y(n_1829) );
AOI33xp33_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_866), .A3(n_869), .B1(n_872), .B2(n_874), .B3(n_876), .Y(n_864) );
AOI33xp33_ASAP7_75t_L g1003 ( .A1(n_865), .A2(n_954), .A3(n_1004), .B1(n_1005), .B2(n_1008), .B3(n_1011), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_865), .B(n_1824), .Y(n_1823) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_R g1300 ( .A(n_871), .Y(n_1300) );
BUFx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx2_ASAP7_75t_L g954 ( .A(n_875), .Y(n_954) );
BUFx2_ASAP7_75t_L g1304 ( .A(n_875), .Y(n_1304) );
BUFx2_ASAP7_75t_L g1400 ( .A(n_875), .Y(n_1400) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g1213 ( .A(n_882), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1421 ( .A(n_882), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_884), .A2(n_886), .B1(n_892), .B2(n_894), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_885), .B(n_1439), .Y(n_1438) );
AOI22xp5_ASAP7_75t_L g1516 ( .A1(n_885), .A2(n_1504), .B1(n_1505), .B2(n_1517), .Y(n_1516) );
AOI22xp33_ASAP7_75t_L g1854 ( .A1(n_885), .A2(n_887), .B1(n_1838), .B2(n_1839), .Y(n_1854) );
INVx2_ASAP7_75t_L g958 ( .A(n_887), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_887), .B(n_1208), .Y(n_1243) );
INVx2_ASAP7_75t_L g1380 ( .A(n_887), .Y(n_1380) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_888), .Y(n_1006) );
INVx3_ASAP7_75t_L g1218 ( .A(n_888), .Y(n_1218) );
INVx2_ASAP7_75t_SL g1393 ( .A(n_888), .Y(n_1393) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_911), .B(n_932), .Y(n_889) );
NAND3xp33_ASAP7_75t_SL g890 ( .A(n_891), .B(n_895), .C(n_909), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_892), .A2(n_987), .B1(n_988), .B2(n_989), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1262 ( .A1(n_892), .A2(n_989), .B1(n_1263), .B2(n_1264), .Y(n_1262) );
AOI22xp5_ASAP7_75t_L g1315 ( .A1(n_892), .A2(n_989), .B1(n_1316), .B2(n_1317), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_892), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
BUFx6f_ASAP7_75t_L g989 ( .A(n_894), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_894), .A2(n_1001), .B1(n_1002), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_894), .A2(n_1024), .B1(n_1360), .B2(n_1361), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1415 ( .A(n_894), .Y(n_1415) );
AOI22xp5_ASAP7_75t_L g1503 ( .A1(n_894), .A2(n_1024), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
AOI22xp5_ASAP7_75t_L g1536 ( .A1(n_894), .A2(n_1024), .B1(n_1537), .B2(n_1538), .Y(n_1536) );
AOI22xp5_ASAP7_75t_L g1574 ( .A1(n_894), .A2(n_1024), .B1(n_1575), .B2(n_1576), .Y(n_1574) );
AOI22xp33_ASAP7_75t_L g1837 ( .A1(n_894), .A2(n_1024), .B1(n_1838), .B2(n_1839), .Y(n_1837) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_903), .B(n_908), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g1842 ( .A(n_898), .Y(n_1842) );
BUFx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g984 ( .A(n_899), .Y(n_984) );
BUFx3_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_908), .A2(n_979), .B(n_981), .Y(n_978) );
AOI21xp5_ASAP7_75t_SL g1015 ( .A1(n_908), .A2(n_1016), .B(n_1021), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g1052 ( .A1(n_908), .A2(n_1053), .B(n_1057), .Y(n_1052) );
INVx1_ASAP7_75t_L g1198 ( .A(n_908), .Y(n_1198) );
AOI21xp5_ASAP7_75t_L g1258 ( .A1(n_908), .A2(n_1259), .B(n_1261), .Y(n_1258) );
AOI21xp5_ASAP7_75t_L g1312 ( .A1(n_908), .A2(n_1313), .B(n_1314), .Y(n_1312) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_908), .A2(n_1356), .B(n_1357), .Y(n_1355) );
AOI21xp5_ASAP7_75t_L g1407 ( .A1(n_908), .A2(n_1408), .B(n_1411), .Y(n_1407) );
AOI221xp5_ASAP7_75t_SL g1840 ( .A1(n_908), .A2(n_910), .B1(n_1831), .B2(n_1841), .C(n_1843), .Y(n_1840) );
INVx2_ASAP7_75t_SL g977 ( .A(n_910), .Y(n_977) );
INVx3_ASAP7_75t_L g1257 ( .A(n_910), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_910), .B(n_1557), .Y(n_1577) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g965 ( .A(n_913), .Y(n_965) );
INVx2_ASAP7_75t_L g1026 ( .A(n_913), .Y(n_1026) );
INVx4_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx4_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_925), .B2(n_926), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g967 ( .A1(n_923), .A2(n_926), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_967) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx5_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
BUFx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g966 ( .A(n_930), .Y(n_966) );
OAI21xp5_ASAP7_75t_SL g1042 ( .A1(n_932), .A2(n_1043), .B(n_1051), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1190 ( .A1(n_932), .A2(n_1191), .B(n_1199), .Y(n_1190) );
OAI21xp5_ASAP7_75t_SL g1247 ( .A1(n_932), .A2(n_1248), .B(n_1256), .Y(n_1247) );
OAI21xp5_ASAP7_75t_L g1353 ( .A1(n_932), .A2(n_1354), .B(n_1362), .Y(n_1353) );
AOI21xp5_ASAP7_75t_L g1534 ( .A1(n_932), .A2(n_1535), .B(n_1545), .Y(n_1534) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1515 ( .A(n_933), .Y(n_1515) );
INVx1_ASAP7_75t_L g1033 ( .A(n_937), .Y(n_1033) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_991), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_940), .B(n_960), .C(n_963), .Y(n_939) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_956), .C(n_959), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_945), .Y(n_941) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g1101 ( .A(n_954), .Y(n_1101) );
INVxp67_ASAP7_75t_L g1517 ( .A(n_958), .Y(n_1517) );
NOR4xp25_ASAP7_75t_L g1375 ( .A(n_959), .B(n_1376), .C(n_1379), .D(n_1381), .Y(n_1375) );
OAI21xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_976), .B(n_990), .Y(n_963) );
BUFx2_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx2_ASAP7_75t_L g1514 ( .A(n_974), .Y(n_1514) );
INVx1_ASAP7_75t_L g1582 ( .A(n_975), .Y(n_1582) );
INVx2_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
HB1xp67_ASAP7_75t_SL g1410 ( .A(n_985), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_989), .A2(n_1024), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1449 ( .A(n_989), .Y(n_1449) );
OAI21xp5_ASAP7_75t_L g1310 ( .A1(n_990), .A2(n_1311), .B(n_1318), .Y(n_1310) );
AOI21xp5_ASAP7_75t_SL g1835 ( .A1(n_990), .A2(n_1836), .B(n_1853), .Y(n_1835) );
AND3x1_ASAP7_75t_L g996 ( .A(n_997), .B(n_1000), .C(n_1003), .Y(n_996) );
INVx2_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
OAI21xp5_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1025), .B(n_1032), .Y(n_1013) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1018), .Y(n_1031) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1018), .Y(n_1194) );
INVx2_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1024), .B(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1024), .Y(n_1455) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1035), .Y(n_1595) );
XNOR2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1424), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1283), .B1(n_1284), .B2(n_1423), .Y(n_1036) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1037), .Y(n_1423) );
AO22x2_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1185), .B1(n_1281), .B2(n_1282), .Y(n_1037) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1038), .Y(n_1281) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1079), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1063), .C(n_1067), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1046), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_1045), .A2(n_1201), .B1(n_1202), .B2(n_1206), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1045), .B(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1045), .Y(n_1852) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1055), .Y(n_1366) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1059), .Y(n_1502) );
INVx2_ASAP7_75t_SL g1848 ( .A(n_1059), .Y(n_1848) );
INVx1_ASAP7_75t_SL g1479 ( .A(n_1066), .Y(n_1479) );
NOR3xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1077), .C(n_1078), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1071), .Y(n_1068) );
NAND3xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1121), .C(n_1151), .Y(n_1080) );
NOR2xp33_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1105), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1085), .A3(n_1090), .B1(n_1094), .B2(n_1101), .B3(n_1102), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1087), .B1(n_1088), .B2(n_1089), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1086), .A2(n_1103), .B1(n_1108), .B2(n_1110), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_1093), .A2(n_1100), .B1(n_1115), .B2(n_1117), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1097), .B1(n_1098), .B2(n_1100), .Y(n_1094) );
INVx2_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
BUFx6f_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1099), .Y(n_1161) );
OAI33xp33_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .A3(n_1112), .B1(n_1113), .B2(n_1114), .B3(n_1118), .Y(n_1105) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
OAI31xp33_ASAP7_75t_SL g1121 ( .A1(n_1122), .A2(n_1134), .A3(n_1144), .B(n_1148), .Y(n_1121) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_1127), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1126) );
BUFx3_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_1130), .A2(n_1165), .B1(n_1169), .B2(n_1172), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx3_ASAP7_75t_SL g1146 ( .A(n_1147), .Y(n_1146) );
BUFx3_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI31xp33_ASAP7_75t_SL g1151 ( .A1(n_1152), .A2(n_1159), .A3(n_1173), .B(n_1180), .Y(n_1151) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
CKINVDCx8_ASAP7_75t_R g1162 ( .A(n_1163), .Y(n_1162) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1167), .B(n_1171), .Y(n_1170) );
BUFx6f_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_SL g1175 ( .A(n_1176), .Y(n_1175) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
BUFx3_ASAP7_75t_L g1468 ( .A(n_1179), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1183), .Y(n_1180) );
INVx1_ASAP7_75t_SL g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1185), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_1186), .A2(n_1187), .B1(n_1245), .B2(n_1280), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
NOR3xp33_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1239), .C(n_1244), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1212), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1195), .Y(n_1192) );
NAND4xp25_ASAP7_75t_L g1568 ( .A(n_1198), .B(n_1569), .C(n_1574), .D(n_1577), .Y(n_1568) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1207), .C(n_1210), .Y(n_1199) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1204), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1214), .B(n_1215), .Y(n_1212) );
AOI21xp5_ASAP7_75t_L g1350 ( .A1(n_1213), .A2(n_1351), .B(n_1352), .Y(n_1350) );
AOI21xp5_ASAP7_75t_SL g1457 ( .A1(n_1213), .A2(n_1458), .B(n_1459), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_1217), .A2(n_1218), .B1(n_1219), .B2(n_1220), .Y(n_1216) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
OAI33xp33_ASAP7_75t_L g1381 ( .A1(n_1222), .A2(n_1382), .A3(n_1386), .B1(n_1392), .B2(n_1396), .B3(n_1399), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B1(n_1226), .B2(n_1227), .Y(n_1223) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_1234), .A2(n_1235), .B1(n_1236), .B2(n_1238), .Y(n_1233) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1245), .Y(n_1280) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1246), .Y(n_1279) );
NAND3xp33_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1265), .C(n_1268), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1272), .Y(n_1269) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
AO22x2_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1286), .B1(n_1372), .B2(n_1422), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1288), .B1(n_1328), .B2(n_1371), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1307), .C(n_1310), .Y(n_1289) );
NOR3xp33_ASAP7_75t_L g1290 ( .A(n_1291), .B(n_1305), .C(n_1306), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1295), .Y(n_1291) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
HB1xp67_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
HB1xp67_ASAP7_75t_L g1445 ( .A(n_1322), .Y(n_1445) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1328), .Y(n_1371) );
NAND2x1p5_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1347), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1345), .Y(n_1330) );
INVxp67_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NOR2xp33_ASAP7_75t_SL g1368 ( .A(n_1332), .B(n_1369), .Y(n_1368) );
INVx2_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1345), .B(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1353), .Y(n_1349) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1372), .Y(n_1422) );
XNOR2xp5_ASAP7_75t_SL g1372 ( .A(n_1373), .B(n_1374), .Y(n_1372) );
AND3x2_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1401), .C(n_1418), .Y(n_1374) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_1384), .A2(n_1387), .B1(n_1397), .B2(n_1398), .Y(n_1396) );
OAI22xp33_ASAP7_75t_L g1462 ( .A1(n_1384), .A2(n_1451), .B1(n_1463), .B2(n_1465), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1389), .B1(n_1390), .B2(n_1391), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
OAI221xp5_ASAP7_75t_L g1466 ( .A1(n_1390), .A2(n_1446), .B1(n_1467), .B2(n_1468), .C(n_1469), .Y(n_1466) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
NAND3xp33_ASAP7_75t_L g1826 ( .A(n_1400), .B(n_1827), .C(n_1828), .Y(n_1826) );
OAI21xp5_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1406), .B(n_1416), .Y(n_1401) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
OAI22xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1548), .B1(n_1549), .B2(n_1594), .Y(n_1424) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1425), .Y(n_1594) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1428), .B1(n_1473), .B2(n_1547), .Y(n_1426) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
XNOR2x1_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1472), .Y(n_1428) );
NOR2x1_ASAP7_75t_L g1429 ( .A(n_1430), .B(n_1440), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1436), .Y(n_1434) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_1436), .A2(n_1478), .B1(n_1479), .B2(n_1480), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_1436), .B(n_1831), .Y(n_1830) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1457), .Y(n_1440) );
OAI31xp33_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1448), .A3(n_1454), .B(n_1456), .Y(n_1441) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OAI221xp5_ASAP7_75t_L g1488 ( .A1(n_1468), .A2(n_1489), .B1(n_1490), .B2(n_1491), .C(n_1492), .Y(n_1488) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1473), .Y(n_1547) );
XNOR2x1_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1518), .Y(n_1473) );
NAND4xp75_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1481), .C(n_1497), .D(n_1516), .Y(n_1475) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
OAI21xp5_ASAP7_75t_L g1497 ( .A1(n_1498), .A2(n_1506), .B(n_1515), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1499), .B(n_1503), .Y(n_1498) );
OAI221xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1509), .B1(n_1510), .B2(n_1512), .C(n_1513), .Y(n_1507) );
BUFx3_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1534), .Y(n_1519) );
AOI22xp5_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1530), .B1(n_1531), .B2(n_1533), .Y(n_1527) );
NAND3xp33_ASAP7_75t_L g1535 ( .A(n_1536), .B(n_1539), .C(n_1542), .Y(n_1535) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
HB1xp67_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
XOR2xp5_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1593), .Y(n_1550) );
NAND3xp33_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1567), .C(n_1591), .Y(n_1551) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
O2A1O1Ixp5_ASAP7_75t_SL g1567 ( .A1(n_1568), .A2(n_1578), .B(n_1588), .C(n_1589), .Y(n_1567) );
OAI211xp5_ASAP7_75t_L g1569 ( .A1(n_1570), .A2(n_1571), .B(n_1572), .C(n_1573), .Y(n_1569) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
OAI221xp5_ASAP7_75t_SL g1596 ( .A1(n_1597), .A2(n_1813), .B1(n_1816), .B2(n_1857), .C(n_1862), .Y(n_1596) );
AND5x1_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1746), .C(n_1761), .D(n_1790), .E(n_1798), .Y(n_1597) );
AOI21xp5_ASAP7_75t_L g1598 ( .A1(n_1599), .A2(n_1695), .B(n_1699), .Y(n_1598) );
NAND5xp2_ASAP7_75t_L g1599 ( .A(n_1600), .B(n_1650), .C(n_1665), .D(n_1678), .E(n_1693), .Y(n_1599) );
AOI21xp5_ASAP7_75t_L g1600 ( .A1(n_1601), .A2(n_1632), .B(n_1641), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1602), .B(n_1617), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1602), .B(n_1619), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1602), .B(n_1635), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1602), .B(n_1667), .Y(n_1694) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_1602), .B(n_1724), .Y(n_1723) );
CKINVDCx14_ASAP7_75t_R g1755 ( .A(n_1602), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1602), .B(n_1673), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1602), .B(n_1676), .Y(n_1789) );
NOR2xp33_ASAP7_75t_L g1805 ( .A(n_1602), .B(n_1672), .Y(n_1805) );
INVx3_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1655 ( .A(n_1603), .B(n_1656), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_1603), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1603), .B(n_1663), .Y(n_1670) );
AOI311xp33_ASAP7_75t_L g1678 ( .A1(n_1603), .A2(n_1679), .A3(n_1681), .B(n_1683), .C(n_1687), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1603), .B(n_1620), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1603), .B(n_1731), .Y(n_1730) );
OR2x2_ASAP7_75t_L g1744 ( .A(n_1603), .B(n_1733), .Y(n_1744) );
AND2x4_ASAP7_75t_SL g1603 ( .A(n_1604), .B(n_1612), .Y(n_1603) );
AND2x4_ASAP7_75t_L g1605 ( .A(n_1606), .B(n_1607), .Y(n_1605) );
AND2x6_ASAP7_75t_L g1610 ( .A(n_1606), .B(n_1611), .Y(n_1610) );
AND2x6_ASAP7_75t_L g1613 ( .A(n_1606), .B(n_1614), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1606), .B(n_1616), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1606), .B(n_1616), .Y(n_1627) );
AND2x2_ASAP7_75t_L g1697 ( .A(n_1606), .B(n_1616), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1608), .B(n_1609), .Y(n_1607) );
INVx2_ASAP7_75t_L g1815 ( .A(n_1613), .Y(n_1815) );
OAI21xp5_ASAP7_75t_L g1870 ( .A1(n_1614), .A2(n_1871), .B(n_1872), .Y(n_1870) );
A2O1A1Ixp33_ASAP7_75t_L g1746 ( .A1(n_1617), .A2(n_1721), .B(n_1747), .C(n_1758), .Y(n_1746) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
NOR2xp33_ASAP7_75t_L g1778 ( .A(n_1618), .B(n_1779), .Y(n_1778) );
NOR2xp33_ASAP7_75t_L g1797 ( .A(n_1618), .B(n_1708), .Y(n_1797) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1623), .Y(n_1618) );
NAND2xp5_ASAP7_75t_L g1711 ( .A(n_1619), .B(n_1663), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1714 ( .A(n_1619), .B(n_1629), .Y(n_1714) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1619), .B(n_1624), .Y(n_1720) );
NOR2xp33_ASAP7_75t_L g1728 ( .A(n_1619), .B(n_1729), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1738 ( .A(n_1619), .B(n_1676), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1619), .B(n_1691), .Y(n_1756) );
OR2x2_ASAP7_75t_L g1765 ( .A(n_1619), .B(n_1657), .Y(n_1765) );
OR2x2_ASAP7_75t_L g1800 ( .A(n_1619), .B(n_1789), .Y(n_1800) );
INVx2_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1620), .B(n_1661), .Y(n_1660) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1620), .B(n_1629), .Y(n_1682) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1620), .B(n_1664), .Y(n_1685) );
OR2x2_ASAP7_75t_L g1733 ( .A(n_1620), .B(n_1624), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1734 ( .A(n_1620), .B(n_1624), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1620), .B(n_1663), .Y(n_1771) );
OR2x2_ASAP7_75t_L g1777 ( .A(n_1620), .B(n_1670), .Y(n_1777) );
OR2x2_ASAP7_75t_L g1786 ( .A(n_1620), .B(n_1657), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1622), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1641 ( .A(n_1623), .B(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1623), .Y(n_1691) );
OR2x2_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1628), .Y(n_1623) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1624), .Y(n_1658) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1624), .B(n_1629), .Y(n_1676) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1629), .B(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1629), .Y(n_1664) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1629), .Y(n_1808) );
NAND2x1_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1631), .Y(n_1629) );
AOI322xp5_ASAP7_75t_L g1726 ( .A1(n_1632), .A2(n_1694), .A3(n_1701), .B1(n_1727), .B2(n_1728), .C1(n_1732), .C2(n_1736), .Y(n_1726) );
OAI21xp33_ASAP7_75t_L g1787 ( .A1(n_1632), .A2(n_1785), .B(n_1788), .Y(n_1787) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1653 ( .A(n_1633), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1633 ( .A(n_1634), .B(n_1638), .Y(n_1633) );
INVx2_ASAP7_75t_L g1680 ( .A(n_1634), .Y(n_1680) );
AOI321xp33_ASAP7_75t_L g1737 ( .A1(n_1634), .A2(n_1718), .A3(n_1738), .B1(n_1739), .B2(n_1741), .C(n_1743), .Y(n_1737) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1648 ( .A(n_1635), .B(n_1649), .Y(n_1648) );
OR2x2_ASAP7_75t_L g1668 ( .A(n_1635), .B(n_1638), .Y(n_1668) );
INVx2_ASAP7_75t_SL g1673 ( .A(n_1635), .Y(n_1673) );
NAND2xp5_ASAP7_75t_L g1772 ( .A(n_1635), .B(n_1707), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1636), .B(n_1637), .Y(n_1635) );
CKINVDCx5p33_ASAP7_75t_R g1649 ( .A(n_1638), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1659 ( .A(n_1638), .B(n_1644), .Y(n_1659) );
HB1xp67_ASAP7_75t_SL g1757 ( .A(n_1638), .Y(n_1757) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1638), .B(n_1645), .Y(n_1794) );
AND2x4_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1640), .Y(n_1638) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1642), .Y(n_1715) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1648), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1643), .B(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1652 ( .A(n_1644), .B(n_1653), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1644), .B(n_1667), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1644), .B(n_1680), .Y(n_1679) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1644), .Y(n_1731) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1644), .B(n_1695), .Y(n_1740) );
NAND3xp33_ASAP7_75t_L g1812 ( .A(n_1644), .B(n_1656), .C(n_1780), .Y(n_1812) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1645), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1718 ( .A(n_1645), .B(n_1649), .Y(n_1718) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1645), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1645 ( .A(n_1646), .B(n_1647), .Y(n_1645) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1648), .Y(n_1760) );
OR2x2_ASAP7_75t_L g1672 ( .A(n_1649), .B(n_1673), .Y(n_1672) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1649), .B(n_1735), .Y(n_1736) );
OAI32xp33_ASAP7_75t_L g1766 ( .A1(n_1649), .A2(n_1661), .A3(n_1710), .B1(n_1722), .B2(n_1767), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1767 ( .A(n_1649), .B(n_1695), .Y(n_1767) );
NAND2xp5_ASAP7_75t_L g1781 ( .A(n_1649), .B(n_1722), .Y(n_1781) );
AOI211xp5_ASAP7_75t_L g1782 ( .A1(n_1649), .A2(n_1680), .B(n_1695), .C(n_1783), .Y(n_1782) );
AOI22xp33_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1654), .B1(n_1659), .B2(n_1660), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
OAI311xp33_ASAP7_75t_L g1716 ( .A1(n_1655), .A2(n_1695), .A3(n_1717), .B1(n_1719), .C1(n_1725), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1656), .B(n_1703), .Y(n_1702) );
OAI211xp5_ASAP7_75t_L g1719 ( .A1(n_1656), .A2(n_1720), .B(n_1721), .C(n_1723), .Y(n_1719) );
NOR2xp33_ASAP7_75t_L g1727 ( .A(n_1656), .B(n_1691), .Y(n_1727) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1658), .B(n_1664), .Y(n_1663) );
NAND3xp33_ASAP7_75t_L g1725 ( .A(n_1659), .B(n_1680), .C(n_1690), .Y(n_1725) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1659), .Y(n_1745) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1660), .Y(n_1759) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1662), .B(n_1663), .Y(n_1661) );
OR2x2_ASAP7_75t_L g1713 ( .A(n_1662), .B(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1662), .Y(n_1752) );
OAI32xp33_ASAP7_75t_L g1790 ( .A1(n_1662), .A2(n_1667), .A3(n_1791), .B1(n_1795), .B2(n_1797), .Y(n_1790) );
AND2x2_ASAP7_75t_L g1811 ( .A(n_1662), .B(n_1685), .Y(n_1811) );
AOI21xp5_ASAP7_75t_L g1665 ( .A1(n_1666), .A2(n_1669), .B(n_1671), .Y(n_1665) );
AOI22xp5_ASAP7_75t_L g1747 ( .A1(n_1667), .A2(n_1748), .B1(n_1753), .B2(n_1757), .Y(n_1747) );
INVx2_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1669), .Y(n_1801) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
NOR2xp33_ASAP7_75t_L g1671 ( .A(n_1672), .B(n_1674), .Y(n_1671) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1672), .Y(n_1689) );
OAI21xp33_ASAP7_75t_L g1762 ( .A1(n_1672), .A2(n_1763), .B(n_1766), .Y(n_1762) );
INVx2_ASAP7_75t_L g1724 ( .A(n_1673), .Y(n_1724) );
NAND2xp5_ASAP7_75t_L g1753 ( .A(n_1673), .B(n_1754), .Y(n_1753) );
NOR2xp33_ASAP7_75t_L g1776 ( .A(n_1673), .B(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1674), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1677), .Y(n_1674) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1693 ( .A(n_1676), .B(n_1694), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1676), .B(n_1692), .Y(n_1742) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1677), .Y(n_1703) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1679), .Y(n_1802) );
A2O1A1Ixp33_ASAP7_75t_L g1700 ( .A1(n_1680), .A2(n_1701), .B(n_1704), .C(n_1708), .Y(n_1700) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1680), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1680), .B(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1686), .Y(n_1684) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1690), .Y(n_1688) );
AOI21xp5_ASAP7_75t_L g1758 ( .A1(n_1689), .A2(n_1759), .B(n_1760), .Y(n_1758) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1691), .B(n_1692), .Y(n_1690) );
INVx3_ASAP7_75t_L g1722 ( .A(n_1695), .Y(n_1722) );
NOR3xp33_ASAP7_75t_L g1743 ( .A(n_1695), .B(n_1744), .C(n_1745), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1698), .Y(n_1695) );
NAND4xp25_ASAP7_75t_SL g1699 ( .A(n_1700), .B(n_1709), .C(n_1726), .D(n_1737), .Y(n_1699) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1707), .Y(n_1705) );
O2A1O1Ixp33_ASAP7_75t_L g1709 ( .A1(n_1710), .A2(n_1712), .B(n_1715), .C(n_1716), .Y(n_1709) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
OAI21xp5_ASAP7_75t_SL g1798 ( .A1(n_1722), .A2(n_1799), .B(n_1803), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1749 ( .A(n_1724), .B(n_1750), .Y(n_1749) );
OAI221xp5_ASAP7_75t_L g1774 ( .A1(n_1724), .A2(n_1775), .B1(n_1782), .B2(n_1784), .C(n_1787), .Y(n_1774) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
AOI21xp33_ASAP7_75t_L g1732 ( .A1(n_1733), .A2(n_1734), .B(n_1735), .Y(n_1732) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1735), .Y(n_1806) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1736), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1738), .B(n_1752), .Y(n_1751) );
NOR2xp33_ASAP7_75t_L g1763 ( .A(n_1738), .B(n_1764), .Y(n_1763) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
OAI311xp33_ASAP7_75t_L g1761 ( .A1(n_1740), .A2(n_1762), .A3(n_1768), .B1(n_1773), .C1(n_1774), .Y(n_1761) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1744), .Y(n_1783) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
NOR4xp25_ASAP7_75t_L g1775 ( .A(n_1751), .B(n_1776), .C(n_1778), .D(n_1781), .Y(n_1775) );
INVx1_ASAP7_75t_L g1773 ( .A(n_1753), .Y(n_1773) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1754), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1755), .B(n_1756), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1755), .B(n_1785), .Y(n_1784) );
INVx2_ASAP7_75t_L g1792 ( .A(n_1756), .Y(n_1792) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1760), .Y(n_1769) );
INVx2_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
OAI21xp33_ASAP7_75t_SL g1768 ( .A1(n_1769), .A2(n_1770), .B(n_1772), .Y(n_1768) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
AOI21xp33_ASAP7_75t_L g1791 ( .A1(n_1772), .A2(n_1792), .B(n_1793), .Y(n_1791) );
AOI21xp33_ASAP7_75t_L g1795 ( .A1(n_1772), .A2(n_1793), .B(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
AOI21xp33_ASAP7_75t_L g1799 ( .A1(n_1800), .A2(n_1801), .B(n_1802), .Y(n_1799) );
OAI321xp33_ASAP7_75t_L g1803 ( .A1(n_1804), .A2(n_1806), .A3(n_1807), .B1(n_1809), .B2(n_1810), .C(n_1812), .Y(n_1803) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1811), .Y(n_1810) );
CKINVDCx20_ASAP7_75t_R g1813 ( .A(n_1814), .Y(n_1813) );
CKINVDCx20_ASAP7_75t_R g1814 ( .A(n_1815), .Y(n_1814) );
INVx2_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
XNOR2x1_ASAP7_75t_L g1817 ( .A(n_1818), .B(n_1819), .Y(n_1817) );
AND3x2_ASAP7_75t_L g1819 ( .A(n_1820), .B(n_1835), .C(n_1855), .Y(n_1819) );
NOR2xp33_ASAP7_75t_SL g1820 ( .A(n_1821), .B(n_1829), .Y(n_1820) );
OAI21xp5_ASAP7_75t_SL g1821 ( .A1(n_1822), .A2(n_1823), .B(n_1826), .Y(n_1821) );
NAND3xp33_ASAP7_75t_L g1836 ( .A(n_1837), .B(n_1840), .C(n_1845), .Y(n_1836) );
AOI31xp33_ASAP7_75t_L g1845 ( .A1(n_1846), .A2(n_1847), .A3(n_1849), .B(n_1850), .Y(n_1845) );
CKINVDCx20_ASAP7_75t_R g1857 ( .A(n_1858), .Y(n_1857) );
CKINVDCx20_ASAP7_75t_R g1858 ( .A(n_1859), .Y(n_1858) );
INVx3_ASAP7_75t_L g1859 ( .A(n_1860), .Y(n_1859) );
HB1xp67_ASAP7_75t_L g1863 ( .A(n_1864), .Y(n_1863) );
BUFx3_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
BUFx3_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
INVxp33_ASAP7_75t_SL g1867 ( .A(n_1868), .Y(n_1867) );
HB1xp67_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
endmodule