module fake_jpeg_14624_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_15),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_19),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_23),
.B(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_21),
.B(n_7),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_69),
.B(n_76),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_15),
.B1(n_17),
.B2(n_33),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_103),
.B(n_0),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_81),
.B(n_83),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_38),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_57),
.B1(n_59),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_109),
.B1(n_86),
.B2(n_73),
.Y(n_144)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_62),
.C(n_51),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_65),
.C(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_45),
.B(n_38),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_36),
.B1(n_29),
.B2(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_32),
.B1(n_25),
.B2(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_36),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_42),
.A2(n_66),
.B1(n_40),
.B2(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_17),
.B1(n_12),
.B2(n_10),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_18),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_114),
.B(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_18),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_135),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_117),
.B(n_91),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_75),
.A2(n_28),
.B1(n_27),
.B2(n_34),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_123),
.B1(n_106),
.B2(n_85),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_130),
.B1(n_141),
.B2(n_100),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_27),
.B1(n_34),
.B2(n_32),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_10),
.B1(n_13),
.B2(n_9),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_140),
.B1(n_145),
.B2(n_3),
.Y(n_173)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_134),
.Y(n_155)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_77),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_72),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_104),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_1),
.B(n_2),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_86),
.A2(n_3),
.B1(n_6),
.B2(n_9),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_147),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_107),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_32),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_159),
.A2(n_173),
.B1(n_184),
.B2(n_188),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_180),
.C(n_147),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_178),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_98),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_154),
.B(n_112),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_118),
.B(n_3),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_175),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_85),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_106),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_78),
.C(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_25),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_100),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_190),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_114),
.B(n_116),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_164),
.A2(n_122),
.B1(n_140),
.B2(n_131),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_191),
.A2(n_212),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_195),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_145),
.B1(n_141),
.B2(n_121),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_196),
.B(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_115),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_137),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_126),
.B1(n_125),
.B2(n_142),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_169),
.B1(n_157),
.B2(n_166),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_214),
.C(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_190),
.B1(n_176),
.B2(n_171),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_143),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_218),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_159),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_157),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_209),
.B(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_148),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_148),
.B(n_124),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_134),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_161),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_223),
.A2(n_237),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_161),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_167),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_167),
.C(n_186),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_238),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_186),
.B(n_166),
.C(n_156),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_240),
.B(n_243),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_230),
.B1(n_212),
.B2(n_226),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_179),
.B(n_155),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_163),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_174),
.B(n_169),
.Y(n_239)
);

AOI221xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_136),
.B1(n_139),
.B2(n_91),
.C(n_189),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_162),
.B(n_68),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_204),
.A2(n_185),
.B1(n_68),
.B2(n_136),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_244),
.A2(n_201),
.B1(n_192),
.B2(n_193),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_273)
);

AO221x1_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_213),
.B1(n_194),
.B2(n_220),
.C(n_197),
.Y(n_249)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_216),
.B1(n_219),
.B2(n_200),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_209),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_205),
.Y(n_255)
);

NAND4xp25_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_260),
.C(n_224),
.D(n_197),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_216),
.B1(n_192),
.B2(n_195),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_256),
.A2(n_223),
.B1(n_228),
.B2(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_261),
.B1(n_226),
.B2(n_242),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_262),
.B(n_241),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_251),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_235),
.B(n_237),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_264),
.A2(n_247),
.B(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_233),
.C(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_268),
.C(n_274),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_271),
.B1(n_275),
.B2(n_253),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_228),
.C(n_225),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_225),
.C(n_238),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_246),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_271),
.B(n_273),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_282),
.B(n_285),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_258),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_242),
.Y(n_283)
);

XOR2x2_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_266),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_267),
.B1(n_275),
.B2(n_264),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_288),
.B(n_276),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_279),
.A2(n_269),
.B(n_263),
.C(n_268),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_291),
.B1(n_274),
.B2(n_276),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_244),
.B1(n_210),
.B2(n_211),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_296),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.C(n_152),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_217),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_292),
.B(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_298),
.Y(n_302)
);


endmodule