module fake_jpeg_359_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_SL g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_21),
.B(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

OR2x4_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_1),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_23),
.B(n_10),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_58),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_60),
.B1(n_22),
.B2(n_6),
.Y(n_74)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_53),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_30),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_85),
.B1(n_74),
.B2(n_65),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_6),
.B1(n_28),
.B2(n_33),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_76),
.B1(n_72),
.B2(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_6),
.B1(n_52),
.B2(n_43),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_90),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_41),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_94),
.C(n_70),
.Y(n_122)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_48),
.C(n_34),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_49),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_110),
.B1(n_76),
.B2(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_90),
.CI(n_91),
.CON(n_107),
.SN(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_78),
.B(n_73),
.C(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_81),
.B1(n_83),
.B2(n_70),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_88),
.B1(n_107),
.B2(n_66),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_103),
.B1(n_106),
.B2(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_92),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_110),
.B(n_108),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_131),
.B1(n_111),
.B2(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_125),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_143),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_112),
.B1(n_111),
.B2(n_120),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_128),
.B1(n_130),
.B2(n_116),
.C(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_149),
.B1(n_137),
.B2(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_153),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_138),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_150),
.C(n_146),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_148),
.B1(n_136),
.B2(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_144),
.Y(n_162)
);

OAI221xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_156),
.B1(n_144),
.B2(n_114),
.C(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_159),
.C(n_123),
.Y(n_164)
);

OAI21x1_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_124),
.B(n_123),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_95),
.C(n_72),
.Y(n_166)
);


endmodule