module fake_jpeg_5483_n_327 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_18),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_13),
.B1(n_15),
.B2(n_27),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_15),
.B1(n_27),
.B2(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_60),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_78),
.B1(n_37),
.B2(n_13),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_66),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_24),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_50),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_26),
.A3(n_23),
.B1(n_22),
.B2(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_76),
.Y(n_89)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_37),
.B1(n_35),
.B2(n_29),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_37),
.B1(n_49),
.B2(n_28),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_95),
.B1(n_101),
.B2(n_71),
.Y(n_122)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_84),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_41),
.B(n_28),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_99),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_17),
.B(n_31),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_27),
.B1(n_15),
.B2(n_14),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_13),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_13),
.B1(n_15),
.B2(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_122),
.B1(n_101),
.B2(n_80),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_101),
.B(n_68),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_107),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_117),
.Y(n_141)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_79),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_140),
.B1(n_149),
.B2(n_15),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_132),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_88),
.C(n_85),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_139),
.C(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_91),
.Y(n_132)
);

OR2x6_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_80),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_162)
);

OAI31xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_93),
.A3(n_101),
.B(n_98),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_90),
.C(n_91),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_93),
.B1(n_92),
.B2(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_25),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_31),
.B(n_17),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_78),
.B(n_19),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_79),
.B1(n_54),
.B2(n_50),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_151),
.A2(n_14),
.B1(n_70),
.B2(n_69),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_109),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_171),
.C(n_142),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_165),
.B1(n_169),
.B2(n_174),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_160),
.B(n_170),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_176),
.B1(n_178),
.B2(n_138),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_27),
.A3(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_173),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_62),
.B1(n_54),
.B2(n_35),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_43),
.B1(n_48),
.B2(n_73),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_38),
.C(n_39),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_138),
.B1(n_140),
.B2(n_128),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_24),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_83),
.B(n_23),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_128),
.B1(n_133),
.B2(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_190),
.C(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_137),
.B1(n_133),
.B2(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_173),
.B1(n_158),
.B2(n_154),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_150),
.B(n_145),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_188),
.B(n_204),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_142),
.B1(n_14),
.B2(n_136),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_52),
.B1(n_48),
.B2(n_123),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_14),
.B1(n_83),
.B2(n_114),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_30),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_200),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_30),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_76),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_218),
.B(n_227),
.Y(n_241)
);

OAI321xp33_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_164),
.A3(n_153),
.B1(n_177),
.B2(n_174),
.C(n_163),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_26),
.B(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_99),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_86),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_224),
.B1(n_226),
.B2(n_200),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_171),
.B1(n_161),
.B2(n_120),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_231),
.B1(n_248),
.B2(n_71),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_215),
.A2(n_182),
.B1(n_180),
.B2(n_191),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_190),
.C(n_195),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_243),
.C(n_244),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_185),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_238),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_198),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_191),
.B1(n_180),
.B2(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_240),
.A2(n_228),
.B1(n_208),
.B2(n_226),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_204),
.C(n_39),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_94),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_94),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_246),
.C(n_223),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_94),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_207),
.A2(n_217),
.B1(n_228),
.B2(n_221),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_214),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_253),
.B(n_259),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_267),
.B1(n_268),
.B2(n_25),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_262),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_223),
.CI(n_21),
.CON(n_258),
.SN(n_258)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_96),
.C(n_77),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_25),
.C(n_17),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_242),
.A2(n_233),
.B1(n_229),
.B2(n_235),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_261),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_245),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_264),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_25),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_247),
.B(n_8),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_8),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_241),
.A2(n_25),
.B1(n_17),
.B2(n_2),
.Y(n_268)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_244),
.B(n_234),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_270),
.A2(n_10),
.B(n_9),
.Y(n_297)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_253),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_17),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_279),
.C(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_25),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_12),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_25),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_25),
.C(n_20),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_258),
.C(n_20),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_285),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_260),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_277),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_261),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_291),
.B(n_294),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_254),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_11),
.C(n_10),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_297),
.B(n_9),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_269),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_303),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_289),
.C(n_284),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_293),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_290),
.A2(n_3),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_4),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_5),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_312),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_311),
.Y(n_318)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_305),
.B1(n_300),
.B2(n_307),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_315),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_304),
.B(n_7),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_310),
.B(n_313),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.C(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_318),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_20),
.C(n_6),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_7),
.B(n_20),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_7),
.B(n_20),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_20),
.Y(n_327)
);


endmodule