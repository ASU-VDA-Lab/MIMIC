module fake_jpeg_22242_n_109 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx5_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_14),
.B(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_31),
.B1(n_29),
.B2(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_41),
.B1(n_47),
.B2(n_17),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_17),
.B1(n_24),
.B2(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_21),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_21),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_20),
.B(n_15),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_36),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_33),
.B(n_34),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_56),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_59),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_61),
.B1(n_40),
.B2(n_11),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_21),
.B(n_11),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_22),
.B1(n_16),
.B2(n_19),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_22),
.B1(n_11),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_66),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_59),
.B(n_56),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_51),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_73),
.C(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_57),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_67),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.C(n_91),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_84),
.C(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_72),
.C(n_68),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_77),
.B(n_83),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_73),
.B(n_85),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_78),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_96),
.C(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_66),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_98),
.B(n_72),
.Y(n_101)
);

XNOR2x1_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_58),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_55),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_104),
.B(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_62),
.CI(n_9),
.CON(n_109),
.SN(n_109)
);


endmodule