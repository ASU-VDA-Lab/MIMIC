module real_jpeg_21071_n_12 (n_5, n_4, n_8, n_0, n_280, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_280;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_244;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_3),
.B1(n_18),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_0),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_0),
.A2(n_9),
.B(n_27),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_0),
.B(n_28),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g187 ( 
.A1(n_0),
.A2(n_10),
.B(n_66),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_0),
.A2(n_40),
.B(n_41),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_1),
.A2(n_3),
.B1(n_18),
.B2(n_19),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_1),
.A2(n_19),
.B1(n_65),
.B2(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_3),
.B1(n_18),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_3),
.A2(n_4),
.B1(n_18),
.B2(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_3),
.A2(n_23),
.B(n_50),
.C(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_30),
.B1(n_39),
.B2(n_40),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_39),
.B1(n_40),
.B2(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

BUFx3_ASAP7_75t_SL g40 ( 
.A(n_11),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_273),
.B(n_276),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_68),
.B(n_272),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_31),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_15),
.B(n_31),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_15),
.B(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_25),
.B(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_22),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_21),
.B(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_38),
.B(n_41),
.C(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_41),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_27),
.A2(n_42),
.B(n_50),
.C(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_48),
.B(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_29),
.B(n_83),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_32),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_32),
.B(n_270),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_46),
.CI(n_51),
.CON(n_32),
.SN(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_34),
.A2(n_37),
.B1(n_43),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_36),
.B(n_95),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_37),
.A2(n_94),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_38),
.A2(n_44),
.B1(n_93),
.B2(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_38),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_38),
.B(n_50),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_40),
.A2(n_50),
.B(n_63),
.C(n_187),
.Y(n_186)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_44),
.B(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_50),
.B(n_79),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_50),
.B(n_64),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_58),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_100),
.C(n_105),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_52),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_52),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_92),
.B1(n_127),
.B2(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_52),
.B(n_154),
.C(n_155),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_52),
.A2(n_105),
.B1(n_127),
.B2(n_165),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_56),
.A2(n_58),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_56),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_60),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_64),
.B1(n_67),
.B2(n_87),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_64),
.B1(n_90),
.B2(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_65),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_269),
.B(n_271),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_122),
.A3(n_133),
.B1(n_267),
.B2(n_268),
.C(n_280),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_107),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_71),
.B(n_107),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_91),
.C(n_98),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_72),
.B(n_91),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_82),
.B2(n_84),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_74),
.A2(n_75),
.B1(n_86),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_82),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_77),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_80),
.B1(n_81),
.B2(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_78),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_78),
.A2(n_79),
.B1(n_148),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_79),
.A2(n_102),
.B(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_96),
.B(n_97),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_92),
.B(n_171),
.C(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_92),
.A2(n_154),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_109),
.C(n_119),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_98),
.A2(n_99),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_100),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_101),
.A2(n_103),
.B1(n_202),
.B2(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_101),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_103),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_103),
.B(n_159),
.C(n_201),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_103),
.A2(n_202),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_103),
.B(n_220),
.C(n_225),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_110),
.C(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_150),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_105),
.A2(n_140),
.B1(n_141),
.B2(n_165),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_105),
.B(n_141),
.C(n_208),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_118),
.B1(n_126),
.B2(n_131),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_118),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_110),
.A2(n_118),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_110),
.B(n_242),
.C(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_117),
.C(n_118),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_118),
.B(n_131),
.C(n_132),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_123),
.B(n_124),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_261),
.B(n_266),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_249),
.B(n_260),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_177),
.B(n_234),
.C(n_248),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_161),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_161),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_139),
.B(n_149),
.C(n_152),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_141),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_140),
.B(n_145),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_141),
.B(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_193),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_169),
.B1(n_199),
.B2(n_203),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.C(n_170),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_162),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_233),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_227),
.B(n_232),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_217),
.B(n_226),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_205),
.B(n_216),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_196),
.B(n_204),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_188),
.B(n_195),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B(n_194),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_207),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_214),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_214),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_236),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_246),
.B2(n_247),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_241),
.C(n_247),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_257),
.C(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);


endmodule