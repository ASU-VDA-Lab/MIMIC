module fake_jpeg_2040_n_159 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_50),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_54),
.B1(n_41),
.B2(n_48),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_47),
.B1(n_56),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_61),
.B1(n_60),
.B2(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_72),
.B1(n_50),
.B2(n_53),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_42),
.B1(n_54),
.B2(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_56),
.B1(n_48),
.B2(n_53),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_48),
.B1(n_53),
.B2(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_44),
.B1(n_47),
.B2(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_90),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_103)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_79),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_93),
.A2(n_76),
.B1(n_73),
.B2(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_104),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_99),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_58),
.B(n_2),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_89),
.C(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_102),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_58),
.B1(n_23),
.B2(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_28),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_4),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_8),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_8),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_122),
.B1(n_125),
.B2(n_17),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_13),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_15),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_39),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_94),
.B(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_131),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_108),
.B(n_19),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_112),
.A2(n_20),
.B1(n_27),
.B2(n_29),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_125),
.B1(n_36),
.B2(n_37),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_31),
.C(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_114),
.A3(n_121),
.B1(n_115),
.B2(n_126),
.C1(n_113),
.C2(n_122),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_140),
.B(n_127),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_138),
.A2(n_35),
.B1(n_38),
.B2(n_128),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_149),
.C(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_135),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_142),
.B1(n_141),
.B2(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_140),
.B1(n_131),
.B2(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_134),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_130),
.B(n_154),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_146),
.Y(n_159)
);


endmodule