module fake_jpeg_12785_n_494 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_494);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_494;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_51),
.B(n_54),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_60),
.B(n_72),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_19),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_71),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_17),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_76),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_29),
.A2(n_16),
.B1(n_13),
.B2(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_44),
.B1(n_33),
.B2(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_83),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_34),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_85),
.Y(n_139)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_89),
.B(n_93),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_26),
.Y(n_104)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_30),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_16),
.B(n_35),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_94),
.A2(n_105),
.B1(n_112),
.B2(n_142),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_29),
.B1(n_42),
.B2(n_26),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_100),
.A2(n_109),
.B(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_117),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_104),
.B(n_115),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_86),
.B1(n_65),
.B2(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_22),
.B1(n_39),
.B2(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_45),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_22),
.B1(n_39),
.B2(n_36),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_45),
.B(n_25),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g198 ( 
.A(n_118),
.B(n_5),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_35),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_32),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_31),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_67),
.B(n_46),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_140),
.B(n_36),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_52),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_73),
.B(n_46),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_18),
.B1(n_20),
.B2(n_39),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_159),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_79),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_41),
.B(n_61),
.C(n_44),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_167),
.B(n_182),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_56),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_168),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_33),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_44),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_184),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_188),
.B1(n_145),
.B2(n_125),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_1),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_181),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_58),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_175),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_62),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_39),
.B1(n_36),
.B2(n_20),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_198),
.B1(n_201),
.B2(n_138),
.Y(n_243)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_180),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_1),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_119),
.B(n_62),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_105),
.A2(n_80),
.B1(n_88),
.B2(n_91),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_82),
.B1(n_78),
.B2(n_76),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_189),
.A2(n_141),
.B(n_124),
.Y(n_241)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_106),
.B(n_3),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_6),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_100),
.B(n_3),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_196),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_94),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_90),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_199),
.B(n_203),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_122),
.A2(n_53),
.B(n_6),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_12),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_109),
.A2(n_69),
.B1(n_6),
.B2(n_7),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_132),
.B(n_5),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_149),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_207),
.Y(n_257)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_129),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_131),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_209),
.Y(n_236)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_210),
.B(n_11),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_211),
.A2(n_141),
.B1(n_129),
.B2(n_124),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_157),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_255),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_152),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_218),
.B(n_241),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_155),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_176),
.A2(n_136),
.B1(n_99),
.B2(n_150),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_176),
.A2(n_136),
.B1(n_99),
.B2(n_123),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_163),
.A2(n_138),
.B1(n_149),
.B2(n_152),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_194),
.A2(n_159),
.B1(n_201),
.B2(n_158),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_243),
.A2(n_208),
.B1(n_168),
.B2(n_185),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_163),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_246),
.B1(n_261),
.B2(n_208),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_173),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_161),
.B(n_169),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_250),
.B(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_154),
.B(n_9),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_259),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_172),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_11),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_206),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_183),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_158),
.A2(n_156),
.B1(n_189),
.B2(n_170),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_263),
.B(n_268),
.Y(n_341)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_233),
.A2(n_184),
.B1(n_166),
.B2(n_199),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_266),
.A2(n_270),
.B1(n_296),
.B2(n_303),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_215),
.B(n_174),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_205),
.B1(n_197),
.B2(n_177),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_225),
.A2(n_249),
.B(n_222),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_257),
.B(n_251),
.Y(n_309)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_218),
.A2(n_198),
.B1(n_187),
.B2(n_167),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_274),
.A2(n_298),
.B(n_292),
.Y(n_332)
);

AO21x1_ASAP7_75t_SL g275 ( 
.A1(n_247),
.A2(n_195),
.B(n_161),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_242),
.B(n_213),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_222),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_276),
.A2(n_304),
.B(n_238),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_277),
.Y(n_311)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_281),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_160),
.B1(n_204),
.B2(n_202),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_212),
.B(n_162),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_212),
.B(n_164),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_214),
.B(n_181),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_221),
.B(n_168),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_295),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_192),
.B1(n_165),
.B2(n_180),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_249),
.A2(n_211),
.B1(n_178),
.B2(n_209),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_161),
.B1(n_190),
.B2(n_171),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_171),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_293),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_190),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_191),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_299),
.B1(n_301),
.B2(n_223),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_218),
.A2(n_175),
.B1(n_177),
.B2(n_186),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_221),
.B(n_175),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_300),
.B(n_307),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_239),
.A2(n_12),
.B1(n_186),
.B2(n_245),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_236),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_305),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_239),
.A2(n_186),
.B1(n_222),
.B2(n_245),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_236),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_227),
.B(n_259),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_226),
.B1(n_241),
.B2(n_230),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_309),
.B(n_334),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_250),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_329),
.C(n_331),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_291),
.A2(n_228),
.B(n_217),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_318),
.A2(n_326),
.B(n_328),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_319),
.B(n_344),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_282),
.A2(n_230),
.B1(n_228),
.B2(n_252),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_321),
.A2(n_281),
.B1(n_278),
.B2(n_267),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_272),
.A2(n_229),
.B1(n_252),
.B2(n_242),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_333),
.B1(n_339),
.B2(n_289),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_330),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_223),
.B(n_220),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_269),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_332),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_223),
.B(n_220),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_271),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_219),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_300),
.B(n_219),
.C(n_231),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_272),
.A2(n_229),
.B1(n_231),
.B2(n_238),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_229),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_346),
.C(n_290),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_296),
.A2(n_253),
.B1(n_269),
.B2(n_274),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_340),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_294),
.A2(n_253),
.B(n_303),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_302),
.C(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_316),
.Y(n_349)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_263),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_357),
.Y(n_400)
);

AO32x1_ASAP7_75t_L g354 ( 
.A1(n_311),
.A2(n_275),
.A3(n_277),
.B1(n_306),
.B2(n_297),
.Y(n_354)
);

OAI21xp33_ASAP7_75t_L g391 ( 
.A1(n_354),
.A2(n_342),
.B(n_314),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_324),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_341),
.B(n_286),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_358),
.B(n_362),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_338),
.Y(n_401)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_320),
.Y(n_361)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_268),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_345),
.Y(n_363)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_295),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_374),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_365),
.A2(n_367),
.B1(n_368),
.B2(n_370),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_301),
.B1(n_285),
.B2(n_275),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_322),
.A2(n_262),
.B1(n_287),
.B2(n_265),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_280),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_372),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_323),
.A2(n_262),
.B1(n_264),
.B2(n_273),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_323),
.A2(n_279),
.B1(n_305),
.B2(n_280),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_371),
.A2(n_380),
.B1(n_377),
.B2(n_368),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_376),
.B(n_379),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_343),
.B1(n_333),
.B2(n_314),
.Y(n_393)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_342),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_346),
.C(n_337),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_384),
.C(n_386),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_379),
.A2(n_311),
.B1(n_319),
.B2(n_317),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_382),
.A2(n_359),
.B1(n_378),
.B2(n_354),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_329),
.C(n_330),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_332),
.C(n_325),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_325),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_398),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_350),
.B(n_315),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_389),
.B(n_371),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_367),
.Y(n_427)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_355),
.B(n_331),
.C(n_309),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_401),
.C(n_381),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_318),
.CI(n_326),
.CON(n_395),
.SN(n_395)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_356),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_375),
.A2(n_328),
.B1(n_317),
.B2(n_344),
.Y(n_397)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_397),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_336),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_375),
.A2(n_338),
.B1(n_336),
.B2(n_278),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_404),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_267),
.B1(n_359),
.B2(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_405),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_410),
.A2(n_415),
.B1(n_422),
.B2(n_413),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_411),
.A2(n_428),
.B(n_395),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_382),
.B1(n_391),
.B2(n_394),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_429),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_387),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_418),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_424),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_366),
.B(n_355),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_423),
.B(n_420),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_402),
.A2(n_349),
.B1(n_351),
.B2(n_361),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_395),
.A2(n_366),
.B(n_370),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_390),
.Y(n_426)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_363),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_365),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_396),
.Y(n_431)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_431),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_403),
.Y(n_434)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_434),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_416),
.A2(n_397),
.B(n_399),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_435),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_420),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_437),
.B(n_441),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_438),
.B(n_389),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_398),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_413),
.A2(n_401),
.B1(n_402),
.B2(n_393),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_443),
.A2(n_423),
.B1(n_421),
.B2(n_427),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_445),
.A2(n_424),
.B1(n_386),
.B2(n_373),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_446),
.A2(n_385),
.B1(n_374),
.B2(n_376),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_388),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_450),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_407),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_444),
.A2(n_415),
.B(n_410),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_455),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_453),
.A2(n_458),
.B1(n_436),
.B2(n_440),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_434),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_456),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_443),
.B1(n_439),
.B2(n_448),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_440),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_459),
.B(n_460),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_444),
.A2(n_419),
.B(n_417),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_L g470 ( 
.A1(n_462),
.A2(n_449),
.B(n_433),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_432),
.B(n_429),
.C(n_417),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_439),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_461),
.A2(n_446),
.B1(n_437),
.B2(n_432),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_471),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_433),
.B1(n_441),
.B2(n_450),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_467),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_468),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_474),
.C(n_454),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_457),
.Y(n_480)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_454),
.A2(n_442),
.B(n_447),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_466),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_473),
.A2(n_464),
.B(n_460),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_480),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_451),
.Y(n_481)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_481),
.Y(n_484)
);

A2O1A1Ixp33_ASAP7_75t_L g482 ( 
.A1(n_475),
.A2(n_473),
.B(n_470),
.C(n_474),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_482),
.A2(n_483),
.B(n_452),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_486),
.A2(n_488),
.B(n_465),
.Y(n_489)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g487 ( 
.A1(n_484),
.A2(n_478),
.B(n_476),
.C(n_479),
.D(n_459),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_487),
.B(n_463),
.Y(n_490)
);

NOR3xp33_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_490),
.C(n_463),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g492 ( 
.A(n_491),
.B(n_442),
.C(n_447),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_448),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_493),
.B(n_472),
.Y(n_494)
);


endmodule