module fake_netlist_6_4330_n_799 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_799);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_799;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_83),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_9),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_56),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_113),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_49),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_36),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_33),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_61),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_32),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_128),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_131),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_18),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_134),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_17),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_77),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_71),
.B(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_42),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_117),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_35),
.B(n_145),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_59),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_80),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_46),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_15),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_86),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_34),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_84),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_191),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

BUFx8_ASAP7_75t_SL g222 ( 
.A(n_171),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_2),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_171),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_163),
.B(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_3),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_164),
.B(n_4),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_159),
.A2(n_5),
.B(n_6),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_162),
.B(n_5),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_179),
.B(n_158),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_165),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_166),
.Y(n_247)
);

AOI22x1_ASAP7_75t_SL g248 ( 
.A1(n_188),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_172),
.B(n_10),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_194),
.B1(n_198),
.B2(n_175),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_174),
.B(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

OAI22x1_ASAP7_75t_L g254 ( 
.A1(n_181),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_182),
.B(n_192),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

AOI22x1_ASAP7_75t_SL g258 ( 
.A1(n_199),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_200),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_208),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_213),
.C(n_210),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_239),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_214),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_169),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_212),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_209),
.C(n_205),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_229),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

AO21x2_ASAP7_75t_L g288 ( 
.A1(n_240),
.A2(n_174),
.B(n_202),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_252),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_239),
.B(n_170),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_242),
.B(n_173),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_216),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_203),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_235),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_225),
.B(n_176),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_229),
.B(n_180),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_215),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_238),
.C(n_215),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_276),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_232),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_232),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_275),
.A2(n_244),
.B1(n_240),
.B2(n_219),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_244),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_242),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_249),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_295),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_253),
.C(n_256),
.Y(n_320)
);

AND2x4_ASAP7_75t_SL g321 ( 
.A(n_266),
.B(n_239),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_242),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_224),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_224),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_231),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_231),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_184),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_275),
.B(n_236),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_266),
.B(n_217),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_275),
.B(n_236),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_277),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_251),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_217),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_217),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_279),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_272),
.B(n_251),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_274),
.B(n_217),
.Y(n_340)
);

NOR2x1p5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_227),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_297),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_293),
.B(n_298),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_285),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_251),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_282),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_287),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_299),
.A2(n_254),
.B1(n_245),
.B2(n_227),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_256),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_287),
.B(n_256),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_290),
.B(n_253),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_299),
.B(n_185),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_282),
.B(n_246),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_223),
.C(n_230),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_288),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_290),
.B(n_246),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_283),
.B(n_246),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_302),
.B(n_247),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_294),
.B(n_247),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_294),
.Y(n_369)
);

AO221x1_ASAP7_75t_L g370 ( 
.A1(n_288),
.A2(n_254),
.B1(n_219),
.B2(n_216),
.C(n_226),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_301),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_288),
.B(n_230),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_302),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_321),
.B(n_303),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_314),
.A2(n_307),
.B(n_303),
.Y(n_376)
);

NAND2x1_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_301),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_312),
.B(n_259),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_307),
.B(n_262),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_317),
.A2(n_322),
.B(n_331),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_313),
.A2(n_273),
.B(n_284),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_314),
.A2(n_247),
.B(n_269),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_338),
.B(n_190),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_312),
.B(n_223),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_336),
.A2(n_337),
.B(n_343),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_346),
.B(n_262),
.Y(n_386)
);

AOI21xp33_ASAP7_75t_L g387 ( 
.A1(n_309),
.A2(n_335),
.B(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_193),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_264),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_340),
.A2(n_273),
.B(n_284),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_363),
.A2(n_269),
.B(n_268),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_326),
.B(n_197),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_328),
.B(n_201),
.Y(n_395)
);

O2A1O1Ixp5_ASAP7_75t_L g396 ( 
.A1(n_372),
.A2(n_264),
.B(n_267),
.C(n_268),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_334),
.B(n_323),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_357),
.A2(n_273),
.B(n_284),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_362),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_273),
.B(n_284),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_267),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_330),
.A2(n_260),
.B1(n_233),
.B2(n_226),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_332),
.A2(n_260),
.B(n_258),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_226),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_339),
.A2(n_284),
.B(n_233),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_319),
.B(n_226),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_319),
.B(n_226),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_308),
.A2(n_284),
.B(n_233),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_310),
.B(n_226),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_370),
.A2(n_233),
.B1(n_258),
.B2(n_248),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_324),
.B(n_233),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_356),
.A2(n_248),
.B(n_233),
.C(n_17),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_329),
.A2(n_273),
.B(n_85),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_315),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_326),
.B(n_15),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_323),
.B(n_16),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_344),
.B(n_21),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_360),
.B(n_16),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_347),
.B(n_22),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_349),
.A2(n_88),
.B1(n_24),
.B2(n_25),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_367),
.A2(n_361),
.B(n_365),
.C(n_366),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_364),
.A2(n_89),
.B(n_26),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_345),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_367),
.B(n_19),
.Y(n_434)
);

OAI321xp33_ASAP7_75t_L g435 ( 
.A1(n_356),
.A2(n_19),
.A3(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_368),
.A2(n_31),
.B(n_37),
.C(n_38),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_361),
.A2(n_40),
.B(n_41),
.C(n_43),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_365),
.A2(n_44),
.B(n_45),
.C(n_48),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_369),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_440)
);

O2A1O1Ixp33_ASAP7_75t_L g441 ( 
.A1(n_351),
.A2(n_54),
.B(n_55),
.C(n_57),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_424),
.A2(n_353),
.B(n_352),
.Y(n_443)
);

AOI21x1_ASAP7_75t_SL g444 ( 
.A1(n_426),
.A2(n_350),
.B(n_371),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_436),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_388),
.B(n_350),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

AO31x2_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_350),
.A3(n_60),
.B(n_62),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_399),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_450)
);

AO21x2_ASAP7_75t_L g451 ( 
.A1(n_376),
.A2(n_65),
.B(n_66),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_376),
.A2(n_67),
.B(n_68),
.Y(n_452)
);

AOI21x1_ASAP7_75t_SL g453 ( 
.A1(n_428),
.A2(n_69),
.B(n_70),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_425),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_72),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_396),
.A2(n_157),
.B(n_75),
.Y(n_457)
);

NOR2x1_ASAP7_75t_SL g458 ( 
.A(n_418),
.B(n_74),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_413),
.B(n_76),
.Y(n_459)
);

AO21x1_ASAP7_75t_L g460 ( 
.A1(n_387),
.A2(n_78),
.B(n_79),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_380),
.A2(n_156),
.B(n_82),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_408),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_402),
.B(n_81),
.Y(n_463)
);

AOI21x1_ASAP7_75t_SL g464 ( 
.A1(n_434),
.A2(n_87),
.B(n_94),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_417),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_404),
.B(n_98),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_373),
.A2(n_99),
.B(n_100),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_384),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_390),
.B(n_103),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_427),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_406),
.B(n_108),
.Y(n_471)
);

AO21x2_ASAP7_75t_L g472 ( 
.A1(n_393),
.A2(n_155),
.B(n_110),
.Y(n_472)
);

AO21x2_ASAP7_75t_L g473 ( 
.A1(n_393),
.A2(n_382),
.B(n_410),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_382),
.A2(n_109),
.B(n_111),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_397),
.B(n_114),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_423),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_115),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_386),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_118),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_420),
.A2(n_389),
.B1(n_432),
.B2(n_375),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_374),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_385),
.A2(n_379),
.B(n_403),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_409),
.B(n_119),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_377),
.A2(n_154),
.B(n_122),
.Y(n_486)
);

OA22x2_ASAP7_75t_L g487 ( 
.A1(n_423),
.A2(n_120),
.B1(n_127),
.B2(n_130),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_418),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_383),
.B(n_132),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_435),
.A2(n_133),
.B(n_136),
.C(n_138),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_412),
.A2(n_414),
.B(n_421),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_438),
.B(n_140),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_410),
.A2(n_141),
.B(n_142),
.Y(n_494)
);

A2O1A1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_144),
.B(n_146),
.C(n_147),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_415),
.A2(n_148),
.B(n_150),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_151),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_441),
.A2(n_153),
.B(n_437),
.C(n_439),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_394),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_407),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_416),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_444),
.A2(n_419),
.B(n_431),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_483),
.A2(n_440),
.B(n_415),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_442),
.B(n_429),
.Y(n_504)
);

NAND2x1p5_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_381),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_492),
.A2(n_398),
.B(n_392),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_457),
.A2(n_400),
.B(n_461),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_478),
.A2(n_483),
.B(n_459),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_468),
.Y(n_512)
);

CKINVDCx11_ASAP7_75t_R g513 ( 
.A(n_475),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_485),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_491),
.A2(n_495),
.B1(n_459),
.B2(n_481),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_469),
.B(n_474),
.Y(n_517)
);

NAND2x1p5_ASAP7_75t_L g518 ( 
.A(n_466),
.B(n_499),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_453),
.B(n_486),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_474),
.A2(n_452),
.B(n_494),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_477),
.Y(n_521)
);

AOI22x1_ASAP7_75t_L g522 ( 
.A1(n_452),
.A2(n_493),
.B1(n_480),
.B2(n_494),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_447),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_484),
.A2(n_473),
.B(n_497),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_490),
.A2(n_467),
.B(n_489),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_455),
.A2(n_443),
.B(n_496),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_473),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_466),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_496),
.A2(n_460),
.B(n_487),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_476),
.A2(n_499),
.B1(n_463),
.B2(n_471),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_487),
.A2(n_450),
.B(n_456),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

OAI221xp5_ASAP7_75t_L g535 ( 
.A1(n_465),
.A2(n_450),
.B1(n_470),
.B2(n_498),
.C(n_493),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_458),
.C(n_451),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_451),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_449),
.A2(n_444),
.B(n_492),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_449),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_472),
.B(n_499),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_472),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_483),
.A2(n_382),
.B(n_474),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_479),
.B(n_401),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_465),
.A2(n_275),
.B1(n_487),
.B2(n_370),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_445),
.Y(n_546)
);

AO21x1_ASAP7_75t_L g547 ( 
.A1(n_452),
.A2(n_474),
.B(n_424),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_465),
.A2(n_275),
.B1(n_487),
.B2(n_370),
.Y(n_548)
);

NAND2x1_ASAP7_75t_L g549 ( 
.A(n_442),
.B(n_374),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_444),
.A2(n_492),
.B(n_457),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_506),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_506),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_514),
.B(n_515),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_518),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_514),
.B(n_500),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_550),
.A2(n_538),
.B(n_508),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_545),
.B(n_548),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_547),
.A2(n_510),
.B(n_517),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_511),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

INVxp33_ASAP7_75t_L g566 ( 
.A(n_543),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_512),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_512),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_522),
.A2(n_535),
.B1(n_520),
.B2(n_545),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_520),
.B(n_540),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_548),
.A2(n_520),
.B1(n_516),
.B2(n_536),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_530),
.B(n_525),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_546),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_551),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_533),
.B(n_524),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_533),
.A2(n_518),
.B1(n_530),
.B2(n_544),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_524),
.B(n_501),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_528),
.Y(n_579)
);

AO21x1_ASAP7_75t_SL g580 ( 
.A1(n_532),
.A2(n_531),
.B(n_534),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_521),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_550),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_530),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_505),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_509),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_505),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_530),
.B(n_523),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_549),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_539),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_513),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_531),
.B(n_504),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_527),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_537),
.A2(n_526),
.B1(n_541),
.B2(n_503),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_558),
.B(n_503),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_558),
.B(n_541),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_588),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_555),
.B(n_513),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_555),
.B(n_519),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_571),
.A2(n_519),
.B1(n_502),
.B2(n_508),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_581),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_578),
.B(n_507),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_578),
.B(n_575),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_581),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_571),
.A2(n_569),
.B1(n_561),
.B2(n_563),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_584),
.B(n_556),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_575),
.B(n_576),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_584),
.B(n_556),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_589),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

OA21x2_ASAP7_75t_L g615 ( 
.A1(n_559),
.A2(n_595),
.B(n_579),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_563),
.B(n_562),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_591),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_568),
.B(n_589),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_591),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_567),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_560),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_564),
.B(n_573),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_560),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_564),
.B(n_573),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_561),
.A2(n_577),
.B1(n_588),
.B2(n_566),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_556),
.B(n_594),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_589),
.B(n_567),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_553),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_584),
.B(n_572),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_554),
.B(n_565),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_583),
.B(n_586),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_560),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_592),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_588),
.A2(n_594),
.B1(n_572),
.B2(n_596),
.Y(n_634)
);

BUFx2_ASAP7_75t_SL g635 ( 
.A(n_572),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_588),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_572),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_583),
.A2(n_586),
.B1(n_593),
.B2(n_570),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

NOR2x1_ASAP7_75t_SL g641 ( 
.A(n_580),
.B(n_593),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_616),
.B(n_563),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_605),
.B(n_563),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_621),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_605),
.B(n_574),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_610),
.B(n_574),
.Y(n_646)
);

NAND2x1p5_ASAP7_75t_L g647 ( 
.A(n_599),
.B(n_587),
.Y(n_647)
);

INVx3_ASAP7_75t_SL g648 ( 
.A(n_633),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_614),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_603),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_622),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_604),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_614),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_621),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_610),
.B(n_580),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_597),
.B(n_579),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_585),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_597),
.B(n_557),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_613),
.B(n_557),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_629),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_613),
.B(n_557),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_616),
.B(n_570),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_SL g663 ( 
.A(n_600),
.B(n_585),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_612),
.B(n_585),
.Y(n_664)
);

BUFx4f_ASAP7_75t_SL g665 ( 
.A(n_603),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_626),
.B(n_587),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_623),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_607),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_623),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_618),
.B(n_587),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_607),
.B(n_587),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_626),
.B(n_590),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_598),
.B(n_570),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_633),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_622),
.Y(n_675)
);

OR2x2_ASAP7_75t_SL g676 ( 
.A(n_620),
.B(n_627),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_632),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_626),
.B(n_590),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_598),
.B(n_595),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_606),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_608),
.B(n_582),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_680),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_652),
.B(n_641),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_641),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_657),
.B(n_664),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_670),
.B(n_628),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_650),
.B(n_628),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_680),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_644),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_644),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_654),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_654),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_668),
.B(n_619),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_615),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_658),
.B(n_604),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_667),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_658),
.B(n_615),
.Y(n_697)
);

AOI211xp5_ASAP7_75t_L g698 ( 
.A1(n_663),
.A2(n_625),
.B(n_634),
.C(n_639),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_667),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_675),
.B(n_619),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_675),
.B(n_617),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_665),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_656),
.B(n_615),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_669),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_672),
.B(n_638),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_677),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_656),
.B(n_615),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_655),
.B(n_640),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_642),
.B(n_601),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_677),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_651),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_660),
.B(n_617),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_659),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_663),
.B(n_602),
.C(n_638),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_692),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_710),
.B(n_662),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_692),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_695),
.B(n_660),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_689),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_699),
.Y(n_722)
);

AO221x1_ASAP7_75t_L g723 ( 
.A1(n_704),
.A2(n_599),
.B1(n_636),
.B2(n_637),
.C(n_649),
.Y(n_723)
);

AND2x4_ASAP7_75t_SL g724 ( 
.A(n_683),
.B(n_660),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_695),
.B(n_655),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_682),
.Y(n_726)
);

OAI33xp33_ASAP7_75t_L g727 ( 
.A1(n_687),
.A2(n_671),
.A3(n_643),
.B1(n_679),
.B2(n_674),
.B3(n_645),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_710),
.B(n_646),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_706),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_709),
.B(n_673),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_694),
.B(n_662),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_698),
.A2(n_666),
.B1(n_629),
.B2(n_678),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_709),
.B(n_673),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_685),
.B(n_703),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_683),
.B(n_661),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_716),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_718),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_727),
.A2(n_715),
.B1(n_705),
.B2(n_666),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_731),
.B(n_694),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_734),
.B(n_713),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_735),
.B(n_684),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_735),
.B(n_684),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_720),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_726),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_732),
.B(n_702),
.Y(n_745)
);

INVxp67_ASAP7_75t_SL g746 ( 
.A(n_726),
.Y(n_746)
);

NOR2x1_ASAP7_75t_L g747 ( 
.A(n_734),
.B(n_702),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_724),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_721),
.Y(n_749)
);

AOI321xp33_ASAP7_75t_L g750 ( 
.A1(n_738),
.A2(n_686),
.A3(n_705),
.B1(n_728),
.B2(n_693),
.C(n_722),
.Y(n_750)
);

OAI222xp33_ASAP7_75t_L g751 ( 
.A1(n_747),
.A2(n_717),
.B1(n_728),
.B2(n_719),
.C1(n_725),
.C2(n_702),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_745),
.A2(n_727),
.B(n_723),
.Y(n_752)
);

OAI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_740),
.A2(n_729),
.B1(n_712),
.B2(n_648),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_748),
.A2(n_701),
.B1(n_700),
.B2(n_714),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

AOI22x1_ASAP7_75t_L g756 ( 
.A1(n_746),
.A2(n_674),
.B1(n_648),
.B2(n_707),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_752),
.A2(n_743),
.B(n_749),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_753),
.A2(n_666),
.B1(n_743),
.B2(n_678),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_754),
.B(n_737),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_751),
.B(n_742),
.Y(n_760)
);

AOI211xp5_ASAP7_75t_L g761 ( 
.A1(n_750),
.A2(n_736),
.B(n_739),
.C(n_744),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_755),
.A2(n_739),
.B(n_711),
.C(n_678),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_759),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_757),
.A2(n_756),
.B(n_724),
.Y(n_764)
);

NAND4xp25_ASAP7_75t_SL g765 ( 
.A(n_761),
.B(n_742),
.C(n_741),
.D(n_733),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_741),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_758),
.B(n_730),
.Y(n_767)
);

NOR3xp33_ASAP7_75t_L g768 ( 
.A(n_763),
.B(n_760),
.C(n_638),
.Y(n_768)
);

NOR3x1_ASAP7_75t_L g769 ( 
.A(n_766),
.B(n_714),
.C(n_676),
.Y(n_769)
);

OAI211xp5_ASAP7_75t_L g770 ( 
.A1(n_764),
.A2(n_624),
.B(n_681),
.C(n_696),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_769),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_770),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_768),
.Y(n_773)
);

NOR2x1_ASAP7_75t_SL g774 ( 
.A(n_771),
.B(n_765),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_773),
.B(n_767),
.Y(n_775)
);

NAND4xp75_ASAP7_75t_L g776 ( 
.A(n_772),
.B(n_624),
.C(n_631),
.D(n_708),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_771),
.B(n_676),
.Y(n_777)
);

OAI22x1_ASAP7_75t_L g778 ( 
.A1(n_771),
.A2(n_611),
.B1(n_609),
.B2(n_672),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_775),
.B(n_672),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_777),
.Y(n_780)
);

OAI221xp5_ASAP7_75t_L g781 ( 
.A1(n_774),
.A2(n_635),
.B1(n_647),
.B2(n_688),
.C(n_682),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_776),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_782),
.A2(n_690),
.B1(n_696),
.B2(n_688),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_781),
.A2(n_609),
.B(n_611),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_783),
.A2(n_611),
.B1(n_609),
.B2(n_629),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_SL g787 ( 
.A1(n_780),
.A2(n_635),
.B1(n_690),
.B2(n_647),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_784),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_786),
.B(n_779),
.C(n_647),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_789),
.A2(n_779),
.B1(n_785),
.B2(n_703),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_788),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_790),
.B(n_708),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_792),
.A2(n_631),
.B(n_637),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_791),
.A2(n_599),
.B1(n_636),
.B2(n_637),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_795),
.B(n_793),
.C(n_794),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_796),
.B(n_636),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_797),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_697),
.B1(n_681),
.B2(n_653),
.Y(n_799)
);


endmodule