module fake_netlist_6_2500_n_2218 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2218);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2218;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_76),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_41),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_144),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_101),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_35),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_117),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_11),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_23),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_122),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_158),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_145),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_92),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_165),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_53),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_73),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_180),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_68),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_5),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_33),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_17),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_118),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_20),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_134),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_186),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_181),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_156),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_36),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_210),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_164),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_162),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_150),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_170),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_42),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_62),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_31),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_39),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_105),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_143),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_18),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_17),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_69),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_184),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_163),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_212),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_69),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_78),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_3),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_171),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_95),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_121),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_213),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_193),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_124),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_119),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_166),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_192),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_61),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_153),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_91),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_136),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_154),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_49),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_141),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_102),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_24),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_51),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_157),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_224),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_191),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_146),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_215),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_61),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_75),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_148),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_175),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_217),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_203),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_219),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_139),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_57),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_188),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_82),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_168),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_220),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_0),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_89),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_107),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_142),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_209),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_155),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_135),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_194),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_87),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_81),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_182),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_30),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_113),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_225),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_206),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_123),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_55),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_4),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_62),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_25),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_29),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_132),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_37),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_3),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_130),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_199),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_50),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_187),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_201),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_108),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_7),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_38),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_8),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_152),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_1),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_36),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_19),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_38),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_75),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_133),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_77),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_80),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_120),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_131),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_88),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_176),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_70),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_67),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_174),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_71),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_128),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_14),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_204),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_1),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_34),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_106),
.Y(n_396)
);

BUFx2_ASAP7_75t_SL g397 ( 
.A(n_96),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_115),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_68),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_197),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_60),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_99),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_8),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_93),
.Y(n_404)
);

BUFx10_ASAP7_75t_L g405 ( 
.A(n_100),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_66),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_50),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_208),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_5),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_52),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_29),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_159),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_39),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_48),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_63),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_127),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_22),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_60),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_70),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_202),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_55),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_19),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_45),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_140),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_2),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_110),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_97),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_126),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_46),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_207),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_112),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_0),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_47),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_7),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_185),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_116),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_32),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_98),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_84),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_216),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_56),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_33),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_9),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_149),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_24),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_114),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_22),
.Y(n_447)
);

INVxp67_ASAP7_75t_SL g448 ( 
.A(n_231),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_263),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_263),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_335),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_263),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_291),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_263),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_388),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_275),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_438),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_263),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_265),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_266),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_283),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_273),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_283),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_277),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_283),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_234),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_283),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_283),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_228),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_285),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_241),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_234),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_287),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_327),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_292),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_297),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_299),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_327),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_327),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_228),
.Y(n_481)
);

INVxp33_ASAP7_75t_SL g482 ( 
.A(n_238),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_327),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_302),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_315),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_237),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_320),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_238),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_243),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_327),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_340),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_307),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_366),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_366),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_246),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_371),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_240),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_326),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_371),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_340),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_340),
.Y(n_504)
);

BUFx6f_ASAP7_75t_SL g505 ( 
.A(n_282),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_329),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_251),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_340),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_351),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_304),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_308),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_340),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_356),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_305),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_356),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_356),
.Y(n_517)
);

INVxp33_ASAP7_75t_SL g518 ( 
.A(n_240),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_247),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_321),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_356),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_356),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_394),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_226),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_247),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_394),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_409),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_358),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_307),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_409),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_359),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_360),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_233),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_362),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_328),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_274),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_256),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_363),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_380),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_375),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_229),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_377),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_257),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_343),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_268),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_293),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_310),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_317),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_333),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_402),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_349),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_319),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_374),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_376),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_411),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_333),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_380),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_274),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_370),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_333),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_370),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_232),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_564),
.B(n_232),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_457),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_460),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_472),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_449),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_455),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_455),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_492),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_513),
.B(n_342),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_470),
.B(n_481),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_492),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_450),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_450),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_461),
.B(n_463),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_463),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_487),
.B(n_282),
.Y(n_593)
);

OA21x2_ASAP7_75t_L g594 ( 
.A1(n_453),
.A2(n_314),
.B(n_296),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_564),
.B(n_342),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_459),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_459),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_490),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_458),
.B(n_354),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_564),
.B(n_354),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_462),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_452),
.A2(n_262),
.B1(n_410),
.B2(n_261),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_493),
.B(n_254),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_462),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_227),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_464),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_467),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_496),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_512),
.B(n_282),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_466),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_466),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_468),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_468),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_469),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_469),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_465),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_545),
.B(n_296),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_489),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_475),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_471),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_475),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_504),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_509),
.B(n_227),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_514),
.B(n_230),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_479),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_494),
.B(n_314),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_480),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_507),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_480),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_483),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_516),
.B(n_230),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_555),
.Y(n_637)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_491),
.B(n_397),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_R g639 ( 
.A(n_471),
.B(n_365),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_473),
.B(n_259),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_517),
.B(n_522),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_474),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_495),
.B(n_254),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_491),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_521),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_521),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_511),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_534),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_523),
.B(n_524),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_534),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_539),
.B(n_352),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_563),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_474),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_476),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_540),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_540),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_526),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_527),
.B(n_236),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_529),
.B(n_236),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_530),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_533),
.B(n_352),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_640),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_644),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_578),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_578),
.Y(n_667)
);

INVx5_ASAP7_75t_L g668 ( 
.A(n_629),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_584),
.B(n_476),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_591),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_584),
.B(n_596),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_579),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

INVx11_ASAP7_75t_L g676 ( 
.A(n_639),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_610),
.A2(n_556),
.B1(n_477),
.B2(n_484),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_620),
.B(n_426),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_607),
.B(n_482),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_644),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_593),
.B(n_525),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_570),
.A2(n_600),
.B1(n_621),
.B2(n_607),
.Y(n_682)
);

AND3x2_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_372),
.C(n_279),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_576),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_590),
.Y(n_685)
);

INVxp33_ASAP7_75t_L g686 ( 
.A(n_573),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_619),
.B(n_451),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_599),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_605),
.B(n_498),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_579),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_605),
.B(n_518),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_582),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_629),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_586),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_623),
.B(n_477),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_612),
.B(n_478),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_582),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_642),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_644),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_603),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_611),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_575),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_633),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_SL g705 ( 
.A(n_571),
.B(n_286),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_644),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_638),
.B(n_426),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_648),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_629),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_654),
.B(n_478),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_603),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_596),
.B(n_497),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_603),
.Y(n_713)
);

CKINVDCx6p67_ASAP7_75t_R g714 ( 
.A(n_572),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_656),
.B(n_484),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_596),
.B(n_486),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_585),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_585),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_629),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_626),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_604),
.B(n_486),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_589),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_625),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_653),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_626),
.B(n_488),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_588),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_581),
.A2(n_485),
.B1(n_508),
.B2(n_456),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_589),
.B(n_488),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_637),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_625),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_625),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_588),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_592),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_592),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_574),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_592),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_627),
.B(n_499),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_574),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_627),
.B(n_506),
.C(n_499),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_653),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_580),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_577),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_636),
.B(n_506),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_597),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_583),
.B(n_510),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_597),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_577),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_613),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_613),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_613),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_618),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_586),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_636),
.A2(n_288),
.B1(n_260),
.B2(n_387),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_630),
.A2(n_429),
.B1(n_415),
.B2(n_515),
.Y(n_758)
);

BUFx10_ASAP7_75t_L g759 ( 
.A(n_583),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_618),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_660),
.A2(n_531),
.B1(n_535),
.B2(n_510),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_583),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_583),
.B(n_531),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_660),
.B(n_536),
.C(n_535),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_598),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_R g766 ( 
.A(n_643),
.B(n_536),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_586),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_618),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_594),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_643),
.B(n_500),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_661),
.B(n_538),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_661),
.B(n_538),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_622),
.Y(n_773)
);

BUFx4f_ASAP7_75t_L g774 ( 
.A(n_594),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_571),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_638),
.B(n_373),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_598),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_580),
.B(n_544),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_663),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_652),
.A2(n_390),
.B1(n_407),
.B2(n_378),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_653),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_622),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_631),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_544),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_631),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_631),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_SL g788 ( 
.A(n_601),
.B(n_379),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_586),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_659),
.B(n_546),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_652),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_606),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_653),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_580),
.B(n_546),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_606),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_587),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_634),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_637),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_652),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_580),
.B(n_548),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_634),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_608),
.B(n_548),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_608),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_659),
.B(n_505),
.Y(n_804)
);

CKINVDCx6p67_ASAP7_75t_R g805 ( 
.A(n_663),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_663),
.B(n_405),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_614),
.B(n_298),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_587),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_663),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_614),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_537),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_662),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_662),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_641),
.B(n_405),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_617),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_634),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_645),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_645),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_594),
.A2(n_568),
.B(n_393),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_617),
.Y(n_820)
);

BUFx6f_ASAP7_75t_SL g821 ( 
.A(n_624),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_624),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_669),
.B(n_547),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_775),
.B(n_632),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_775),
.B(n_632),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_738),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_671),
.B(n_519),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_664),
.B(n_520),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_738),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_721),
.B(n_647),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_785),
.B(n_647),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_741),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_759),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_679),
.B(n_657),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_726),
.B(n_657),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_776),
.B(n_426),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_779),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_740),
.B(n_587),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_724),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_741),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_771),
.A2(n_444),
.B1(n_550),
.B2(n_541),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_791),
.B(n_333),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_709),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_766),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_772),
.B(n_557),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_724),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_716),
.B(n_528),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_769),
.B(n_426),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_732),
.Y(n_849)
);

INVx4_ASAP7_75t_L g850 ( 
.A(n_779),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_788),
.A2(n_336),
.B1(n_369),
.B2(n_347),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_769),
.B(n_426),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_712),
.B(n_501),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_769),
.B(n_333),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_746),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_682),
.A2(n_567),
.B(n_235),
.C(n_401),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_746),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_665),
.B(n_587),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_759),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_774),
.B(n_333),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_774),
.B(n_333),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_665),
.B(n_587),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_732),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_709),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_747),
.A2(n_422),
.B(n_390),
.C(n_407),
.Y(n_865)
);

BUFx3_ASAP7_75t_L g866 ( 
.A(n_701),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_774),
.B(n_333),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_751),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_712),
.B(n_770),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_680),
.B(n_587),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_680),
.B(n_602),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_699),
.B(n_602),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_699),
.B(n_602),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_706),
.A2(n_594),
.B1(n_393),
.B2(n_383),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_706),
.B(n_602),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_791),
.B(n_602),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_689),
.B(n_454),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_733),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_733),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_751),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_799),
.B(n_602),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_701),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_759),
.B(n_383),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_SL g884 ( 
.A(n_696),
.B(n_262),
.C(n_261),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_799),
.A2(n_245),
.B1(n_249),
.B2(n_244),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_L g886 ( 
.A(n_779),
.B(n_250),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_779),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_691),
.B(n_609),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_805),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_762),
.B(n_258),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_762),
.B(n_809),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_743),
.B(n_505),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_705),
.A2(n_269),
.B1(n_271),
.B2(n_267),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_711),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_762),
.B(n_809),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_713),
.B(n_609),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_749),
.B(n_502),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_815),
.B(n_609),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_764),
.B(n_505),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_763),
.B(n_239),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_723),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_765),
.B(n_609),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_765),
.B(n_609),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_777),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_757),
.A2(n_378),
.B(n_432),
.C(n_425),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_777),
.B(n_609),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_792),
.B(n_615),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_792),
.B(n_615),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_809),
.B(n_270),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_795),
.B(n_615),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_770),
.B(n_543),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_795),
.B(n_615),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_813),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_803),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_803),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_810),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_810),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_811),
.B(n_549),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_820),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_820),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_822),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_822),
.A2(n_424),
.B1(n_301),
.B2(n_312),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_685),
.B(n_272),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_666),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_666),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_812),
.B(n_790),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_778),
.B(n_284),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_794),
.B(n_800),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_811),
.B(n_551),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_761),
.B(n_239),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_709),
.B(n_615),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_745),
.B(n_325),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_720),
.B(n_615),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_813),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_705),
.B(n_395),
.C(n_392),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_720),
.B(n_725),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_720),
.B(n_616),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_808),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_811),
.B(n_337),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_667),
.Y(n_940)
);

NAND3xp33_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_406),
.C(n_399),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_725),
.B(n_616),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_667),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_673),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_811),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_758),
.B(n_553),
.C(n_552),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_744),
.B(n_616),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_782),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_782),
.B(n_338),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_782),
.B(n_344),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_805),
.A2(n_309),
.B1(n_280),
.B2(n_278),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_672),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_722),
.A2(n_311),
.B1(n_276),
.B2(n_281),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_793),
.A2(n_431),
.B1(n_435),
.B2(n_416),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_793),
.B(n_616),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_793),
.B(n_616),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_673),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_685),
.B(n_641),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_674),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_727),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_807),
.B(n_616),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_674),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_735),
.B(n_554),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_767),
.B(n_628),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_675),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_727),
.Y(n_966)
);

AOI22x1_ASAP7_75t_SL g967 ( 
.A1(n_688),
.A2(n_441),
.B1(n_414),
.B2(n_418),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_735),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_729),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_SL g970 ( 
.A1(n_681),
.A2(n_405),
.B1(n_410),
.B2(n_413),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_686),
.B(n_242),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_684),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_675),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_729),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_703),
.B(n_242),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_672),
.B(n_346),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_672),
.B(n_350),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_690),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_677),
.B(n_248),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_672),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_734),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_684),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_683),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_730),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_678),
.A2(n_404),
.B1(n_400),
.B2(n_391),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_678),
.A2(n_389),
.B1(n_386),
.B2(n_364),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_767),
.B(n_789),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_734),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_789),
.B(n_628),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_681),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_681),
.A2(n_568),
.B1(n_445),
.B2(n_443),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_672),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_844),
.B(n_670),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_823),
.B(n_695),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_826),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_952),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_835),
.B(n_806),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_831),
.B(n_681),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_913),
.B(n_670),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_843),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_930),
.A2(n_715),
.B(n_710),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_963),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_834),
.B(n_796),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_826),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_829),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_901),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_913),
.B(n_670),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_843),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_928),
.A2(n_821),
.B1(n_687),
.B2(n_814),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_829),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_832),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_926),
.B(n_796),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_832),
.Y(n_1013)
);

AND2x2_ASAP7_75t_SL g1014 ( 
.A(n_886),
.B(n_707),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_901),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_928),
.A2(n_821),
.B1(n_804),
.B2(n_728),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_843),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_864),
.B(n_838),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_840),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_855),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_848),
.A2(n_717),
.B(n_694),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_857),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_934),
.B(n_676),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_888),
.B(n_904),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_866),
.B(n_702),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_963),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_827),
.B(n_698),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_857),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_836),
.A2(n_781),
.B1(n_707),
.B2(n_737),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_915),
.B(n_796),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_845),
.B(n_676),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_868),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_911),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_968),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_880),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_880),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_916),
.B(n_694),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_874),
.A2(n_821),
.B1(n_714),
.B2(n_819),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_836),
.A2(n_736),
.B1(n_818),
.B2(n_817),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_884),
.A2(n_736),
.B1(n_818),
.B2(n_817),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_864),
.B(n_698),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_971),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_914),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_917),
.B(n_919),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_920),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_921),
.B(n_827),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_848),
.A2(n_750),
.B1(n_816),
.B2(n_737),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_918),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_911),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_869),
.B(n_698),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_972),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_847),
.B(n_714),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

INVx5_ASAP7_75t_L g1054 ( 
.A(n_837),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_846),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_849),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_866),
.B(n_704),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_869),
.B(n_853),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_952),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_864),
.B(n_694),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_824),
.B(n_694),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_825),
.B(n_694),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_863),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_900),
.B(n_717),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_924),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_837),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_878),
.B(n_717),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_852),
.A2(n_961),
.B(n_862),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_925),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_927),
.A2(n_728),
.B1(n_723),
.B2(n_345),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_879),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_882),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_830),
.B(n_717),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_927),
.A2(n_396),
.B1(n_332),
.B2(n_331),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_918),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_889),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_984),
.B(n_688),
.Y(n_1078)
);

BUFx4f_ASAP7_75t_L g1079 ( 
.A(n_983),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_925),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_833),
.B(n_717),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_853),
.B(n_756),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_877),
.B(n_708),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_948),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_894),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_897),
.B(n_756),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_940),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_940),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_897),
.B(n_756),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_943),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_833),
.B(n_859),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_952),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_943),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_944),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_944),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_952),
.Y(n_1096)
);

AO22x1_ASAP7_75t_L g1097 ( 
.A1(n_979),
.A2(n_437),
.B1(n_413),
.B2(n_414),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_890),
.A2(n_330),
.B1(n_385),
.B2(n_384),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_957),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_929),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_828),
.B(n_708),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_958),
.B(n_739),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_837),
.B(n_668),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_957),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_842),
.A2(n_752),
.B1(n_742),
.B2(n_801),
.Y(n_1105)
);

BUFx4f_ASAP7_75t_L g1106 ( 
.A(n_983),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_959),
.Y(n_1107)
);

NAND2x1_ASAP7_75t_L g1108 ( 
.A(n_850),
.B(n_887),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_850),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_859),
.B(n_808),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_850),
.B(n_808),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_972),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_851),
.B(n_418),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_959),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_929),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_890),
.A2(n_322),
.B1(n_361),
.B2(n_355),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_909),
.A2(n_883),
.B1(n_941),
.B2(n_895),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_887),
.B(n_808),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_923),
.Y(n_1119)
);

NOR2xp67_ASAP7_75t_L g1120 ( 
.A(n_892),
.B(n_558),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_975),
.B(n_559),
.Y(n_1121)
);

NAND2x1p5_ASAP7_75t_L g1122 ( 
.A(n_887),
.B(n_889),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_962),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_992),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_992),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_992),
.B(n_808),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_980),
.B(n_742),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_962),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_982),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_965),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_965),
.B(n_748),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_982),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_973),
.B(n_748),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_973),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_841),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_935),
.B(n_421),
.C(n_419),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_992),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_978),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_752),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_938),
.Y(n_1140)
);

NOR2x1p5_ASAP7_75t_L g1141 ( 
.A(n_939),
.B(n_419),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_909),
.A2(n_819),
.B1(n_446),
.B2(n_440),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_858),
.A2(n_871),
.B(n_870),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_938),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_960),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_966),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_854),
.B(n_668),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_967),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_991),
.B(n_753),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_969),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_974),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_981),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_938),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_988),
.B(n_754),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_936),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_902),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_903),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_906),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_872),
.B(n_754),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_907),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_945),
.B(n_421),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_873),
.B(n_755),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_905),
.B(n_434),
.C(n_433),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_875),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_908),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_910),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_842),
.A2(n_801),
.B1(n_797),
.B2(n_787),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_860),
.B(n_668),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_990),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_970),
.B(n_560),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_912),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_939),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_939),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1054),
.A2(n_886),
.B(n_891),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1025),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1051),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1004),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1058),
.A2(n_946),
.B1(n_867),
.B2(n_861),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1048),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1004),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_1140),
.B(n_1144),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_1129),
.B(n_891),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1054),
.A2(n_895),
.B(n_987),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_L g1184 ( 
.A1(n_1018),
.A2(n_867),
.B(n_977),
.C(n_976),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_998),
.B(n_856),
.Y(n_1185)
);

OAI22x1_ASAP7_75t_L g1186 ( 
.A1(n_1083),
.A2(n_899),
.B1(n_893),
.B2(n_953),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1169),
.A2(n_1083),
.B1(n_1006),
.B2(n_1015),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1054),
.A2(n_881),
.B(n_876),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1011),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1054),
.A2(n_964),
.B(n_989),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1002),
.B(n_865),
.Y(n_1191)
);

AO21x1_ASAP7_75t_L g1192 ( 
.A1(n_1018),
.A2(n_977),
.B(n_976),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1034),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_SL g1194 ( 
.A(n_1066),
.B(n_248),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_997),
.A2(n_951),
.B1(n_885),
.B2(n_985),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1026),
.B(n_932),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1046),
.B(n_922),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1042),
.B(n_898),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1001),
.A2(n_949),
.B(n_950),
.C(n_896),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1066),
.A2(n_933),
.B(n_931),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1033),
.B(n_954),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1049),
.B(n_1121),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_994),
.A2(n_932),
.B(n_949),
.C(n_950),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1025),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_996),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1066),
.A2(n_942),
.B(n_937),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1024),
.A2(n_986),
.B1(n_956),
.B2(n_955),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_994),
.B(n_947),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_1068),
.A2(n_755),
.B(n_797),
.C(n_787),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1109),
.A2(n_798),
.B(n_731),
.Y(n_1210)
);

INVx4_ASAP7_75t_L g1211 ( 
.A(n_996),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1013),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_R g1213 ( 
.A(n_1119),
.B(n_252),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1109),
.A2(n_798),
.B(n_731),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1164),
.B(n_760),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1109),
.A2(n_798),
.B(n_731),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_996),
.Y(n_1217)
);

NOR3xp33_ASAP7_75t_SL g1218 ( 
.A(n_1113),
.B(n_434),
.C(n_433),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1144),
.A2(n_637),
.B(n_668),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1020),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1135),
.A2(n_1027),
.B1(n_1115),
.B2(n_1050),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1048),
.A2(n_353),
.B1(n_295),
.B2(n_300),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_L g1223 ( 
.A1(n_1064),
.A2(n_786),
.B(n_784),
.C(n_783),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1164),
.B(n_760),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1009),
.B(n_252),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1044),
.A2(n_1053),
.B1(n_1056),
.B2(n_1055),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_996),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1113),
.A2(n_446),
.B(n_255),
.C(n_264),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1117),
.B(n_768),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1153),
.A2(n_637),
.B(n_668),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_L g1231 ( 
.A(n_1070),
.B(n_650),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1020),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_1122),
.B(n_303),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1057),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1022),
.Y(n_1235)
);

OA22x2_ASAP7_75t_L g1236 ( 
.A1(n_1071),
.A2(n_437),
.B1(n_441),
.B2(n_447),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1156),
.B(n_768),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1157),
.B(n_773),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1112),
.Y(n_1239)
);

OAI21xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1014),
.A2(n_561),
.B(n_562),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1136),
.B(n_253),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1153),
.A2(n_637),
.B(n_693),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1101),
.B(n_442),
.Y(n_1243)
);

O2A1O1Ixp5_ASAP7_75t_L g1244 ( 
.A1(n_1143),
.A2(n_1081),
.B(n_1110),
.C(n_1147),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1158),
.B(n_773),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1038),
.A2(n_786),
.B(n_784),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1022),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1082),
.A2(n_637),
.B(n_693),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1028),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1076),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1160),
.B(n_780),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1165),
.B(n_780),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1014),
.A2(n_442),
.B1(n_447),
.B2(n_253),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1016),
.A2(n_436),
.B(n_264),
.C(n_334),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1086),
.A2(n_693),
.B(n_783),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1089),
.A2(n_693),
.B(n_719),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1101),
.B(n_255),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1028),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1032),
.Y(n_1259)
);

OAI21xp33_ASAP7_75t_L g1260 ( 
.A1(n_1052),
.A2(n_436),
.B(n_334),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_993),
.A2(n_650),
.B(n_719),
.C(n_718),
.Y(n_1261)
);

NAND2xp33_ASAP7_75t_R g1262 ( 
.A(n_1163),
.B(n_339),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1059),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1132),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1061),
.A2(n_700),
.B(n_697),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1166),
.B(n_690),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1172),
.B(n_339),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1171),
.B(n_692),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1172),
.B(n_412),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1172),
.B(n_412),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1045),
.Y(n_1271)
);

AOI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1045),
.A2(n_1155),
.B1(n_1005),
.B2(n_1010),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1012),
.A2(n_428),
.B1(n_420),
.B2(n_427),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1063),
.B(n_692),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1072),
.B(n_697),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_995),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1155),
.B(n_420),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1000),
.B(n_306),
.Y(n_1278)
);

AOI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1081),
.A2(n_1110),
.B(n_1147),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1000),
.B(n_313),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1031),
.A2(n_430),
.B(n_427),
.C(n_428),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1076),
.B(n_542),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1057),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1062),
.A2(n_316),
.B(n_318),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1003),
.B(n_430),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1100),
.B(n_1052),
.Y(n_1286)
);

AO32x1_ASAP7_75t_L g1287 ( 
.A1(n_1142),
.A2(n_542),
.A3(n_565),
.B1(n_566),
.B2(n_569),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1079),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1168),
.A2(n_323),
.B(n_324),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1168),
.A2(n_341),
.B(n_348),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1008),
.A2(n_440),
.B1(n_439),
.B2(n_381),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1100),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1059),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_993),
.A2(n_565),
.B(n_566),
.C(n_569),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1031),
.B(n_439),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1078),
.B(n_367),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1074),
.B(n_368),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1172),
.B(n_382),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1127),
.A2(n_398),
.B(n_408),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1008),
.A2(n_658),
.B1(n_655),
.B2(n_651),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1159),
.A2(n_628),
.B(n_635),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_999),
.A2(n_658),
.B(n_655),
.C(n_651),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1078),
.B(n_635),
.C(n_628),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1077),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1085),
.B(n_651),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1019),
.B(n_645),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1161),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1017),
.A2(n_649),
.B1(n_646),
.B2(n_635),
.Y(n_1309)
);

INVx3_ASAP7_75t_SL g1310 ( 
.A(n_1148),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1035),
.B(n_649),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1036),
.B(n_649),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1170),
.B(n_2),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1162),
.A2(n_635),
.B(n_628),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1043),
.B(n_646),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1120),
.B(n_1070),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1047),
.A2(n_646),
.B(n_635),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1065),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1161),
.B(n_6),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1017),
.A2(n_635),
.B1(n_628),
.B2(n_211),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1077),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1145),
.B(n_6),
.Y(n_1322)
);

OAI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1023),
.A2(n_9),
.B(n_10),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1073),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1059),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1239),
.B(n_1023),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1276),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1209),
.A2(n_1021),
.B(n_1108),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1257),
.A2(n_1141),
.B1(n_1173),
.B2(n_999),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1229),
.A2(n_1041),
.B(n_1091),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1185),
.B(n_1073),
.Y(n_1331)
);

BUFx4f_ASAP7_75t_L g1332 ( 
.A(n_1310),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1185),
.B(n_1097),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1257),
.B(n_1091),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1223),
.A2(n_1118),
.B(n_1111),
.Y(n_1335)
);

OAI21xp33_ASAP7_75t_L g1336 ( 
.A1(n_1243),
.A2(n_1007),
.B(n_1075),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1243),
.B(n_1007),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1223),
.A2(n_1133),
.B(n_1131),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1202),
.B(n_1041),
.Y(n_1339)
);

BUFx4f_ASAP7_75t_L g1340 ( 
.A(n_1310),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1229),
.A2(n_1102),
.B(n_1125),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1174),
.A2(n_1125),
.B(n_1149),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1272),
.A2(n_1139),
.B(n_1030),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1188),
.A2(n_1060),
.B(n_1096),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1208),
.B(n_1146),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1226),
.B(n_1150),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1226),
.B(n_1151),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1190),
.A2(n_1154),
.B(n_1037),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1205),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1183),
.A2(n_1096),
.B(n_1126),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1175),
.B(n_1084),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1205),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_SL g1353 ( 
.A1(n_1192),
.A2(n_1067),
.B(n_1040),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1265),
.A2(n_1167),
.B(n_1105),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1286),
.B(n_1079),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1282),
.B(n_1152),
.Y(n_1356)
);

NOR2xp67_ASAP7_75t_SL g1357 ( 
.A(n_1305),
.B(n_1096),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1319),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1308),
.B(n_1193),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1200),
.A2(n_1167),
.B(n_1105),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1207),
.A2(n_1103),
.B(n_1029),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1205),
.B(n_1092),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1197),
.B(n_1069),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_1213),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1184),
.A2(n_1040),
.B(n_1039),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1199),
.A2(n_1103),
.B(n_1029),
.Y(n_1366)
);

OAI21xp33_ASAP7_75t_L g1367 ( 
.A1(n_1319),
.A2(n_1098),
.B(n_1116),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1179),
.B(n_1087),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1313),
.A2(n_1122),
.B(n_1104),
.C(n_1090),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1308),
.B(n_1313),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1179),
.B(n_1106),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1206),
.A2(n_1093),
.B(n_1069),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1297),
.B(n_1080),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1244),
.A2(n_1107),
.B(n_1093),
.Y(n_1374)
);

BUFx2_ASAP7_75t_R g1375 ( 
.A(n_1176),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_1107),
.B(n_1080),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1180),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1203),
.A2(n_1106),
.B(n_1114),
.C(n_1138),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1184),
.A2(n_1039),
.B(n_1134),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1279),
.A2(n_1123),
.B(n_1134),
.Y(n_1380)
);

AO31x2_ASAP7_75t_L g1381 ( 
.A1(n_1186),
.A2(n_1099),
.A3(n_1095),
.B(n_1088),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1302),
.A2(n_1099),
.B(n_1095),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1250),
.B(n_1094),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1191),
.B(n_1088),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1253),
.A2(n_1130),
.B1(n_1128),
.B2(n_1123),
.C(n_1124),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1250),
.B(n_1092),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1314),
.A2(n_1137),
.B(n_1124),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1293),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1240),
.A2(n_1137),
.B(n_205),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1177),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1178),
.A2(n_200),
.B(n_198),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1213),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1221),
.B(n_10),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1189),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1220),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1178),
.A2(n_189),
.B(n_183),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1233),
.A2(n_177),
.B(n_173),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1235),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1187),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1246),
.A2(n_172),
.B(n_169),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1181),
.A2(n_161),
.B(n_160),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1255),
.A2(n_151),
.B(n_137),
.Y(n_1402)
);

INVx5_ASAP7_75t_L g1403 ( 
.A(n_1205),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1296),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1404)
);

AOI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1195),
.A2(n_15),
.B(n_16),
.Y(n_1405)
);

AOI221x1_ASAP7_75t_L g1406 ( 
.A1(n_1254),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1321),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1211),
.Y(n_1408)
);

AO22x2_ASAP7_75t_L g1409 ( 
.A1(n_1225),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1298),
.A2(n_129),
.B(n_125),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1234),
.B(n_111),
.Y(n_1411)
);

CKINVDCx6p67_ASAP7_75t_R g1412 ( 
.A(n_1264),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1211),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1204),
.Y(n_1414)
);

AOI21xp33_ASAP7_75t_L g1415 ( 
.A1(n_1236),
.A2(n_26),
.B(n_27),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1283),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1293),
.B(n_26),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1256),
.A2(n_94),
.B(n_90),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1212),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1196),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1228),
.A2(n_1281),
.B(n_1260),
.C(n_1322),
.Y(n_1421)
);

BUFx2_ASAP7_75t_R g1422 ( 
.A(n_1324),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1247),
.B(n_27),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1249),
.B(n_28),
.Y(n_1424)
);

NAND2xp33_ASAP7_75t_R g1425 ( 
.A(n_1218),
.B(n_86),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1218),
.B(n_28),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1198),
.B(n_31),
.Y(n_1427)
);

NAND3x1_ASAP7_75t_L g1428 ( 
.A(n_1222),
.B(n_32),
.C(n_34),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1258),
.B(n_35),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1317),
.A2(n_85),
.B(n_83),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1201),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1253),
.B(n_44),
.C(n_45),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1289),
.B(n_47),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1241),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.C(n_53),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1217),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1215),
.A2(n_54),
.B(n_57),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1262),
.B(n_58),
.C(n_59),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1277),
.B(n_58),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1259),
.B(n_59),
.Y(n_1439)
);

INVx5_ASAP7_75t_L g1440 ( 
.A(n_1217),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1262),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1261),
.A2(n_63),
.B(n_64),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_SL g1443 ( 
.A1(n_1320),
.A2(n_64),
.B(n_65),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1236),
.B(n_65),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1304),
.A2(n_74),
.B1(n_67),
.B2(n_72),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1285),
.B(n_66),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1182),
.B(n_72),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1224),
.A2(n_73),
.B(n_74),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1232),
.B(n_1271),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1182),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1182),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1237),
.B(n_1251),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1325),
.Y(n_1453)
);

A2O1A1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1278),
.A2(n_1280),
.B(n_1300),
.C(n_1284),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1248),
.A2(n_1311),
.B(n_1307),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1278),
.A2(n_1280),
.B(n_1291),
.C(n_1290),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1325),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1312),
.A2(n_1315),
.B(n_1245),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1318),
.Y(n_1459)
);

NAND3xp33_ASAP7_75t_L g1460 ( 
.A(n_1273),
.B(n_1295),
.C(n_1292),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1274),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1238),
.B(n_1252),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1227),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1275),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1263),
.A2(n_1268),
.B(n_1266),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1231),
.B(n_1306),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1219),
.A2(n_1242),
.B(n_1230),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1194),
.A2(n_1301),
.B(n_1299),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1316),
.A2(n_1309),
.B(n_1303),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1267),
.B(n_1269),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1287),
.A2(n_1210),
.A3(n_1214),
.B(n_1216),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1472)
);

AOI221x1_ASAP7_75t_L g1473 ( 
.A1(n_1287),
.A2(n_1323),
.B1(n_1319),
.B2(n_1313),
.C(n_1186),
.Y(n_1473)
);

INVx6_ASAP7_75t_SL g1474 ( 
.A(n_1288),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1294),
.A2(n_1184),
.B(n_1244),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1294),
.B(n_1287),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1209),
.A2(n_1223),
.B(n_1272),
.Y(n_1477)
);

INVx5_ASAP7_75t_L g1478 ( 
.A(n_1205),
.Y(n_1478)
);

O2A1O1Ixp5_ASAP7_75t_L g1479 ( 
.A1(n_1257),
.A2(n_836),
.B(n_1243),
.C(n_1296),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1184),
.A2(n_1244),
.B(n_1229),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1209),
.A2(n_1223),
.B(n_1272),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1243),
.A2(n_664),
.B(n_1319),
.C(n_1257),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1229),
.A2(n_1066),
.B(n_1054),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1209),
.A2(n_1223),
.B(n_1272),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1185),
.B(n_1058),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1276),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1184),
.A2(n_1244),
.B(n_1068),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1276),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1286),
.B(n_1002),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1490)
);

AO31x2_ASAP7_75t_L g1491 ( 
.A1(n_1473),
.A2(n_1361),
.A3(n_1366),
.B(n_1378),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1388),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1374),
.A2(n_1376),
.B(n_1477),
.Y(n_1494)
);

NAND2xp33_ASAP7_75t_L g1495 ( 
.A(n_1336),
.B(n_1367),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1457),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1403),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1391),
.A2(n_1396),
.B(n_1487),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1407),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1333),
.B(n_1370),
.Y(n_1500)
);

OA21x2_ASAP7_75t_L g1501 ( 
.A1(n_1481),
.A2(n_1484),
.B(n_1487),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1407),
.Y(n_1502)
);

AO32x2_ASAP7_75t_L g1503 ( 
.A1(n_1450),
.A2(n_1406),
.A3(n_1405),
.B1(n_1445),
.B2(n_1385),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_L g1504 ( 
.A(n_1403),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1337),
.B(n_1334),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1367),
.B(n_1336),
.C(n_1437),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1327),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1419),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1451),
.B(n_1355),
.Y(n_1509)
);

BUFx12f_ASAP7_75t_L g1510 ( 
.A(n_1407),
.Y(n_1510)
);

CKINVDCx11_ASAP7_75t_R g1511 ( 
.A(n_1364),
.Y(n_1511)
);

AO21x1_ASAP7_75t_L g1512 ( 
.A1(n_1391),
.A2(n_1442),
.B(n_1405),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1403),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_SL g1514 ( 
.A1(n_1442),
.A2(n_1347),
.B(n_1346),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1372),
.A2(n_1342),
.B(n_1343),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1416),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1357),
.B(n_1478),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1485),
.A2(n_1389),
.B(n_1475),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1455),
.A2(n_1387),
.B(n_1380),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1432),
.A2(n_1415),
.B1(n_1409),
.B2(n_1437),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1389),
.A2(n_1465),
.B(n_1341),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1353),
.A2(n_1379),
.B(n_1400),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1348),
.A2(n_1350),
.B(n_1344),
.Y(n_1523)
);

AOI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1432),
.A2(n_1415),
.B1(n_1431),
.B2(n_1434),
.C(n_1409),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_SL g1525 ( 
.A(n_1346),
.B(n_1347),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1331),
.B(n_1384),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1427),
.B(n_1421),
.C(n_1329),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1453),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1420),
.B(n_1489),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1420),
.B(n_1444),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1335),
.A2(n_1379),
.B(n_1338),
.Y(n_1531)
);

OAI222xp33_ASAP7_75t_L g1532 ( 
.A1(n_1393),
.A2(n_1448),
.B1(n_1436),
.B2(n_1438),
.C1(n_1345),
.C2(n_1446),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1358),
.B(n_1417),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1445),
.A2(n_1358),
.B1(n_1426),
.B2(n_1460),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1371),
.Y(n_1535)
);

INVx8_ASAP7_75t_L g1536 ( 
.A(n_1478),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1412),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_SL g1538 ( 
.A1(n_1369),
.A2(n_1443),
.B(n_1345),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1399),
.A2(n_1441),
.B1(n_1447),
.B2(n_1470),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1488),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1478),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1363),
.B(n_1461),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1375),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1414),
.B(n_1326),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1332),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1483),
.A2(n_1454),
.B(n_1360),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_L g1548 ( 
.A(n_1425),
.B(n_1404),
.C(n_1402),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1363),
.B(n_1464),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1354),
.A2(n_1330),
.B(n_1468),
.Y(n_1550)
);

OA21x2_ASAP7_75t_L g1551 ( 
.A1(n_1402),
.A2(n_1418),
.B(n_1476),
.Y(n_1551)
);

AO221x2_ASAP7_75t_L g1552 ( 
.A1(n_1418),
.A2(n_1428),
.B1(n_1460),
.B2(n_1339),
.C(n_1424),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1459),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1480),
.A2(n_1430),
.B(n_1458),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1362),
.Y(n_1555)
);

BUFx4f_ASAP7_75t_L g1556 ( 
.A(n_1435),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1368),
.B(n_1356),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1377),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1452),
.B(n_1462),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1332),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1373),
.A2(n_1451),
.B1(n_1429),
.B2(n_1424),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1394),
.Y(n_1562)
);

AO21x2_ASAP7_75t_L g1563 ( 
.A1(n_1456),
.A2(n_1469),
.B(n_1466),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1386),
.B(n_1457),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_R g1565 ( 
.A(n_1392),
.B(n_1451),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1395),
.B(n_1398),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1383),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1449),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1480),
.A2(n_1430),
.B(n_1458),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1365),
.A2(n_1397),
.B(n_1423),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1410),
.A2(n_1429),
.B(n_1423),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1439),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1381),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1401),
.A2(n_1439),
.B(n_1472),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1351),
.A2(n_1411),
.B(n_1471),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1381),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1381),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1359),
.A2(n_1433),
.B1(n_1351),
.B2(n_1340),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1413),
.A2(n_1471),
.B(n_1362),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1411),
.A2(n_1413),
.B(n_1422),
.C(n_1474),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1362),
.A2(n_1463),
.B(n_1440),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1408),
.B(n_1435),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1349),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1349),
.Y(n_1584)
);

AOI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1440),
.A2(n_1474),
.B(n_1352),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1440),
.A2(n_1352),
.B(n_1408),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1337),
.A2(n_1083),
.B1(n_828),
.B2(n_1101),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1388),
.Y(n_1589)
);

OR2x6_ASAP7_75t_L g1590 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1327),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1487),
.A2(n_1361),
.B(n_1475),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1435),
.Y(n_1594)
);

INVx4_ASAP7_75t_L g1595 ( 
.A(n_1440),
.Y(n_1595)
);

CKINVDCx16_ASAP7_75t_R g1596 ( 
.A(n_1364),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1485),
.B(n_1331),
.Y(n_1598)
);

OAI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1599)
);

AO21x2_ASAP7_75t_L g1600 ( 
.A1(n_1487),
.A2(n_1361),
.B(n_1475),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1391),
.B(n_1396),
.Y(n_1601)
);

A2O1A1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1482),
.A2(n_1396),
.B(n_1391),
.C(n_1319),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1482),
.A2(n_1243),
.B1(n_1319),
.B2(n_1405),
.C(n_1313),
.Y(n_1603)
);

BUFx8_ASAP7_75t_L g1604 ( 
.A(n_1407),
.Y(n_1604)
);

AND2x6_ASAP7_75t_L g1605 ( 
.A(n_1346),
.B(n_1347),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1388),
.Y(n_1606)
);

BUFx10_ASAP7_75t_L g1607 ( 
.A(n_1359),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1608)
);

NAND2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1357),
.B(n_1403),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1327),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1364),
.Y(n_1611)
);

BUFx4_ASAP7_75t_SL g1612 ( 
.A(n_1453),
.Y(n_1612)
);

AOI22x1_ASAP7_75t_L g1613 ( 
.A1(n_1391),
.A2(n_1186),
.B1(n_1396),
.B2(n_1442),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1403),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1477),
.A2(n_1484),
.B(n_1481),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1617)
);

O2A1O1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1482),
.A2(n_1243),
.B(n_1319),
.C(n_1405),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1619)
);

CKINVDCx8_ASAP7_75t_R g1620 ( 
.A(n_1364),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1390),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1432),
.A2(n_1313),
.B1(n_1482),
.B2(n_1257),
.Y(n_1624)
);

AO21x2_ASAP7_75t_L g1625 ( 
.A1(n_1487),
.A2(n_1361),
.B(n_1475),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1450),
.B(n_1451),
.Y(n_1626)
);

INVx5_ASAP7_75t_L g1627 ( 
.A(n_1362),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1477),
.A2(n_1484),
.B(n_1481),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1327),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1489),
.B(n_1027),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1453),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1453),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1407),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1432),
.A2(n_1319),
.B1(n_1313),
.B2(n_1405),
.Y(n_1634)
);

AOI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1366),
.A2(n_1361),
.B(n_1229),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1327),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1332),
.Y(n_1637)
);

A2O1A1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1482),
.A2(n_1396),
.B(n_1391),
.C(n_1319),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1328),
.A2(n_1467),
.B(n_1382),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_SL g1642 ( 
.A1(n_1391),
.A2(n_1396),
.B(n_1442),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1432),
.A2(n_1319),
.B1(n_1313),
.B2(n_1405),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1479),
.A2(n_1482),
.B(n_1396),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1432),
.A2(n_1319),
.B1(n_1313),
.B2(n_1405),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1485),
.B(n_1331),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1337),
.A2(n_1083),
.B1(n_828),
.B2(n_1101),
.Y(n_1647)
);

AO32x2_ASAP7_75t_L g1648 ( 
.A1(n_1450),
.A2(n_1406),
.A3(n_1473),
.B1(n_1273),
.B2(n_1405),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1366),
.A2(n_1361),
.B(n_1391),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1327),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1375),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1432),
.A2(n_1370),
.B1(n_1333),
.B2(n_1406),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1370),
.B(n_1420),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1388),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1541),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1588),
.A2(n_1601),
.B1(n_1590),
.B2(n_1587),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_SL g1659 ( 
.A1(n_1602),
.A2(n_1638),
.B(n_1590),
.Y(n_1659)
);

CKINVDCx14_ASAP7_75t_R g1660 ( 
.A(n_1511),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1611),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1496),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1507),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1533),
.B(n_1567),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1535),
.B(n_1505),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1588),
.A2(n_1590),
.B1(n_1601),
.B2(n_1647),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1511),
.Y(n_1667)
);

AOI21x1_ASAP7_75t_SL g1668 ( 
.A1(n_1598),
.A2(n_1646),
.B(n_1526),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1505),
.B(n_1598),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1500),
.B(n_1509),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1618),
.A2(n_1638),
.B(n_1602),
.C(n_1603),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1529),
.B(n_1622),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1499),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1498),
.A2(n_1601),
.B(n_1588),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1554),
.A2(n_1569),
.B(n_1521),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1500),
.B(n_1557),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1651),
.B(n_1654),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1534),
.B(n_1539),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1564),
.B(n_1496),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1534),
.B(n_1578),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1578),
.B(n_1508),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1605),
.B(n_1543),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1633),
.B(n_1581),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1605),
.B(n_1543),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1634),
.A2(n_1643),
.B1(n_1645),
.B2(n_1603),
.Y(n_1685)
);

OA22x2_ASAP7_75t_L g1686 ( 
.A1(n_1624),
.A2(n_1642),
.B1(n_1644),
.B2(n_1490),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1493),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1624),
.A2(n_1618),
.B(n_1498),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_SL g1689 ( 
.A1(n_1517),
.A2(n_1609),
.B(n_1559),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1690)
);

BUFx4f_ASAP7_75t_SL g1691 ( 
.A(n_1510),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1493),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1605),
.B(n_1572),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1581),
.B(n_1502),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1525),
.B(n_1653),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1634),
.A2(n_1643),
.B1(n_1645),
.B2(n_1520),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1506),
.A2(n_1527),
.B1(n_1524),
.B2(n_1653),
.C(n_1520),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1623),
.B(n_1552),
.Y(n_1699)
);

O2A1O1Ixp5_ASAP7_75t_L g1700 ( 
.A1(n_1512),
.A2(n_1608),
.B(n_1621),
.C(n_1639),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1589),
.B(n_1606),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1613),
.A2(n_1524),
.B1(n_1649),
.B2(n_1548),
.Y(n_1702)
);

OA22x2_ASAP7_75t_L g1703 ( 
.A1(n_1599),
.A2(n_1644),
.B1(n_1640),
.B2(n_1621),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1552),
.B(n_1568),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1640),
.A2(n_1627),
.B1(n_1555),
.B2(n_1655),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_SL g1706 ( 
.A1(n_1571),
.A2(n_1521),
.B(n_1518),
.C(n_1582),
.Y(n_1706)
);

OA21x2_ASAP7_75t_L g1707 ( 
.A1(n_1494),
.A2(n_1550),
.B(n_1547),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1555),
.A2(n_1627),
.B1(n_1655),
.B2(n_1591),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1607),
.B(n_1528),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1561),
.B(n_1518),
.Y(n_1711)
);

AOI21x1_ASAP7_75t_SL g1712 ( 
.A1(n_1566),
.A2(n_1648),
.B(n_1503),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1553),
.B(n_1631),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1632),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1540),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1563),
.A2(n_1547),
.B(n_1571),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1515),
.A2(n_1519),
.B(n_1492),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1563),
.A2(n_1600),
.B(n_1592),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1558),
.B(n_1562),
.Y(n_1719)
);

O2A1O1Ixp5_ASAP7_75t_L g1720 ( 
.A1(n_1532),
.A2(n_1635),
.B(n_1575),
.C(n_1570),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1594),
.B(n_1545),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1555),
.A2(n_1627),
.B1(n_1629),
.B2(n_1650),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1555),
.A2(n_1627),
.B1(n_1636),
.B2(n_1610),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1532),
.A2(n_1538),
.B1(n_1522),
.B2(n_1580),
.C(n_1592),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1607),
.B(n_1583),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1544),
.B(n_1652),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1600),
.A2(n_1625),
.B(n_1523),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1517),
.A2(n_1609),
.B(n_1580),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1593),
.A2(n_1597),
.B(n_1641),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1576),
.Y(n_1730)
);

O2A1O1Ixp5_ASAP7_75t_L g1731 ( 
.A1(n_1595),
.A2(n_1577),
.B(n_1573),
.C(n_1582),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1560),
.A2(n_1537),
.B(n_1551),
.C(n_1516),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1584),
.B(n_1596),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1556),
.B(n_1585),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1491),
.B(n_1574),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1497),
.B(n_1513),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1565),
.A2(n_1504),
.B(n_1497),
.Y(n_1737)
);

NOR2xp67_ASAP7_75t_L g1738 ( 
.A(n_1546),
.B(n_1637),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1504),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1504),
.B(n_1614),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1513),
.B(n_1614),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1604),
.B(n_1614),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1513),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1491),
.B(n_1579),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1503),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1536),
.A2(n_1586),
.B(n_1648),
.C(n_1542),
.Y(n_1746)
);

AOI21x1_ASAP7_75t_SL g1747 ( 
.A1(n_1612),
.A2(n_1620),
.B(n_1604),
.Y(n_1747)
);

INVxp67_ASAP7_75t_L g1748 ( 
.A(n_1542),
.Y(n_1748)
);

OR2x6_ASAP7_75t_L g1749 ( 
.A(n_1542),
.B(n_1615),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1501),
.B(n_1531),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1542),
.B(n_1616),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1617),
.B(n_1619),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1628),
.A2(n_1569),
.B(n_1554),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1529),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1618),
.A2(n_1482),
.B(n_1638),
.C(n_1602),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1604),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1602),
.A2(n_1396),
.B(n_1391),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1588),
.A2(n_1601),
.B1(n_1590),
.B2(n_1587),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1587),
.B(n_1647),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1505),
.B(n_1500),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_SL g1763 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1763)
);

O2A1O1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1602),
.A2(n_1482),
.B(n_1638),
.C(n_1624),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1529),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1498),
.A2(n_1590),
.B(n_1588),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1505),
.B(n_1598),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1507),
.Y(n_1768)
);

O2A1O1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1602),
.A2(n_1482),
.B(n_1638),
.C(n_1624),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1505),
.B(n_1598),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1529),
.B(n_1622),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1588),
.A2(n_1601),
.B1(n_1590),
.B2(n_1587),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1529),
.B(n_1622),
.Y(n_1774)
);

AND2x2_ASAP7_75t_SL g1775 ( 
.A(n_1495),
.B(n_1634),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1507),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1604),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_SL g1778 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1778)
);

INVx3_ASAP7_75t_SL g1779 ( 
.A(n_1546),
.Y(n_1779)
);

O2A1O1Ixp5_ASAP7_75t_L g1780 ( 
.A1(n_1512),
.A2(n_1638),
.B(n_1602),
.C(n_1599),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1602),
.A2(n_1482),
.B(n_1638),
.C(n_1624),
.Y(n_1782)
);

INVx6_ASAP7_75t_L g1783 ( 
.A(n_1604),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1530),
.B(n_1630),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1498),
.A2(n_1590),
.B(n_1588),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1505),
.B(n_1598),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1683),
.Y(n_1788)
);

OR2x6_ASAP7_75t_L g1789 ( 
.A(n_1757),
.B(n_1659),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1715),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1730),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1753),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1689),
.B(n_1688),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1749),
.B(n_1763),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1704),
.B(n_1699),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1663),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1674),
.B(n_1766),
.Y(n_1797)
);

AO21x2_ASAP7_75t_L g1798 ( 
.A1(n_1716),
.A2(n_1727),
.B(n_1671),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1669),
.Y(n_1799)
);

NAND4xp25_ASAP7_75t_L g1800 ( 
.A(n_1698),
.B(n_1782),
.C(n_1769),
.D(n_1764),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1683),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_L g1802 ( 
.A(n_1728),
.B(n_1732),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1662),
.Y(n_1803)
);

AO21x2_ASAP7_75t_L g1804 ( 
.A1(n_1718),
.A2(n_1755),
.B(n_1702),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_SL g1805 ( 
.A(n_1705),
.B(n_1722),
.Y(n_1805)
);

AO21x2_ASAP7_75t_L g1806 ( 
.A1(n_1702),
.A2(n_1786),
.B(n_1750),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1696),
.B(n_1746),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1682),
.B(n_1684),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1768),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1751),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1751),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1682),
.B(n_1684),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1776),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1687),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1690),
.B(n_1693),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1775),
.A2(n_1685),
.B1(n_1697),
.B2(n_1759),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1690),
.B(n_1693),
.Y(n_1817)
);

AO21x2_ASAP7_75t_L g1818 ( 
.A1(n_1735),
.A2(n_1696),
.B(n_1685),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1694),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1729),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1687),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1749),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1719),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1749),
.B(n_1778),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1752),
.B(n_1695),
.Y(n_1825)
);

OA21x2_ASAP7_75t_L g1826 ( 
.A1(n_1720),
.A2(n_1700),
.B(n_1780),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1745),
.B(n_1703),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1703),
.B(n_1686),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1701),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1719),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1669),
.B(n_1767),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1709),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_SL g1833 ( 
.A(n_1767),
.B(n_1770),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1711),
.B(n_1709),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1692),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1657),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1679),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1711),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1686),
.Y(n_1839)
);

AO21x2_ASAP7_75t_L g1840 ( 
.A1(n_1705),
.A2(n_1706),
.B(n_1658),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1744),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1787),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1676),
.B(n_1658),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1675),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1677),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1731),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1754),
.B(n_1765),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1672),
.Y(n_1848)
);

AO21x2_ASAP7_75t_L g1849 ( 
.A1(n_1666),
.A2(n_1772),
.B(n_1758),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1717),
.Y(n_1850)
);

INVx1_ASAP7_75t_SL g1851 ( 
.A(n_1714),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1666),
.A2(n_1772),
.B(n_1758),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1708),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1752),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1771),
.B(n_1774),
.Y(n_1855)
);

AO21x2_ASAP7_75t_L g1856 ( 
.A1(n_1697),
.A2(n_1722),
.B(n_1723),
.Y(n_1856)
);

NAND2x1p5_ASAP7_75t_L g1857 ( 
.A(n_1707),
.B(n_1734),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1723),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1665),
.B(n_1680),
.Y(n_1859)
);

OA21x2_ASAP7_75t_L g1860 ( 
.A1(n_1724),
.A2(n_1708),
.B(n_1681),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1670),
.B(n_1656),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1664),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1717),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1760),
.B(n_1781),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1726),
.B(n_1710),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1713),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1743),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1791),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1791),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1792),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1800),
.A2(n_1678),
.B1(n_1785),
.B2(n_1761),
.C(n_1773),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1816),
.A2(n_1784),
.B1(n_1660),
.B2(n_1733),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1810),
.B(n_1725),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1857),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1792),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1792),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1838),
.B(n_1832),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1838),
.B(n_1712),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1796),
.Y(n_1879)
);

INVx4_ASAP7_75t_L g1880 ( 
.A(n_1789),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1810),
.B(n_1673),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1815),
.B(n_1740),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1789),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1832),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1820),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1815),
.B(n_1817),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1811),
.B(n_1806),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1811),
.Y(n_1888)
);

NAND2x1p5_ASAP7_75t_L g1889 ( 
.A(n_1793),
.B(n_1739),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1817),
.B(n_1741),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1812),
.B(n_1673),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1806),
.B(n_1748),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1834),
.B(n_1833),
.Y(n_1893)
);

INVxp67_ASAP7_75t_L g1894 ( 
.A(n_1819),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1808),
.B(n_1739),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_1857),
.Y(n_1896)
);

BUFx3_ASAP7_75t_L g1897 ( 
.A(n_1794),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1854),
.B(n_1736),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1819),
.B(n_1721),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1806),
.B(n_1742),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1868),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1871),
.A2(n_1789),
.B1(n_1793),
.B2(n_1849),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1897),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1871),
.A2(n_1789),
.B1(n_1849),
.B2(n_1804),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1868),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1893),
.B(n_1865),
.Y(n_1906)
);

AOI21xp33_ASAP7_75t_L g1907 ( 
.A1(n_1900),
.A2(n_1804),
.B(n_1807),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1893),
.B(n_1834),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1897),
.B(n_1794),
.Y(n_1909)
);

OAI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1872),
.A2(n_1802),
.B1(n_1852),
.B2(n_1839),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1897),
.B(n_1794),
.Y(n_1911)
);

OAI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1872),
.A2(n_1802),
.B1(n_1797),
.B2(n_1839),
.C(n_1828),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1880),
.A2(n_1849),
.B1(n_1828),
.B2(n_1840),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1869),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1898),
.B(n_1794),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1886),
.B(n_1827),
.Y(n_1916)
);

OR2x2_ASAP7_75t_SL g1917 ( 
.A(n_1900),
.B(n_1826),
.Y(n_1917)
);

CKINVDCx16_ASAP7_75t_R g1918 ( 
.A(n_1882),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1878),
.A2(n_1831),
.B1(n_1799),
.B2(n_1846),
.C(n_1845),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1869),
.Y(n_1920)
);

AOI33xp33_ASAP7_75t_L g1921 ( 
.A1(n_1888),
.A2(n_1827),
.A3(n_1846),
.B1(n_1851),
.B2(n_1859),
.B3(n_1866),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1884),
.Y(n_1922)
);

INVx5_ASAP7_75t_L g1923 ( 
.A(n_1880),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1889),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1899),
.B(n_1855),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1888),
.B(n_1818),
.Y(n_1926)
);

OAI211xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1899),
.A2(n_1842),
.B(n_1847),
.C(n_1866),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1886),
.B(n_1837),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1870),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1870),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1886),
.B(n_1825),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1879),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1880),
.A2(n_1840),
.B1(n_1797),
.B2(n_1856),
.Y(n_1933)
);

OAI221xp5_ASAP7_75t_SL g1934 ( 
.A1(n_1887),
.A2(n_1797),
.B1(n_1853),
.B2(n_1843),
.C(n_1855),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1882),
.B(n_1825),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1870),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1891),
.B(n_1848),
.Y(n_1937)
);

OA332x1_ASAP7_75t_L g1938 ( 
.A1(n_1878),
.A2(n_1818),
.A3(n_1747),
.B1(n_1859),
.B2(n_1667),
.B3(n_1668),
.C1(n_1840),
.C2(n_1795),
.Y(n_1938)
);

OA21x2_ASAP7_75t_L g1939 ( 
.A1(n_1875),
.A2(n_1844),
.B(n_1863),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1884),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1887),
.B(n_1818),
.Y(n_1941)
);

OR2x6_ASAP7_75t_L g1942 ( 
.A(n_1880),
.B(n_1797),
.Y(n_1942)
);

AND2x4_ASAP7_75t_L g1943 ( 
.A(n_1898),
.B(n_1824),
.Y(n_1943)
);

AO21x2_ASAP7_75t_L g1944 ( 
.A1(n_1885),
.A2(n_1850),
.B(n_1844),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1880),
.A2(n_1797),
.B1(n_1856),
.B2(n_1843),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1877),
.A2(n_1795),
.B1(n_1803),
.B2(n_1814),
.C(n_1821),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1894),
.A2(n_1853),
.B1(n_1858),
.B2(n_1841),
.C(n_1830),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1883),
.A2(n_1856),
.B1(n_1860),
.B2(n_1824),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1873),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1881),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1876),
.Y(n_1951)
);

OAI33xp33_ASAP7_75t_L g1952 ( 
.A1(n_1877),
.A2(n_1830),
.A3(n_1823),
.B1(n_1841),
.B2(n_1809),
.B3(n_1813),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1889),
.A2(n_1801),
.B1(n_1788),
.B2(n_1783),
.Y(n_1953)
);

AOI222xp33_ASAP7_75t_L g1954 ( 
.A1(n_1894),
.A2(n_1805),
.B1(n_1864),
.B2(n_1861),
.C1(n_1858),
.C2(n_1862),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1883),
.A2(n_1798),
.B1(n_1860),
.B2(n_1801),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1882),
.B(n_1825),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1879),
.Y(n_1957)
);

INVxp67_ASAP7_75t_SL g1958 ( 
.A(n_1887),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1889),
.A2(n_1829),
.B1(n_1790),
.B2(n_1822),
.C(n_1835),
.Y(n_1959)
);

OR2x6_ASAP7_75t_L g1960 ( 
.A(n_1942),
.B(n_1883),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1939),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1901),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1905),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1918),
.B(n_1890),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1906),
.B(n_1779),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1914),
.Y(n_1966)
);

BUFx12f_ASAP7_75t_L g1967 ( 
.A(n_1924),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1920),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1923),
.B(n_1874),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1919),
.B(n_1883),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1932),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1939),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_SL g1973 ( 
.A(n_1904),
.B(n_1874),
.C(n_1896),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1957),
.Y(n_1974)
);

AND4x1_ASAP7_75t_L g1975 ( 
.A(n_1902),
.B(n_1913),
.C(n_1921),
.D(n_1933),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1909),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1908),
.B(n_1661),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1922),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1915),
.B(n_1890),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1944),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1944),
.Y(n_1981)
);

INVx4_ASAP7_75t_SL g1982 ( 
.A(n_1924),
.Y(n_1982)
);

AND2x4_ASAP7_75t_L g1983 ( 
.A(n_1923),
.B(n_1874),
.Y(n_1983)
);

OA21x2_ASAP7_75t_L g1984 ( 
.A1(n_1907),
.A2(n_1947),
.B(n_1948),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1926),
.B(n_1873),
.Y(n_1985)
);

NOR3xp33_ASAP7_75t_SL g1986 ( 
.A(n_1912),
.B(n_1867),
.C(n_1836),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1940),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1949),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1915),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1923),
.B(n_1896),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1944),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1929),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1930),
.Y(n_1993)
);

INVx11_ASAP7_75t_L g1994 ( 
.A(n_1938),
.Y(n_1994)
);

BUFx8_ASAP7_75t_L g1995 ( 
.A(n_1924),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1950),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1936),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1925),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1923),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1951),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1950),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1946),
.B(n_1895),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1962),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1962),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1989),
.B(n_1915),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1989),
.B(n_1943),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1979),
.B(n_1976),
.Y(n_2007)
);

NOR3xp33_ASAP7_75t_L g2008 ( 
.A(n_1973),
.B(n_1910),
.C(n_1934),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1976),
.B(n_1943),
.Y(n_2009)
);

AOI33xp33_ASAP7_75t_L g2010 ( 
.A1(n_1975),
.A2(n_1955),
.A3(n_1945),
.B1(n_1829),
.B2(n_1938),
.B3(n_1864),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1964),
.B(n_1909),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1995),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1964),
.B(n_1909),
.Y(n_2013)
);

NAND2xp33_ASAP7_75t_SL g2014 ( 
.A(n_1986),
.B(n_1921),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1963),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1980),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1970),
.A2(n_1952),
.B(n_1927),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1975),
.B(n_1954),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1987),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1980),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1963),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1998),
.B(n_1937),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1966),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1985),
.B(n_1941),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1999),
.B(n_1953),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1978),
.B(n_1931),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1985),
.B(n_1941),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1988),
.B(n_1917),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1982),
.B(n_1911),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1966),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1999),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1978),
.B(n_1931),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1968),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1988),
.B(n_1917),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2002),
.B(n_1916),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1968),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_1995),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1971),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1984),
.B(n_1935),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1971),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1996),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1974),
.Y(n_2042)
);

NAND2xp33_ASAP7_75t_SL g2043 ( 
.A(n_1999),
.B(n_1924),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_2001),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1999),
.Y(n_2045)
);

OAI322xp33_ASAP7_75t_L g2046 ( 
.A1(n_1994),
.A2(n_1958),
.A3(n_1974),
.B1(n_1959),
.B2(n_1977),
.C1(n_1892),
.C2(n_1993),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1997),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1994),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1980),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1984),
.B(n_1935),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1982),
.B(n_1903),
.Y(n_2051)
);

NOR3xp33_ASAP7_75t_SL g2052 ( 
.A(n_1965),
.B(n_1867),
.C(n_1928),
.Y(n_2052)
);

OAI21xp33_ASAP7_75t_L g2053 ( 
.A1(n_1960),
.A2(n_1892),
.B(n_1942),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1995),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1984),
.B(n_1873),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1967),
.B(n_1691),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_2008),
.B(n_1999),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2029),
.B(n_1982),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2016),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2017),
.B(n_1984),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2018),
.B(n_1992),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2003),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2029),
.B(n_1982),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2016),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2003),
.Y(n_2065)
);

OAI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_2048),
.A2(n_1999),
.B1(n_1923),
.B2(n_1942),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2011),
.B(n_1982),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2020),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2019),
.B(n_1992),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2004),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_2010),
.B(n_1924),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2004),
.Y(n_2072)
);

AND2x4_ASAP7_75t_L g2073 ( 
.A(n_2051),
.B(n_1960),
.Y(n_2073)
);

CKINVDCx16_ASAP7_75t_R g2074 ( 
.A(n_2012),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2020),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2015),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2015),
.Y(n_2077)
);

AOI21xp33_ASAP7_75t_SL g2078 ( 
.A1(n_2056),
.A2(n_1756),
.B(n_1960),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2022),
.B(n_1956),
.Y(n_2079)
);

NOR2x1_ASAP7_75t_L g2080 ( 
.A(n_2031),
.B(n_1969),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2052),
.B(n_2014),
.Y(n_2081)
);

OAI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2055),
.A2(n_1942),
.B1(n_1960),
.B2(n_1883),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_2031),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2049),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_2043),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_2041),
.Y(n_2086)
);

NOR4xp25_ASAP7_75t_L g2087 ( 
.A(n_2046),
.B(n_1980),
.C(n_1961),
.D(n_1972),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2012),
.B(n_2037),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2035),
.B(n_2000),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2011),
.B(n_1969),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_SL g2091 ( 
.A(n_2046),
.B(n_1967),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_2037),
.B(n_1777),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2044),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2049),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2013),
.B(n_1969),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_2051),
.B(n_1960),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2013),
.B(n_1969),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2086),
.B(n_2054),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_2085),
.Y(n_2099)
);

INVx1_ASAP7_75t_SL g2100 ( 
.A(n_2085),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2080),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2093),
.B(n_2081),
.Y(n_2102)
);

AOI22xp33_ASAP7_75t_L g2103 ( 
.A1(n_2091),
.A2(n_2053),
.B1(n_2025),
.B2(n_2039),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2062),
.Y(n_2104)
);

NAND2x1_ASAP7_75t_SL g2105 ( 
.A(n_2080),
.B(n_2031),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2062),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_2083),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2074),
.B(n_2054),
.Y(n_2108)
);

AO21x2_ASAP7_75t_L g2109 ( 
.A1(n_2060),
.A2(n_2055),
.B(n_2034),
.Y(n_2109)
);

INVx1_ASAP7_75t_SL g2110 ( 
.A(n_2058),
.Y(n_2110)
);

AND2x4_ASAP7_75t_L g2111 ( 
.A(n_2058),
.B(n_2045),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2063),
.B(n_2067),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_2063),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_2091),
.A2(n_2053),
.B1(n_2050),
.B2(n_1798),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2067),
.B(n_2007),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2090),
.B(n_2007),
.Y(n_2116)
);

INVxp67_ASAP7_75t_L g2117 ( 
.A(n_2057),
.Y(n_2117)
);

NAND3xp33_ASAP7_75t_L g2118 ( 
.A(n_2060),
.B(n_2045),
.C(n_2034),
.Y(n_2118)
);

NAND4xp75_ASAP7_75t_L g2119 ( 
.A(n_2061),
.B(n_1738),
.C(n_2005),
.D(n_2006),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_2071),
.A2(n_1798),
.B1(n_2045),
.B2(n_2006),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_SL g2121 ( 
.A1(n_2061),
.A2(n_2005),
.B1(n_2028),
.B2(n_2009),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_2073),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2069),
.B(n_2028),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2065),
.Y(n_2124)
);

NAND3x1_ASAP7_75t_SL g2125 ( 
.A(n_2074),
.B(n_2087),
.C(n_1783),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2073),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2065),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2099),
.B(n_2088),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2103),
.A2(n_2096),
.B1(n_2073),
.B2(n_2087),
.Y(n_2129)
);

OAI21xp5_ASAP7_75t_SL g2130 ( 
.A1(n_2114),
.A2(n_2078),
.B(n_2066),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2100),
.B(n_2110),
.Y(n_2131)
);

OAI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2118),
.A2(n_2078),
.B(n_2082),
.Y(n_2132)
);

AOI222xp33_ASAP7_75t_L g2133 ( 
.A1(n_2117),
.A2(n_2073),
.B1(n_2096),
.B2(n_2069),
.C1(n_2083),
.C2(n_2077),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2107),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2113),
.B(n_2079),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2112),
.B(n_2090),
.Y(n_2136)
);

NAND3xp33_ASAP7_75t_L g2137 ( 
.A(n_2102),
.B(n_2072),
.C(n_2070),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2112),
.B(n_2095),
.Y(n_2138)
);

AO22x1_ASAP7_75t_L g2139 ( 
.A1(n_2125),
.A2(n_2096),
.B1(n_2092),
.B2(n_1995),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2127),
.Y(n_2140)
);

NAND2x1_ASAP7_75t_SL g2141 ( 
.A(n_2122),
.B(n_2096),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2127),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2105),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_2109),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2104),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2115),
.B(n_2095),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2104),
.Y(n_2147)
);

OAI21xp5_ASAP7_75t_SL g2148 ( 
.A1(n_2108),
.A2(n_2097),
.B(n_2089),
.Y(n_2148)
);

AOI222xp33_ASAP7_75t_L g2149 ( 
.A1(n_2120),
.A2(n_2070),
.B1(n_2072),
.B2(n_2077),
.C1(n_2076),
.C2(n_2097),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2105),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2144),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2141),
.Y(n_2152)
);

HB1xp67_ASAP7_75t_L g2153 ( 
.A(n_2144),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2131),
.B(n_2098),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2146),
.B(n_2122),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2129),
.A2(n_2109),
.B1(n_2121),
.B2(n_2126),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2133),
.B(n_2134),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2146),
.B(n_2122),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2136),
.B(n_2115),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2138),
.B(n_2111),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2128),
.B(n_2116),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2135),
.B(n_2123),
.Y(n_2162)
);

OAI21xp5_ASAP7_75t_SL g2163 ( 
.A1(n_2130),
.A2(n_2132),
.B(n_2148),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2143),
.B(n_2116),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2140),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2149),
.B(n_2111),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_2155),
.B(n_2111),
.Y(n_2167)
);

OAI22xp33_ASAP7_75t_SL g2168 ( 
.A1(n_2152),
.A2(n_2150),
.B1(n_2143),
.B2(n_2125),
.Y(n_2168)
);

O2A1O1Ixp33_ASAP7_75t_L g2169 ( 
.A1(n_2163),
.A2(n_2157),
.B(n_2156),
.C(n_2166),
.Y(n_2169)
);

OAI211xp5_ASAP7_75t_L g2170 ( 
.A1(n_2156),
.A2(n_2150),
.B(n_2137),
.C(n_2125),
.Y(n_2170)
);

OAI321xp33_ASAP7_75t_L g2171 ( 
.A1(n_2158),
.A2(n_2101),
.A3(n_2123),
.B1(n_2145),
.B2(n_2142),
.C(n_2147),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2155),
.B(n_2111),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2153),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2155),
.B(n_2101),
.Y(n_2174)
);

OAI221xp5_ASAP7_75t_L g2175 ( 
.A1(n_2154),
.A2(n_2106),
.B1(n_2124),
.B2(n_2139),
.C(n_2089),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2164),
.B(n_2109),
.Y(n_2176)
);

OA21x2_ASAP7_75t_L g2177 ( 
.A1(n_2153),
.A2(n_2124),
.B(n_2106),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2162),
.B(n_2119),
.Y(n_2178)
);

OAI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_2160),
.A2(n_2076),
.B1(n_2021),
.B2(n_2040),
.Y(n_2179)
);

OAI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2169),
.A2(n_2119),
.B1(n_2161),
.B2(n_2159),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2177),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2177),
.Y(n_2182)
);

AOI22x1_ASAP7_75t_L g2183 ( 
.A1(n_2178),
.A2(n_2159),
.B1(n_2165),
.B2(n_2151),
.Y(n_2183)
);

AOI221xp5_ASAP7_75t_L g2184 ( 
.A1(n_2171),
.A2(n_2094),
.B1(n_2084),
.B2(n_2075),
.C(n_2068),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2170),
.A2(n_1983),
.B1(n_1990),
.B2(n_2075),
.Y(n_2185)
);

OAI322xp33_ASAP7_75t_L g2186 ( 
.A1(n_2176),
.A2(n_2094),
.A3(n_2059),
.B1(n_2084),
.B2(n_2075),
.C1(n_2068),
.C2(n_2064),
.Y(n_2186)
);

AOI221xp5_ASAP7_75t_L g2187 ( 
.A1(n_2168),
.A2(n_2094),
.B1(n_2059),
.B2(n_2084),
.C(n_2068),
.Y(n_2187)
);

AOI221xp5_ASAP7_75t_L g2188 ( 
.A1(n_2175),
.A2(n_2064),
.B1(n_2059),
.B2(n_2033),
.C(n_2042),
.Y(n_2188)
);

NOR2x1_ASAP7_75t_L g2189 ( 
.A(n_2181),
.B(n_2173),
.Y(n_2189)
);

INVx1_ASAP7_75t_SL g2190 ( 
.A(n_2183),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2180),
.B(n_2167),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2182),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2186),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2185),
.B(n_2174),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2188),
.B(n_2172),
.Y(n_2195)
);

AOI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_2190),
.A2(n_2179),
.B1(n_2184),
.B2(n_2187),
.C(n_2064),
.Y(n_2196)
);

NOR2x1_ASAP7_75t_L g2197 ( 
.A(n_2189),
.B(n_2021),
.Y(n_2197)
);

INVx2_ASAP7_75t_SL g2198 ( 
.A(n_2194),
.Y(n_2198)
);

INVx2_ASAP7_75t_SL g2199 ( 
.A(n_2191),
.Y(n_2199)
);

OAI21xp5_ASAP7_75t_L g2200 ( 
.A1(n_2193),
.A2(n_2030),
.B(n_2023),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2192),
.Y(n_2201)
);

OAI222xp33_ASAP7_75t_L g2202 ( 
.A1(n_2199),
.A2(n_2198),
.B1(n_2197),
.B2(n_2195),
.C1(n_2201),
.C2(n_2196),
.Y(n_2202)
);

AND3x2_ASAP7_75t_L g2203 ( 
.A(n_2200),
.B(n_1737),
.C(n_1783),
.Y(n_2203)
);

AOI311xp33_ASAP7_75t_L g2204 ( 
.A1(n_2200),
.A2(n_2047),
.A3(n_2042),
.B(n_2040),
.C(n_2038),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2202),
.B(n_2024),
.Y(n_2205)
);

OAI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2205),
.A2(n_2204),
.B1(n_2203),
.B2(n_2030),
.C(n_2036),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2206),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2206),
.Y(n_2208)
);

XNOR2xp5_ASAP7_75t_L g2209 ( 
.A(n_2208),
.B(n_2009),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2207),
.Y(n_2210)
);

INVx1_ASAP7_75t_SL g2211 ( 
.A(n_2209),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2210),
.Y(n_2212)
);

OAI22xp33_ASAP7_75t_L g2213 ( 
.A1(n_2211),
.A2(n_2038),
.B1(n_2036),
.B2(n_2033),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_2213),
.Y(n_2214)
);

OAI21xp5_ASAP7_75t_L g2215 ( 
.A1(n_2214),
.A2(n_2212),
.B(n_2023),
.Y(n_2215)
);

AOI222xp33_ASAP7_75t_L g2216 ( 
.A1(n_2215),
.A2(n_2047),
.B1(n_1981),
.B2(n_2026),
.C1(n_2032),
.C2(n_1991),
.Y(n_2216)
);

AOI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2216),
.A2(n_1981),
.B1(n_1972),
.B2(n_1961),
.C(n_1991),
.Y(n_2217)
);

AOI211xp5_ASAP7_75t_L g2218 ( 
.A1(n_2217),
.A2(n_2027),
.B(n_2024),
.C(n_1990),
.Y(n_2218)
);


endmodule