module fake_jpeg_3475_n_126 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_33),
.Y(n_60)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_45),
.Y(n_61)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_65),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_38),
.B1(n_45),
.B2(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_44),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.C(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_0),
.Y(n_83)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_51),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_50),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_73),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_4),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_51),
.B1(n_41),
.B2(n_39),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_13),
.B1(n_28),
.B2(n_27),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_92),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_80),
.B1(n_81),
.B2(n_79),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_101),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_17),
.B(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_11),
.C(n_23),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_103),
.A3(n_95),
.B1(n_102),
.B2(n_96),
.C(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_117),
.C(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_114),
.C(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_118),
.C(n_113),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_117),
.Y(n_126)
);


endmodule