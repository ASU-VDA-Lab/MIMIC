module fake_jpeg_17111_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_4),
.B(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_25),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_2),
.C(n_3),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_17),
.B(n_7),
.C(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_10),
.C(n_17),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_34),
.C(n_15),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_16),
.B(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_16),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_39),
.B(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_15),
.B1(n_35),
.B2(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_29),
.B1(n_31),
.B2(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_46),
.B1(n_38),
.B2(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_47),
.A2(n_15),
.B1(n_42),
.B2(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_53),
.B1(n_51),
.B2(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_57),
.Y(n_61)
);


endmodule