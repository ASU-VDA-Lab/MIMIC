module real_jpeg_9547_n_12 (n_5, n_4, n_8, n_0, n_327, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_327;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_4),
.B(n_21),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_4),
.A2(n_11),
.B(n_25),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_9),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_38),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_5),
.A2(n_21),
.B1(n_32),
.B2(n_38),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_5),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_21),
.B1(n_32),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_7),
.A2(n_41),
.B(n_54),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_7),
.B(n_41),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_7),
.A2(n_11),
.B(n_41),
.C(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_9),
.B1(n_37),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_8),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_104),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_8),
.A2(n_21),
.B1(n_32),
.B2(n_104),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_10),
.B1(n_37),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_47),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_21),
.B1(n_32),
.B2(n_47),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_11),
.A2(n_21),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_11),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_37),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_11),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_70),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_53),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_80),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_78),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_72),
.Y(n_14)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_15),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_63),
.C(n_65),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_16),
.A2(n_17),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_50),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_18),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_18),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_18),
.A2(n_106),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_18),
.A2(n_50),
.B1(n_51),
.B2(n_106),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_29),
.B(n_30),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_19),
.A2(n_97),
.B(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_20),
.B(n_170),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_20),
.B(n_98),
.Y(n_206)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_21),
.A2(n_33),
.B(n_55),
.Y(n_201)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_24),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_24),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_24),
.B(n_31),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_91),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_28),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_29),
.B(n_33),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_29),
.A2(n_206),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_33),
.B(n_91),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_34),
.A2(n_35),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B(n_44),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_36),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_39),
.B(n_40),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_39),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_39),
.A2(n_48),
.B(n_76),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_39)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_41),
.B(n_43),
.Y(n_131)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_42),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_45),
.B(n_102),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_48),
.B(n_76),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_49),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_59),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_54),
.B(n_62),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_54),
.A2(n_57),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_56),
.B(n_58),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_58),
.A2(n_144),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_59),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_63),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_63),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_63),
.A2(n_65),
.B1(n_249),
.B2(n_322),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_69),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_74),
.B(n_115),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_77),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_318),
.B(n_324),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_294),
.A3(n_313),
.B1(n_316),
.B2(n_317),
.C(n_327),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_272),
.B(n_293),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_253),
.B(n_271),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_152),
.B(n_235),
.C(n_252),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_135),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_86),
.B(n_135),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_111),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_100),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_88),
.B(n_100),
.C(n_111),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_89),
.B(n_96),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_94),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_90),
.A2(n_91),
.B(n_150),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_93),
.B(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_92),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_92),
.B(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_94),
.B(n_175),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_97),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_107),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_101),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_105),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_106),
.B(n_298),
.C(n_303),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_109),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_122),
.B1(n_123),
.B2(n_134),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_121),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_113),
.B(n_121),
.C(n_122),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_126),
.B(n_192),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_136),
.A2(n_137),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_231)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_143),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_144),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_234),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_228),
.B(n_233),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_213),
.B(n_227),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_194),
.B(n_212),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_182),
.B(n_193),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_171),
.B(n_181),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_163),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_165),
.B(n_167),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_180),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B1(n_204),
.B2(n_211),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_197),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_198),
.A2(n_199),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_198),
.A2(n_199),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_198),
.A2(n_286),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_199),
.B(n_268),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_223),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_222),
.C(n_226),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_222),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_236),
.B(n_237),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_250),
.B2(n_251),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_244),
.C(n_251),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_242),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_248),
.C(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_250),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_255),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_267),
.C(n_270),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_261),
.C(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_274),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_291),
.B2(n_292),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_282),
.B1(n_289),
.B2(n_290),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_290),
.C(n_292),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B(n_281),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_279),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_296),
.C(n_305),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_281),
.B(n_296),
.CI(n_305),
.CON(n_315),
.SN(n_315)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_287),
.B2(n_288),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_306),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_298),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_308),
.C(n_312),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_314),
.B(n_315),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_315),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_321),
.Y(n_323)
);


endmodule