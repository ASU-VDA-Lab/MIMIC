module fake_jpeg_27676_n_58 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_27),
.B1(n_25),
.B2(n_5),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_8),
.C(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_2),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_43),
.B(n_35),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_27),
.B1(n_25),
.B2(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_48),
.C(n_49),
.Y(n_53)
);

NOR4xp25_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_4),
.C(n_6),
.D(n_7),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_39),
.B(n_41),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_38),
.C(n_50),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_52),
.C(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_43),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_44),
.B(n_51),
.C(n_11),
.Y(n_57)
);

AOI321xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_4),
.A3(n_7),
.B1(n_18),
.B2(n_51),
.C(n_41),
.Y(n_58)
);


endmodule