module real_aes_6832_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_516;
wire n_177;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_0), .A2(n_127), .B1(n_133), .B2(n_721), .C1(n_722), .C2(n_725), .Y(n_126) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g462 ( .A(n_2), .Y(n_462) );
INVx1_ASAP7_75t_L g266 ( .A(n_3), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_4), .A2(n_37), .B1(n_216), .B2(n_501), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g227 ( .A1(n_5), .A2(n_149), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_6), .B(n_171), .Y(n_487) );
AND2x6_ASAP7_75t_L g154 ( .A(n_7), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_8), .A2(n_148), .B(n_156), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_9), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_9), .B(n_38), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_10), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g233 ( .A(n_11), .Y(n_233) );
INVx1_ASAP7_75t_L g146 ( .A(n_12), .Y(n_146) );
INVx1_ASAP7_75t_L g456 ( .A(n_13), .Y(n_456) );
INVx1_ASAP7_75t_L g166 ( .A(n_14), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_15), .B(n_240), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_16), .B(n_172), .Y(n_489) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_17), .A2(n_171), .A3(n_187), .B1(n_475), .B2(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_18), .B(n_216), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_19), .B(n_183), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_20), .B(n_172), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_48), .B1(n_216), .B2(n_501), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_22), .B(n_149), .Y(n_176) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_23), .A2(n_77), .B1(n_216), .B2(n_240), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_24), .B(n_216), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_25), .B(n_226), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_26), .A2(n_163), .B(n_165), .C(n_167), .Y(n_162) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_27), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_28), .B(n_142), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_29), .B(n_198), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_30), .A2(n_101), .B1(n_129), .B2(n_130), .Y(n_128) );
INVx1_ASAP7_75t_L g130 ( .A(n_30), .Y(n_130) );
INVx1_ASAP7_75t_L g245 ( .A(n_31), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_32), .B(n_142), .Y(n_513) );
INVx2_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_34), .B(n_216), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_35), .B(n_142), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_36), .A2(n_154), .B(n_159), .C(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g113 ( .A(n_38), .Y(n_113) );
INVx1_ASAP7_75t_L g243 ( .A(n_39), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_40), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_41), .B(n_216), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_42), .A2(n_87), .B1(n_168), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_43), .B(n_216), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_44), .B(n_216), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_45), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_46), .B(n_461), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_47), .B(n_149), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_49), .A2(n_59), .B1(n_216), .B2(n_240), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_50), .A2(n_734), .B1(n_737), .B2(n_738), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_50), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_51), .A2(n_159), .B1(n_240), .B2(n_242), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_52), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_53), .B(n_216), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_54), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_55), .B(n_216), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_56), .A2(n_231), .B(n_232), .C(n_234), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_57), .Y(n_202) );
INVx1_ASAP7_75t_L g229 ( .A(n_58), .Y(n_229) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_61), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_61), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_62), .B(n_216), .Y(n_463) );
INVx1_ASAP7_75t_L g145 ( .A(n_63), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_64), .A2(n_75), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_64), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
AO32x2_ASAP7_75t_L g498 ( .A1(n_66), .A2(n_171), .A3(n_208), .B1(n_475), .B2(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
INVx1_ASAP7_75t_L g508 ( .A(n_68), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_SL g253 ( .A1(n_69), .A2(n_183), .B(n_234), .C(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_L g255 ( .A(n_70), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_71), .B(n_240), .Y(n_509) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_73), .Y(n_248) );
INVx1_ASAP7_75t_L g193 ( .A(n_74), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_75), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_76), .A2(n_104), .B1(n_114), .B2(n_741), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_78), .A2(n_154), .B(n_159), .C(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_79), .B(n_501), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_80), .B(n_240), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_81), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_83), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_84), .B(n_240), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_85), .A2(n_154), .B(n_159), .C(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g108 ( .A(n_86), .Y(n_108) );
OR2x2_ASAP7_75t_L g121 ( .A(n_86), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g134 ( .A(n_86), .B(n_123), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_88), .A2(n_102), .B1(n_240), .B2(n_241), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_89), .B(n_142), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_90), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_91), .A2(n_154), .B(n_159), .C(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_92), .Y(n_219) );
INVx1_ASAP7_75t_L g252 ( .A(n_93), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g157 ( .A(n_94), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_95), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_96), .B(n_180), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_97), .B(n_240), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_98), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_100), .A2(n_149), .B(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_101), .Y(n_129) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g742 ( .A(n_105), .Y(n_742) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g123 ( .A(n_107), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g445 ( .A(n_108), .B(n_123), .Y(n_445) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_108), .B(n_122), .Y(n_727) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_126), .B1(n_728), .B2(n_730), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_119), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g729 ( .A(n_118), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_119), .A2(n_731), .B(n_739), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g119 ( .A(n_120), .B(n_125), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g740 ( .A(n_121), .Y(n_740) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g721 ( .A(n_127), .Y(n_721) );
INVx1_ASAP7_75t_L g131 ( .A(n_128), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B1(n_443), .B2(n_446), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_134), .A2(n_445), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_135), .Y(n_723) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_135), .A2(n_723), .B1(n_732), .B2(n_733), .Y(n_731) );
OR4x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_339), .C(n_398), .D(n_425), .Y(n_135) );
NAND3xp33_ASAP7_75t_SL g136 ( .A(n_137), .B(n_281), .C(n_306), .Y(n_136) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_204), .B(n_224), .C(n_257), .Y(n_137) );
AOI211xp5_ASAP7_75t_SL g429 ( .A1(n_138), .A2(n_430), .B(n_432), .C(n_435), .Y(n_429) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_173), .Y(n_138) );
INVx1_ASAP7_75t_L g304 ( .A(n_139), .Y(n_304) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g279 ( .A(n_140), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g311 ( .A(n_140), .Y(n_311) );
AND2x2_ASAP7_75t_L g366 ( .A(n_140), .B(n_335), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_140), .B(n_222), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_140), .B(n_223), .Y(n_424) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g285 ( .A(n_141), .Y(n_285) );
AND2x2_ASAP7_75t_L g328 ( .A(n_141), .B(n_191), .Y(n_328) );
AND2x2_ASAP7_75t_L g346 ( .A(n_141), .B(n_223), .Y(n_346) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_170), .Y(n_141) );
INVx1_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
INVx2_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_142), .A2(n_506), .B(n_513), .Y(n_505) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_142), .A2(n_515), .B(n_523), .Y(n_514) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_L g172 ( .A(n_143), .B(n_144), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_154), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_150), .B(n_154), .Y(n_194) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
INVx1_ASAP7_75t_L g461 ( .A(n_151), .Y(n_461) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g241 ( .A(n_152), .Y(n_241) );
INVx1_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
INVx3_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
INVx1_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
INVx4_ASAP7_75t_SL g169 ( .A(n_154), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_154), .A2(n_455), .B(n_459), .Y(n_454) );
BUFx3_ASAP7_75t_L g475 ( .A(n_154), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_154), .A2(n_481), .B(n_484), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_154), .A2(n_507), .B(n_510), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_154), .A2(n_516), .B(n_520), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_162), .C(n_169), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_158), .A2(n_169), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_158), .A2(n_169), .B(n_252), .C(n_253), .Y(n_251) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx3_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVx1_ASAP7_75t_L g501 ( .A(n_160), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_163), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g458 ( .A(n_163), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_163), .A2(n_511), .B(n_512), .Y(n_510) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g242 ( .A1(n_164), .A2(n_243), .B1(n_244), .B2(n_245), .Y(n_242) );
INVx2_ASAP7_75t_L g244 ( .A(n_164), .Y(n_244) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_169), .A2(n_194), .B1(n_239), .B2(n_246), .Y(n_238) );
INVx4_ASAP7_75t_L g190 ( .A(n_171), .Y(n_190) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_171), .A2(n_250), .B(n_256), .Y(n_249) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_171), .A2(n_480), .B(n_487), .Y(n_479) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g187 ( .A(n_172), .Y(n_187) );
INVx4_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_173), .A2(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g414 ( .A(n_173), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_191), .Y(n_173) );
INVx1_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
AND2x2_ASAP7_75t_L g283 ( .A(n_174), .B(n_223), .Y(n_283) );
OR2x2_ASAP7_75t_L g312 ( .A(n_174), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g326 ( .A(n_174), .Y(n_326) );
INVx3_ASAP7_75t_L g335 ( .A(n_174), .Y(n_335) );
AND2x2_ASAP7_75t_L g345 ( .A(n_174), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g378 ( .A(n_174), .B(n_284), .Y(n_378) );
AND2x2_ASAP7_75t_L g402 ( .A(n_174), .B(n_358), .Y(n_402) );
OR2x6_ASAP7_75t_L g174 ( .A(n_175), .B(n_188), .Y(n_174) );
AOI21xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_186), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_184), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_180), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
INVx2_ASAP7_75t_L g464 ( .A(n_180), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_180), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_180), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_SL g507 ( .A1(n_180), .A2(n_234), .B(n_508), .C(n_509), .Y(n_507) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_181), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_181), .B(n_255), .Y(n_254) );
OAI22xp5_ASAP7_75t_SL g499 ( .A1(n_181), .A2(n_198), .B1(n_500), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_183), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_184), .A2(n_197), .B(n_199), .Y(n_196) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g200 ( .A(n_186), .Y(n_200) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_186), .A2(n_454), .B(n_465), .Y(n_453) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_186), .A2(n_468), .B(n_476), .Y(n_467) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_187), .A2(n_238), .B(n_247), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_187), .B(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_187), .A2(n_262), .B(n_269), .Y(n_261) );
NOR2xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx3_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_190), .B(n_475), .C(n_491), .Y(n_490) );
AO21x1_ASAP7_75t_L g569 ( .A1(n_190), .A2(n_491), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g223 ( .A(n_191), .Y(n_223) );
AND2x2_ASAP7_75t_L g438 ( .A(n_191), .B(n_280), .Y(n_438) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_200), .B(n_201), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_194), .A2(n_263), .B(n_264), .Y(n_262) );
INVx4_ASAP7_75t_L g214 ( .A(n_198), .Y(n_214) );
INVx2_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_198), .A2(n_464), .B1(n_492), .B2(n_493), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_198), .A2(n_464), .B1(n_537), .B2(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_203), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_203), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_220), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_206), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g358 ( .A(n_206), .B(n_346), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_206), .B(n_335), .Y(n_420) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
AND2x2_ASAP7_75t_L g284 ( .A(n_207), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g325 ( .A(n_207), .B(n_326), .Y(n_325) );
AO21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_218), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_217), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_215), .Y(n_211) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g234 ( .A(n_216), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_220), .B(n_321), .Y(n_343) );
INVx1_ASAP7_75t_L g382 ( .A(n_220), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_220), .B(n_309), .Y(n_426) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g289 ( .A(n_221), .B(n_284), .Y(n_289) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_223), .B(n_280), .Y(n_313) );
INVx1_ASAP7_75t_L g392 ( .A(n_223), .Y(n_392) );
AOI322xp5_ASAP7_75t_L g416 ( .A1(n_224), .A2(n_331), .A3(n_391), .B1(n_417), .B2(n_419), .C1(n_421), .C2(n_423), .Y(n_416) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_225), .B(n_236), .Y(n_224) );
AND2x2_ASAP7_75t_L g271 ( .A(n_225), .B(n_249), .Y(n_271) );
INVx1_ASAP7_75t_SL g274 ( .A(n_225), .Y(n_274) );
AND2x2_ASAP7_75t_L g276 ( .A(n_225), .B(n_237), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_225), .B(n_293), .Y(n_299) );
INVx2_ASAP7_75t_L g318 ( .A(n_225), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_225), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g369 ( .A(n_225), .B(n_293), .Y(n_369) );
BUFx2_ASAP7_75t_L g386 ( .A(n_225), .Y(n_386) );
AND2x2_ASAP7_75t_L g400 ( .A(n_225), .B(n_260), .Y(n_400) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g472 ( .A1(n_231), .A2(n_460), .B(n_473), .C(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_231), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_236), .B(n_288), .Y(n_315) );
AND2x2_ASAP7_75t_L g442 ( .A(n_236), .B(n_318), .Y(n_442) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_249), .Y(n_236) );
OR2x2_ASAP7_75t_L g287 ( .A(n_237), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g293 ( .A(n_237), .Y(n_293) );
AND2x2_ASAP7_75t_L g338 ( .A(n_237), .B(n_261), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_237), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_237), .Y(n_422) );
INVx2_ASAP7_75t_L g268 ( .A(n_240), .Y(n_268) );
INVx3_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g273 ( .A(n_249), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g295 ( .A(n_249), .Y(n_295) );
BUFx2_ASAP7_75t_L g301 ( .A(n_249), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_249), .B(n_293), .Y(n_320) );
INVx3_ASAP7_75t_L g332 ( .A(n_249), .Y(n_332) );
OR2x2_ASAP7_75t_L g342 ( .A(n_249), .B(n_293), .Y(n_342) );
AOI31xp33_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_272), .A3(n_275), .B(n_277), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_271), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_259), .B(n_294), .Y(n_305) );
OR2x2_ASAP7_75t_L g329 ( .A(n_259), .B(n_299), .Y(n_329) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_260), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g350 ( .A(n_260), .B(n_342), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_260), .B(n_332), .Y(n_360) );
AND2x2_ASAP7_75t_L g367 ( .A(n_260), .B(n_368), .Y(n_367) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_260), .B(n_331), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_260), .B(n_386), .Y(n_396) );
AND2x2_ASAP7_75t_L g408 ( .A(n_260), .B(n_293), .Y(n_408) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g288 ( .A(n_261), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_268), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g354 ( .A(n_271), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_271), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_273), .B(n_349), .Y(n_383) );
AND2x4_ASAP7_75t_L g294 ( .A(n_274), .B(n_295), .Y(n_294) );
CKINVDCx16_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g373 ( .A(n_279), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_279), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_311), .Y(n_321) );
AND2x2_ASAP7_75t_L g415 ( .A(n_280), .B(n_285), .Y(n_415) );
INVx1_ASAP7_75t_L g440 ( .A(n_280), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_286), .B1(n_289), .B2(n_290), .C(n_296), .Y(n_281) );
CKINVDCx14_ASAP7_75t_R g302 ( .A(n_282), .Y(n_302) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_283), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_286), .B(n_337), .Y(n_356) );
INVx3_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g405 ( .A(n_287), .B(n_301), .Y(n_405) );
AND2x2_ASAP7_75t_L g319 ( .A(n_288), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_288), .B(n_332), .Y(n_377) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_288), .B(n_389), .C(n_420), .Y(n_419) );
AOI211xp5_ASAP7_75t_SL g352 ( .A1(n_289), .A2(n_353), .B(n_355), .C(n_363), .Y(n_352) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_342), .B1(n_343), .B2(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_292), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_292), .B(n_376), .Y(n_375) );
BUFx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g434 ( .A(n_294), .B(n_408), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_302), .B1(n_303), .B2(n_305), .Y(n_296) );
NOR2xp33_ASAP7_75t_SL g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_300), .B(n_349), .Y(n_380) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_303), .A2(n_395), .B1(n_426), .B2(n_433), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_314), .B1(n_316), .B2(n_321), .C(n_322), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_312), .A2(n_323), .B1(n_329), .B2(n_330), .C(n_333), .Y(n_322) );
INVx1_ASAP7_75t_L g365 ( .A(n_313), .Y(n_365) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_SL g337 ( .A(n_318), .Y(n_337) );
OR2x2_ASAP7_75t_L g410 ( .A(n_318), .B(n_342), .Y(n_410) );
AND2x2_ASAP7_75t_L g412 ( .A(n_318), .B(n_320), .Y(n_412) );
INVx1_ASAP7_75t_L g351 ( .A(n_321), .Y(n_351) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_324), .A2(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g388 ( .A(n_324), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g362 ( .A(n_325), .B(n_346), .Y(n_362) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp33_ASAP7_75t_SL g379 ( .A(n_330), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_331), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_332), .B(n_368), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_335), .A2(n_348), .B(n_350), .C(n_351), .Y(n_347) );
NAND2x1_ASAP7_75t_SL g372 ( .A(n_335), .B(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_336), .A2(n_385), .B1(n_387), .B2(n_390), .Y(n_384) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_338), .B(n_428), .Y(n_427) );
NAND5xp2_ASAP7_75t_L g339 ( .A(n_340), .B(n_352), .C(n_370), .D(n_384), .E(n_393), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_347), .Y(n_340) );
INVx1_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_345), .A2(n_364), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_346), .B(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_349), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_349), .B(n_415), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_361), .Y(n_355) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g437 ( .A(n_366), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B1(n_378), .B2(n_379), .C(n_381), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g421 ( .A(n_376), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g428 ( .A(n_386), .Y(n_428) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_396), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_401), .B(n_403), .C(n_416), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_401), .A2(n_426), .B(n_427), .C(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_405), .B(n_407), .Y(n_406) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g724 ( .A(n_446), .Y(n_724) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR5x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_612), .C(n_670), .D(n_706), .E(n_713), .Y(n_448) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_558), .C(n_582), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_494), .B1(n_524), .B2(n_529), .C(n_539), .Y(n_450) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_451), .A2(n_693), .B(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_477), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_452), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_466), .Y(n_452) );
INVx2_ASAP7_75t_L g528 ( .A(n_453), .Y(n_528) );
AND2x2_ASAP7_75t_L g541 ( .A(n_453), .B(n_479), .Y(n_541) );
AND2x2_ASAP7_75t_L g595 ( .A(n_453), .B(n_478), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_453), .B(n_467), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B(n_463), .C(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_464), .A2(n_485), .B(n_486), .Y(n_484) );
AND2x2_ASAP7_75t_L g628 ( .A(n_466), .B(n_569), .Y(n_628) );
AND2x2_ASAP7_75t_L g661 ( .A(n_466), .B(n_479), .Y(n_661) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g568 ( .A(n_467), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g581 ( .A(n_467), .B(n_479), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_467), .B(n_569), .Y(n_588) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_467), .Y(n_597) );
AND2x2_ASAP7_75t_L g604 ( .A(n_467), .B(n_478), .Y(n_604) );
INVx1_ASAP7_75t_L g635 ( .A(n_467), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g611 ( .A(n_477), .Y(n_611) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
INVx2_ASAP7_75t_L g567 ( .A(n_478), .Y(n_567) );
AND2x2_ASAP7_75t_L g589 ( .A(n_478), .B(n_528), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_478), .B(n_635), .Y(n_640) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_479), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g712 ( .A(n_479), .B(n_676), .Y(n_712) );
INVx2_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
INVx3_ASAP7_75t_L g627 ( .A(n_488), .Y(n_627) );
OR2x2_ASAP7_75t_L g657 ( .A(n_488), .B(n_658), .Y(n_657) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_488), .B(n_567), .Y(n_683) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g570 ( .A(n_489), .Y(n_570) );
AOI33xp33_ASAP7_75t_L g703 ( .A1(n_494), .A2(n_541), .A3(n_555), .B1(n_627), .B2(n_704), .B3(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .Y(n_495) );
OR2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_496), .B(n_553), .Y(n_615) );
OR2x2_ASAP7_75t_L g668 ( .A(n_496), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g594 ( .A(n_497), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g619 ( .A(n_497), .B(n_503), .Y(n_619) );
AND2x2_ASAP7_75t_L g686 ( .A(n_497), .B(n_531), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_497), .A2(n_586), .B(n_712), .Y(n_711) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g533 ( .A(n_498), .Y(n_533) );
INVx1_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
AND2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_535), .Y(n_565) );
AND2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_534), .Y(n_614) );
INVx2_ASAP7_75t_SL g656 ( .A(n_503), .Y(n_656) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
INVx2_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
INVx1_ASAP7_75t_L g707 ( .A(n_504), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_504), .B(n_601), .Y(n_720) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g547 ( .A(n_505), .Y(n_547) );
OR2x2_ASAP7_75t_L g553 ( .A(n_505), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_514), .Y(n_531) );
AND2x2_ASAP7_75t_L g548 ( .A(n_514), .B(n_534), .Y(n_548) );
INVx1_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_514), .B(n_535), .Y(n_586) );
INVx2_ASAP7_75t_L g602 ( .A(n_514), .Y(n_602) );
AND2x2_ASAP7_75t_L g695 ( .A(n_514), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_514), .B(n_576), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g550 ( .A(n_526), .Y(n_550) );
INVx1_ASAP7_75t_L g579 ( .A(n_526), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_526), .B(n_610), .Y(n_676) );
INVx1_ASAP7_75t_SL g636 ( .A(n_527), .Y(n_636) );
INVx2_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
AND2x2_ASAP7_75t_L g626 ( .A(n_528), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g642 ( .A(n_528), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g704 ( .A(n_530), .Y(n_704) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g559 ( .A(n_532), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g662 ( .A(n_532), .B(n_652), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_532), .A2(n_673), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_L g575 ( .A(n_533), .B(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g600 ( .A(n_533), .Y(n_600) );
INVx1_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
OR2x2_ASAP7_75t_L g688 ( .A(n_534), .B(n_547), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_534), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .B1(n_549), .B2(n_551), .Y(n_539) );
OR2x2_ASAP7_75t_L g618 ( .A(n_540), .B(n_568), .Y(n_618) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_541), .A2(n_660), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g606 ( .A(n_545), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_547), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_547), .Y(n_631) );
AND2x2_ASAP7_75t_L g679 ( .A(n_547), .B(n_548), .Y(n_679) );
INVx1_ASAP7_75t_L g697 ( .A(n_547), .Y(n_697) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g663 ( .A(n_550), .B(n_589), .Y(n_663) );
AND2x2_ASAP7_75t_L g705 ( .A(n_550), .B(n_581), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_552), .B(n_600), .Y(n_687) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_553), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g580 ( .A(n_557), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g648 ( .A(n_557), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_566), .C(n_571), .Y(n_558) );
INVxp67_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_560), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_560), .B(n_607), .Y(n_702) );
BUFx3_ASAP7_75t_L g666 ( .A(n_561), .Y(n_666) );
INVx1_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g592 ( .A(n_564), .B(n_586), .Y(n_592) );
INVx1_ASAP7_75t_SL g632 ( .A(n_565), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
AND2x2_ASAP7_75t_L g645 ( .A(n_567), .B(n_628), .Y(n_645) );
INVx1_ASAP7_75t_SL g616 ( .A(n_568), .Y(n_616) );
INVx1_ASAP7_75t_L g643 ( .A(n_569), .Y(n_643) );
AOI31xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .A3(n_574), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g664 ( .A(n_575), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g638 ( .A(n_576), .Y(n_638) );
BUFx2_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
AND2x2_ASAP7_75t_L g680 ( .A(n_576), .B(n_601), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g653 ( .A(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_581), .B(n_648), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_581), .B(n_627), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B(n_590), .C(n_605), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_587), .A2(n_614), .B1(n_615), .B2(n_616), .C(n_617), .Y(n_613) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g621 ( .A(n_588), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
OAI32xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_596), .B1(n_598), .B2(n_603), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_592), .A2(n_645), .B(n_646), .C(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_600), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g669 ( .A(n_601), .Y(n_669) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_607), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g655 ( .A(n_607), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g672 ( .A(n_609), .Y(n_672) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_625), .C(n_644), .D(n_659), .Y(n_612) );
AND2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g673 ( .A(n_614), .B(n_666), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_616), .B(n_648), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_620), .B2(n_623), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_618), .A2(n_669), .B1(n_700), .B2(n_702), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_618), .A2(n_707), .B(n_708), .C(n_711), .Y(n_706) );
INVx2_ASAP7_75t_L g677 ( .A(n_619), .Y(n_677) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_621), .A2(n_655), .B1(n_672), .B2(n_673), .C1(n_674), .C2(n_677), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_629), .C(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g691 ( .A(n_626), .Y(n_691) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_630), .A2(n_634), .B1(n_637), .B2(n_639), .Y(n_633) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g660 ( .A(n_642), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g718 ( .A(n_645), .Y(n_718) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_654), .B2(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_652), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g709 ( .A(n_657), .Y(n_709) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g717 ( .A(n_663), .Y(n_717) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND5xp2_ASAP7_75t_L g670 ( .A(n_671), .B(n_678), .C(n_692), .D(n_698), .E(n_703), .Y(n_670) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_681), .C(n_684), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI31xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .A3(n_688), .B(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g710 ( .A(n_686), .Y(n_710) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI222xp33_ASAP7_75t_L g713 ( .A1(n_700), .A2(n_702), .B1(n_714), .B2(n_717), .C1(n_718), .C2(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_734), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
endmodule