module fake_aes_9639_n_14 (n_1, n_2, n_4, n_3, n_5, n_0, n_14);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_7;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_2), .B(n_0), .Y(n_7) );
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_5), .B(n_1), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
BUFx4f_ASAP7_75t_SL g10 ( .A(n_7), .Y(n_10) );
AND2x4_ASAP7_75t_L g11 ( .A(n_9), .B(n_8), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_11), .B(n_9), .Y(n_12) );
OA22x2_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_11), .B1(n_10), .B2(n_2), .Y(n_13) );
AOI21xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_4), .B(n_1), .Y(n_14) );
endmodule