module fake_jpeg_25527_n_147 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_82),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_62),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_65),
.B(n_49),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_54),
.B(n_67),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_60),
.B(n_55),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_56),
.B(n_64),
.C(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_49),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_7),
.C(n_8),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_48),
.B1(n_50),
.B2(n_65),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_96),
.B1(n_4),
.B2(n_5),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_97),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_77),
.B1(n_73),
.B2(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_89),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_7),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_63),
.B1(n_58),
.B2(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_68),
.B1(n_51),
.B2(n_64),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_57),
.B1(n_20),
.B2(n_45),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_44),
.B1(n_21),
.B2(n_22),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_19),
.B1(n_42),
.B2(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_8),
.Y(n_121)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_18),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_9),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_106),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_105),
.C(n_24),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_132),
.C(n_133),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_113),
.B(n_93),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_114),
.B1(n_93),
.B2(n_9),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_115),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_139),
.C(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_134),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_124),
.C(n_11),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_34),
.B(n_15),
.C(n_17),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_30),
.A3(n_36),
.B1(n_43),
.B2(n_118),
.C(n_10),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_145),
.B(n_10),
.CI(n_132),
.CON(n_146),
.SN(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_146),
.Y(n_147)
);


endmodule