module fake_aes_12329_n_755 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_755);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_755;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_87), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_22), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_93), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_0), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_62), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_51), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_7), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_57), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_81), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_18), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_54), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_39), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_45), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_77), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_42), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_98), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_73), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_1), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_21), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_22), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_16), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_63), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_10), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_9), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_36), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_33), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_50), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_14), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_21), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_23), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_78), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_109), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_134), .B(n_0), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_134), .B(n_2), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_131), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_114), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_127), .B(n_3), .Y(n_148) );
OR2x6_ASAP7_75t_L g149 ( .A(n_136), .B(n_5), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_109), .B(n_5), .Y(n_150) );
OAI22xp5_ASAP7_75t_L g151 ( .A1(n_105), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_115), .B(n_6), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_103), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_115), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
OAI21x1_ASAP7_75t_L g156 ( .A1(n_141), .A2(n_58), .B(n_100), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_104), .B(n_106), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_110), .Y(n_159) );
NAND2xp33_ASAP7_75t_L g160 ( .A(n_102), .B(n_56), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_161), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_149), .B(n_105), .Y(n_164) );
INVxp67_ASAP7_75t_SL g165 ( .A(n_157), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_157), .B(n_112), .Y(n_166) );
OR2x2_ASAP7_75t_L g167 ( .A(n_148), .B(n_118), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_143), .B(n_128), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_113), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_161), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_143), .B(n_117), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_149), .A2(n_107), .B1(n_126), .B2(n_139), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_154), .Y(n_174) );
AOI22xp33_ASAP7_75t_SL g175 ( .A1(n_144), .A2(n_138), .B1(n_126), .B2(n_139), .Y(n_175) );
BUFx8_ASAP7_75t_SL g176 ( .A(n_149), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_149), .B(n_107), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_144), .B(n_119), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_150), .B(n_125), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_154), .B(n_135), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx2_ASAP7_75t_SL g183 ( .A(n_158), .Y(n_183) );
INVxp33_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_154), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_161), .Y(n_186) );
INVx3_ASAP7_75t_R g187 ( .A(n_149), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_146), .B(n_155), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_156), .A2(n_123), .B(n_140), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_147), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_164), .A2(n_158), .B1(n_152), .B2(n_132), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_164), .A2(n_158), .B1(n_129), .B2(n_133), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_164), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_190), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_165), .B(n_158), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_166), .B(n_158), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_190), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_173), .B(n_137), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_184), .A2(n_173), .B1(n_164), .B2(n_177), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_164), .B(n_129), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_171), .A2(n_156), .B(n_121), .C(n_108), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_167), .B(n_158), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_178), .B(n_122), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_190), .A2(n_160), .B(n_106), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_177), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_167), .B(n_110), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_169), .B(n_158), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_177), .A2(n_145), .B1(n_153), .B2(n_158), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_183), .B(n_110), .Y(n_213) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_124), .B(n_121), .C(n_111), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_177), .B(n_132), .Y(n_215) );
BUFx8_ASAP7_75t_L g216 ( .A(n_176), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_177), .B(n_133), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_172), .B(n_108), .Y(n_219) );
AND2x6_ASAP7_75t_SL g220 ( .A(n_168), .B(n_111), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_179), .B(n_116), .Y(n_221) );
INVxp67_ASAP7_75t_SL g222 ( .A(n_174), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_174), .B(n_116), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_175), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_185), .B(n_120), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_189), .B(n_120), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_187), .B(n_123), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_189), .B(n_130), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_191), .A2(n_151), .B1(n_155), .B2(n_146), .Y(n_231) );
AND2x6_ASAP7_75t_SL g232 ( .A(n_188), .B(n_130), .Y(n_232) );
BUFx12f_ASAP7_75t_L g233 ( .A(n_216), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_209), .B(n_187), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_199), .A2(n_182), .B(n_180), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_209), .B(n_153), .Y(n_236) );
AND3x2_ASAP7_75t_L g237 ( .A(n_216), .B(n_136), .C(n_140), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_146), .Y(n_238) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_141), .B1(n_146), .B2(n_155), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_204), .B(n_155), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_226), .Y(n_241) );
BUFx2_ASAP7_75t_SL g242 ( .A(n_196), .Y(n_242) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_196), .B(n_147), .Y(n_243) );
NAND3xp33_ASAP7_75t_SL g244 ( .A(n_212), .B(n_182), .C(n_180), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_207), .B(n_11), .Y(n_245) );
INVxp33_ASAP7_75t_SL g246 ( .A(n_203), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_214), .A2(n_159), .B(n_147), .C(n_163), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_202), .B(n_11), .Y(n_248) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_197), .A2(n_186), .B(n_170), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g250 ( .A(n_224), .B(n_159), .C(n_170), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_226), .Y(n_251) );
INVx11_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_199), .A2(n_186), .B(n_170), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_214), .A2(n_159), .B(n_163), .C(n_186), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_206), .A2(n_163), .B(n_155), .Y(n_256) );
NOR2x1p5_ASAP7_75t_L g257 ( .A(n_196), .B(n_155), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_215), .B(n_159), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_196), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_206), .A2(n_161), .B(n_59), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_222), .B(n_12), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
CKINVDCx14_ASAP7_75t_R g264 ( .A(n_216), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_194), .B(n_161), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_217), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_211), .A2(n_161), .B(n_60), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
NAND3xp33_ASAP7_75t_SL g269 ( .A(n_250), .B(n_212), .C(n_231), .Y(n_269) );
AO31x2_ASAP7_75t_L g270 ( .A1(n_267), .A2(n_205), .A3(n_201), .B(n_197), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_263), .B(n_236), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g272 ( .A(n_233), .B(n_245), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_249), .A2(n_197), .B(n_201), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_211), .B(n_201), .Y(n_274) );
AND2x2_ASAP7_75t_SL g275 ( .A(n_246), .B(n_217), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_262), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_249), .A2(n_208), .B(n_200), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_248), .A2(n_210), .B(n_219), .C(n_223), .Y(n_279) );
AND2x6_ASAP7_75t_L g280 ( .A(n_261), .B(n_193), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_261), .Y(n_281) );
OAI22x1_ASAP7_75t_L g282 ( .A1(n_257), .A2(n_220), .B1(n_232), .B2(n_228), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_235), .A2(n_208), .B(n_198), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_266), .B(n_193), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_247), .A2(n_195), .B(n_200), .C(n_225), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_254), .A2(n_198), .B(n_195), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_244), .A2(n_230), .B(n_221), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_258), .Y(n_288) );
AO32x2_ASAP7_75t_L g289 ( .A1(n_239), .A2(n_232), .A3(n_220), .B1(n_225), .B2(n_223), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_246), .B(n_230), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_238), .A2(n_229), .B(n_227), .C(n_192), .Y(n_291) );
AO31x2_ASAP7_75t_L g292 ( .A1(n_285), .A2(n_260), .A3(n_240), .B(n_229), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_280), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_275), .B(n_251), .Y(n_294) );
NAND2x1p5_ASAP7_75t_L g295 ( .A(n_281), .B(n_251), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_277), .A2(n_227), .B(n_241), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_273), .A2(n_255), .B(n_257), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_280), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_283), .A2(n_274), .B(n_286), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_280), .B(n_259), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_286), .A2(n_243), .B(n_265), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_271), .A2(n_239), .B1(n_264), .B2(n_241), .C(n_242), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_287), .A2(n_253), .B(n_234), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_268), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_288), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
OR2x6_ASAP7_75t_L g311 ( .A(n_290), .B(n_242), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_287), .A2(n_243), .B(n_253), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_291), .A2(n_259), .B(n_213), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_289), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_309), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_309), .Y(n_316) );
BUFx2_ASAP7_75t_SL g317 ( .A(n_293), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_310), .B(n_276), .Y(n_318) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_296), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_300), .A2(n_269), .B(n_279), .Y(n_320) );
AND2x4_ASAP7_75t_SL g321 ( .A(n_301), .B(n_281), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_300), .A2(n_271), .B(n_289), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_302), .B(n_278), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_299), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_308), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_310), .B(n_270), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_308), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_297), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
AO21x2_ASAP7_75t_L g340 ( .A1(n_306), .A2(n_289), .B(n_270), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_293), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_292), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_311), .B(n_282), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_336), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_331), .B(n_314), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_319), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_333), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_336), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_333), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_329), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_334), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_325), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_334), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_331), .B(n_314), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_334), .B(n_292), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_329), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_342), .B(n_292), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_342), .B(n_292), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_311), .B1(n_304), .B2(n_294), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_342), .B(n_292), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_345), .B(n_311), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_345), .B(n_303), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_341), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_315), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_330), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_315), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_345), .B(n_303), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_316), .B(n_299), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_341), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_330), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_344), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_323), .B(n_303), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_332), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_332), .B(n_298), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_323), .B(n_298), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_335), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_343), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_318), .B(n_304), .Y(n_394) );
INVx2_ASAP7_75t_SL g395 ( .A(n_344), .Y(n_395) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_322), .B(n_298), .Y(n_396) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_322), .B(n_301), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_337), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_322), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_323), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_337), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_364), .B(n_339), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_347), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_398), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_347), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_351), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_323), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_364), .B(n_340), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_368), .B(n_340), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_353), .B(n_340), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_354), .Y(n_413) );
AND2x4_ASAP7_75t_SL g414 ( .A(n_375), .B(n_322), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_387), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_394), .B(n_307), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_354), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_387), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_368), .B(n_339), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_368), .B(n_340), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_371), .B(n_338), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_394), .B(n_324), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_371), .B(n_338), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_350), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_371), .B(n_338), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_373), .B(n_320), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_373), .B(n_320), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_373), .B(n_320), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_361), .B(n_320), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_361), .B(n_346), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_379), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_382), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_353), .B(n_346), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_349), .B(n_324), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_361), .B(n_326), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_355), .B(n_326), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_357), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_392), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_355), .B(n_318), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_358), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_392), .B(n_321), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_352), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_352), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_395), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_375), .B(n_317), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_350), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_374), .B(n_321), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_355), .B(n_317), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_356), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_355), .B(n_321), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_349), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_367), .B(n_312), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_375), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_367), .B(n_237), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_398), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_356), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_372), .B(n_312), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_398), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_356), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_372), .B(n_306), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_374), .B(n_294), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_401), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_374), .B(n_13), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_400), .B(n_272), .C(n_313), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_362), .B(n_13), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_359), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_380), .B(n_301), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_401), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_395), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_362), .B(n_301), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_348), .B(n_15), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_395), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_359), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_359), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_380), .B(n_15), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_348), .B(n_16), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_401), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_399), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_445), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_458), .B(n_375), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_437), .B(n_360), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_407), .B(n_360), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_433), .B(n_399), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_466), .B(n_376), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_458), .B(n_396), .Y(n_490) );
OAI211xp5_ASAP7_75t_L g491 ( .A1(n_416), .A2(n_370), .B(n_397), .C(n_396), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_412), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_413), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_412), .Y(n_494) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_450), .A2(n_370), .B(n_400), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_413), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_426), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_407), .B(n_388), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_443), .B(n_397), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_441), .B(n_363), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_466), .B(n_376), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_408), .B(n_388), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_443), .B(n_376), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_417), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_417), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_472), .B(n_384), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_443), .B(n_384), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_452), .B(n_384), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_408), .B(n_388), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_426), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_472), .B(n_390), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_409), .B(n_393), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_409), .B(n_393), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_472), .B(n_390), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_421), .B(n_380), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_427), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_425), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_421), .B(n_363), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_452), .B(n_391), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_432), .B(n_403), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_432), .B(n_363), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_472), .B(n_390), .Y(n_524) );
AND3x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_252), .C(n_390), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_427), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_403), .B(n_365), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_434), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_444), .B(n_365), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_434), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_435), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_444), .B(n_365), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_436), .B(n_366), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_435), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_452), .B(n_391), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_436), .B(n_366), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_415), .B(n_381), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_468), .B(n_381), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_414), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_480), .B(n_366), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_425), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_439), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_423), .B(n_369), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_419), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_480), .B(n_369), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_418), .B(n_369), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_439), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_405), .B(n_389), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_414), .B(n_389), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_405), .B(n_389), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_438), .B(n_386), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_452), .B(n_386), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_451), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_459), .B(n_17), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_453), .B(n_386), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_406), .B(n_385), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_442), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_438), .B(n_378), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_451), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_478), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_406), .B(n_385), .Y(n_561) );
NOR2x1p5_ASAP7_75t_L g562 ( .A(n_470), .B(n_385), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_422), .B(n_378), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_455), .B(n_378), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_455), .B(n_383), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_422), .B(n_383), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_481), .B(n_17), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_424), .B(n_383), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_474), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_478), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_442), .Y(n_571) );
INVx2_ASAP7_75t_SL g572 ( .A(n_414), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_410), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_481), .B(n_18), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_483), .B(n_429), .Y(n_575) );
NOR2xp33_ASAP7_75t_SL g576 ( .A(n_549), .B(n_449), .Y(n_576) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_490), .A2(n_453), .B1(n_477), .B2(n_447), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_488), .B(n_429), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_485), .B(n_446), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_544), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_484), .B(n_476), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_567), .A2(n_470), .B(n_469), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_521), .B(n_410), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_546), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_516), .B(n_402), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_520), .B(n_430), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_485), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_521), .B(n_430), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_522), .B(n_431), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_562), .A2(n_475), .B1(n_469), .B2(n_448), .Y(n_590) );
AOI21xp33_ASAP7_75t_L g591 ( .A1(n_574), .A2(n_554), .B(n_491), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_487), .B(n_447), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_569), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_516), .B(n_402), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_485), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_544), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_402), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_549), .A2(n_448), .B(n_479), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_520), .B(n_431), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_402), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_487), .B(n_411), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_494), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_493), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_497), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_500), .B(n_420), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_535), .B(n_420), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_496), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_563), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_495), .B(n_411), .C(n_465), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_486), .B(n_420), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_539), .B(n_572), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
INVx4_ASAP7_75t_L g614 ( .A(n_499), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_501), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_555), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_568), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_555), .B(n_420), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_498), .B(n_457), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_511), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_503), .B(n_424), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_498), .B(n_465), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_428), .Y(n_623) );
INVxp67_ASAP7_75t_SL g624 ( .A(n_537), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_495), .A2(n_428), .B(n_440), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_510), .B(n_457), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g627 ( .A1(n_499), .A2(n_461), .B(n_479), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_517), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_526), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_515), .B(n_440), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_528), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_510), .B(n_454), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_513), .A2(n_462), .B1(n_454), .B2(n_471), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_519), .B(n_462), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_524), .B(n_461), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_530), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_489), .B(n_464), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_531), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_513), .B(n_19), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_534), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_514), .A2(n_471), .B(n_464), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_542), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_504), .B(n_482), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_499), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_514), .B(n_482), .Y(n_645) );
OAI22xp33_ASAP7_75t_L g646 ( .A1(n_555), .A2(n_482), .B1(n_473), .B2(n_467), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_547), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_502), .B(n_473), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_557), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_580), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_587), .A2(n_509), .B1(n_519), .B2(n_504), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_583), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_602), .B(n_523), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_601), .B(n_565), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_576), .A2(n_523), .B1(n_509), .B2(n_532), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_593), .B(n_543), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_583), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_602), .B(n_529), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_589), .B(n_533), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_576), .A2(n_508), .B1(n_536), .B2(n_552), .Y(n_660) );
O2A1O1Ixp5_ASAP7_75t_SL g661 ( .A1(n_591), .A2(n_573), .B(n_571), .C(n_561), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_639), .A2(n_550), .B(n_561), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_627), .A2(n_508), .B(n_538), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_633), .B(n_540), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_591), .A2(n_507), .B1(n_552), .B2(n_564), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_592), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_625), .A2(n_545), .B1(n_551), .B2(n_558), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_592), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_596), .B(n_525), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_600), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_603), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_624), .B(n_527), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_596), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_605), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_620), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_577), .A2(n_527), .B(n_548), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_622), .A2(n_548), .A3(n_550), .B1(n_556), .B2(n_570), .C1(n_553), .C2(n_559), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g678 ( .A1(n_616), .A2(n_556), .B1(n_560), .B2(n_541), .C(n_518), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_616), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_618), .A2(n_506), .B(n_505), .C(n_473), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_614), .A2(n_463), .B1(n_460), .B2(n_404), .Y(n_681) );
OAI32xp33_ASAP7_75t_L g682 ( .A1(n_614), .A2(n_463), .A3(n_460), .B1(n_404), .B2(n_467), .Y(n_682) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_590), .A2(n_463), .B(n_460), .C(n_404), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_579), .A2(n_467), .B1(n_252), .B2(n_383), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_628), .Y(n_685) );
AOI322xp5_ASAP7_75t_L g686 ( .A1(n_622), .A2(n_383), .A3(n_20), .B1(n_19), .B2(n_313), .C1(n_295), .C2(n_27), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_629), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_581), .B(n_20), .Y(n_688) );
AOI322xp5_ASAP7_75t_L g689 ( .A1(n_619), .A2(n_626), .A3(n_611), .B1(n_588), .B2(n_634), .C1(n_615), .C2(n_575), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_634), .B(n_383), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_584), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_631), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_641), .B(n_383), .Y(n_693) );
CKINVDCx14_ASAP7_75t_R g694 ( .A(n_612), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_590), .A2(n_295), .B1(n_25), .B2(n_26), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_672), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_689), .B(n_641), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_688), .B(n_582), .C(n_610), .D(n_598), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_663), .A2(n_618), .B1(n_579), .B2(n_644), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_663), .B(n_644), .Y(n_700) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_694), .A2(n_582), .B(n_646), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_665), .A2(n_579), .B1(n_597), .B2(n_594), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_662), .A2(n_606), .B1(n_642), .B2(n_647), .C(n_649), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_660), .B(n_595), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_676), .A2(n_643), .B(n_608), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_677), .B(n_637), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_669), .A2(n_607), .B(n_585), .C(n_621), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_679), .A2(n_632), .B(n_645), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_683), .A2(n_599), .B(n_586), .C(n_635), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_652), .B(n_578), .Y(n_710) );
AOI222xp33_ASAP7_75t_L g711 ( .A1(n_679), .A2(n_640), .B1(n_638), .B2(n_636), .C1(n_604), .C2(n_648), .Y(n_711) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_678), .B(n_617), .C(n_613), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_651), .A2(n_623), .B(n_609), .C(n_630), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_655), .A2(n_24), .B(n_28), .C(n_29), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_673), .A2(n_295), .B1(n_31), .B2(n_32), .C1(n_34), .C2(n_35), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_667), .A2(n_30), .B1(n_37), .B2(n_38), .C(n_40), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_680), .A2(n_41), .B(n_43), .C(n_46), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_657), .B(n_47), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_650), .A2(n_48), .B1(n_52), .B2(n_53), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_656), .A2(n_55), .B1(n_61), .B2(n_64), .C(n_65), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_684), .B(n_66), .C(n_67), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_673), .A2(n_68), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_722) );
AO221x1_ASAP7_75t_L g723 ( .A1(n_681), .A2(n_74), .B1(n_75), .B2(n_76), .C(n_79), .Y(n_723) );
O2A1O1Ixp33_ASAP7_75t_SL g724 ( .A1(n_664), .A2(n_80), .B(n_82), .C(n_83), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_666), .A2(n_84), .B1(n_85), .B2(n_86), .C(n_88), .Y(n_725) );
OAI311xp33_ASAP7_75t_L g726 ( .A1(n_695), .A2(n_89), .A3(n_91), .B1(n_92), .C1(n_94), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_686), .A2(n_95), .B(n_96), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_682), .A2(n_99), .B(n_101), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g729 ( .A1(n_668), .A2(n_218), .B(n_690), .Y(n_729) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_670), .A2(n_218), .B1(n_674), .B2(n_692), .C(n_687), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_693), .A2(n_218), .B(n_691), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_653), .B(n_671), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_675), .B(n_685), .C(n_661), .Y(n_733) );
OAI211xp5_ASAP7_75t_SL g734 ( .A1(n_701), .A2(n_700), .B(n_697), .C(n_727), .Y(n_734) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_722), .B(n_698), .C(n_716), .Y(n_735) );
NAND3x1_ASAP7_75t_L g736 ( .A(n_733), .B(n_705), .C(n_706), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_704), .A2(n_699), .B(n_709), .C(n_713), .Y(n_737) );
NAND3x1_ASAP7_75t_SL g738 ( .A(n_703), .B(n_720), .C(n_723), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_704), .A2(n_696), .B1(n_702), .B2(n_712), .Y(n_739) );
NAND3xp33_ASAP7_75t_SL g740 ( .A(n_737), .B(n_715), .C(n_714), .Y(n_740) );
NAND4xp75_ASAP7_75t_L g741 ( .A(n_736), .B(n_728), .C(n_725), .D(n_730), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_734), .B(n_711), .C(n_718), .Y(n_742) );
AND5x1_ASAP7_75t_L g743 ( .A(n_735), .B(n_707), .C(n_724), .D(n_726), .E(n_721), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_742), .B(n_739), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_740), .Y(n_745) );
NAND5xp2_ASAP7_75t_L g746 ( .A(n_741), .B(n_738), .C(n_717), .D(n_729), .E(n_731), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_745), .B(n_732), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_744), .Y(n_748) );
OR2x6_ASAP7_75t_L g749 ( .A(n_748), .B(n_746), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_747), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_750), .B(n_748), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_751), .A2(n_749), .B(n_748), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_752), .A2(n_719), .B(n_708), .Y(n_753) );
OA22x2_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_743), .B1(n_710), .B2(n_654), .Y(n_754) );
AOI21xp33_ASAP7_75t_L g755 ( .A1(n_754), .A2(n_658), .B(n_659), .Y(n_755) );
endmodule