module fake_jpeg_24406_n_305 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_181;
wire n_26;
wire n_38;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_282;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_39),
.B(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_54),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_28),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_64),
.Y(n_92)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_52),
.B1(n_32),
.B2(n_36),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_33),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_50),
.B1(n_40),
.B2(n_51),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_17),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_86),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_87),
.B1(n_96),
.B2(n_64),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_65),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_72),
.Y(n_122)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_119),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_68),
.B1(n_55),
.B2(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_112),
.B1(n_73),
.B2(n_37),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_65),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_117),
.Y(n_138)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_108),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_74),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_55),
.B1(n_36),
.B2(n_37),
.Y(n_112)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_65),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_97),
.B1(n_98),
.B2(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_122),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_129),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_100),
.B1(n_80),
.B2(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_133),
.B1(n_137),
.B2(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_117),
.B(n_109),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_144),
.B(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_80),
.B1(n_79),
.B2(n_60),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_101),
.B(n_79),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_140),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_90),
.B1(n_75),
.B2(n_42),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_61),
.C(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_146),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_75),
.B1(n_41),
.B2(n_77),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_17),
.B(n_13),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_61),
.B(n_88),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_88),
.B1(n_71),
.B2(n_77),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_111),
.B1(n_121),
.B2(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_152),
.Y(n_178)
);

NAND2x1p5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_167),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_173),
.B1(n_175),
.B2(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_R g162 ( 
.A(n_138),
.B(n_121),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_130),
.C(n_140),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_131),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_165),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_113),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_85),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_69),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_69),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_139),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_81),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_99),
.C(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_120),
.B1(n_108),
.B2(n_106),
.Y(n_175)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_187),
.C(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_142),
.B1(n_161),
.B2(n_162),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_184),
.B1(n_188),
.B2(n_198),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_143),
.B1(n_128),
.B2(n_126),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_144),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_120),
.B1(n_113),
.B2(n_108),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_106),
.B1(n_104),
.B2(n_102),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_99),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_169),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_135),
.B1(n_104),
.B2(n_149),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_13),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_13),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_160),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_173),
.B1(n_175),
.B2(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_213),
.B1(n_214),
.B2(n_184),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_207),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_218),
.C(n_219),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_176),
.B(n_18),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_135),
.B1(n_16),
.B2(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_16),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_53),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_16),
.B1(n_21),
.B2(n_24),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_24),
.B1(n_26),
.B2(n_53),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_15),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_195),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_27),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_190),
.C(n_183),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_238),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_215),
.A2(n_192),
.B1(n_187),
.B2(n_188),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_230),
.B1(n_217),
.B2(n_206),
.Y(n_246)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_177),
.B(n_186),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_240),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_233),
.C(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_203),
.A2(n_186),
.B1(n_23),
.B2(n_18),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_53),
.C(n_38),
.Y(n_233)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_38),
.C(n_34),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_210),
.B(n_34),
.CI(n_20),
.CON(n_238),
.SN(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_26),
.B(n_25),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_38),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_229),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_218),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_252),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_22),
.C(n_20),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_236),
.C(n_225),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_27),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_222),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_263),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_238),
.C(n_12),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_11),
.B(n_1),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_22),
.C(n_20),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_22),
.C(n_19),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_11),
.B(n_1),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_243),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_27),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_269),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_27),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_274),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_277),
.Y(n_290)
);

OAI221xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_254),
.B1(n_243),
.B2(n_248),
.C(n_253),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_3),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_257),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_22),
.B1(n_19),
.B2(n_2),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_265),
.C(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_27),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_281),
.A2(n_282),
.B(n_1),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_0),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_259),
.C(n_2),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_288),
.C(n_7),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_289),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_2),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_291),
.B(n_6),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_275),
.C(n_278),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_7),
.C(n_8),
.Y(n_296)
);

AOI21xp33_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_7),
.B(n_8),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_298),
.A2(n_285),
.B(n_297),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_299),
.B(n_293),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_285),
.C(n_9),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_8),
.B(n_9),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_9),
.B(n_10),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_9),
.B(n_10),
.Y(n_305)
);


endmodule