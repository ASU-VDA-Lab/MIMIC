module real_jpeg_13473_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_42),
.B1(n_64),
.B2(n_67),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_5),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_5),
.A2(n_57),
.B1(n_64),
.B2(n_67),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_28),
.B1(n_32),
.B2(n_57),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_64),
.B1(n_67),
.B2(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_28),
.B1(n_32),
.B2(n_72),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_8),
.A2(n_64),
.B1(n_67),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_8),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_8),
.A2(n_51),
.B1(n_53),
.B2(n_79),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_79),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_79),
.Y(n_287)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_32),
.B(n_35),
.C(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_10),
.B(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_31),
.B1(n_51),
.B2(n_53),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_10),
.A2(n_88),
.B1(n_117),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_55),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_11),
.A2(n_64),
.B1(n_67),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_11),
.A2(n_51),
.B1(n_53),
.B2(n_81),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_81),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_81),
.Y(n_297)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_13),
.A2(n_46),
.B1(n_51),
.B2(n_53),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_13),
.A2(n_46),
.B1(n_64),
.B2(n_67),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_51),
.B1(n_53),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_14),
.A2(n_28),
.B1(n_32),
.B2(n_69),
.Y(n_247)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_318),
.C(n_322),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_316),
.B(n_320),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_308),
.B(n_315),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_274),
.B(n_305),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_252),
.B(n_273),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_225),
.B(n_251),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_126),
.B(n_204),
.C(n_224),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_99),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_24),
.B(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_73),
.C(n_86),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_25),
.B(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_44),
.C(n_58),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_26)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_31),
.A2(n_36),
.B(n_38),
.Y(n_83)
);

HAxp5_ASAP7_75t_SL g136 ( 
.A(n_31),
.B(n_39),
.CON(n_136),
.SN(n_136)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_31),
.B(n_62),
.C(n_67),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_31),
.B(n_88),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_31),
.B(n_63),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_33),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_33),
.A2(n_40),
.B1(n_108),
.B2(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_33),
.B(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_33),
.A2(n_40),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_33),
.A2(n_40),
.B(n_247),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_37),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_37),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_38),
.B(n_50),
.C(n_51),
.Y(n_137)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_40),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_40),
.B(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_58),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_47),
.A2(n_55),
.B1(n_96),
.B2(n_136),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_47),
.A2(n_112),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_47),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_47),
.A2(n_55),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_47),
.A2(n_55),
.B(n_112),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_48),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_48),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_48),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

OA22x2_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_49),
.A2(n_53),
.B(n_135),
.C(n_137),
.Y(n_134)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_51),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_53),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_68),
.B(n_70),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_59),
.A2(n_143),
.B1(n_145),
.B2(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_59),
.A2(n_145),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_59),
.A2(n_145),
.B1(n_153),
.B2(n_163),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_59),
.A2(n_145),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_59),
.A2(n_70),
.B(n_213),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_59),
.A2(n_68),
.B(n_145),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_63),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

CKINVDCx6p67_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_67),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_73),
.B(n_86),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_80),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_75),
.A2(n_120),
.B(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_75),
.A2(n_76),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_76),
.B(n_139),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_94),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_91),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_88),
.A2(n_117),
.B1(n_168),
.B2(n_176),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_88),
.A2(n_117),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_186),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_94),
.B(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_97),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_114),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_100),
.B(n_115),
.C(n_125),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_113),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_109),
.C(n_113),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_105),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_105),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_105),
.A2(n_269),
.B(n_312),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_111),
.B(n_242),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_116),
.B(n_121),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_170),
.B(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_122),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_123),
.B(n_144),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_199),
.B(n_203),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_154),
.B(n_198),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_149),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_149),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_146),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_140),
.C(n_146),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_138),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B(n_144),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_152),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_193),
.B(n_197),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_182),
.B(n_192),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_171),
.B(n_181),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_164),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_180),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_179),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_188),
.C(n_191),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_196),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_223),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_208),
.C(n_215),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_214),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_214),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_227),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_250),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_235),
.B1(n_248),
.B2(n_249),
.Y(n_228)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_249),
.C(n_250),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_231),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_233),
.Y(n_264)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_231),
.A2(n_264),
.B(n_266),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_240),
.C(n_244),
.Y(n_255)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_288),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_272),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_272),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_271),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_257),
.C(n_263),
.Y(n_303)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_261),
.B(n_262),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_261),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_277),
.C(n_290),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_262),
.B(n_277),
.CI(n_290),
.CON(n_304),
.SN(n_304)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_302),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_291),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_291),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_289),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_285),
.C(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_285),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_295),
.C(n_300),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_289),
.B1(n_294),
.B2(n_301),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_292),
.C(n_301),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_294),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_297),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_314),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_318),
.Y(n_321)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.CI(n_313),
.CON(n_309),
.SN(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);


endmodule