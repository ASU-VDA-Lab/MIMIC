module fake_jpeg_8289_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_66),
.Y(n_71)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_56),
.B1(n_51),
.B2(n_42),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_81),
.B1(n_86),
.B2(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_51),
.B1(n_42),
.B2(n_48),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_90),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_40),
.B1(n_47),
.B2(n_46),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_45),
.C(n_41),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_50),
.B1(n_43),
.B2(n_37),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_105),
.C(n_106),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_100),
.B(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_5),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_36),
.B1(n_10),
.B2(n_11),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_16),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_98),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_111),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_87),
.C(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_100),
.C(n_80),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_20),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_119),
.B(n_24),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_102),
.B(n_26),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_121),
.A2(n_97),
.B(n_27),
.C(n_28),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_R g123 ( 
.A(n_122),
.B(n_101),
.Y(n_123)
);

AOI332xp33_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_105),
.A3(n_93),
.B1(n_104),
.B2(n_99),
.B3(n_103),
.C1(n_77),
.C2(n_94),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_107),
.Y(n_125)
);


endmodule