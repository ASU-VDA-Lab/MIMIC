module fake_jpeg_5146_n_285 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_28),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_57),
.B(n_22),
.C(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_25),
.B1(n_31),
.B2(n_20),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_56),
.B1(n_30),
.B2(n_16),
.Y(n_87)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_32),
.B1(n_22),
.B2(n_26),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_76),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_27),
.B(n_18),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_82),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_37),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_26),
.B1(n_18),
.B2(n_30),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_45),
.B1(n_64),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_98),
.B1(n_105),
.B2(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_68),
.B(n_80),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_37),
.B(n_29),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_47),
.B1(n_65),
.B2(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_51),
.B1(n_66),
.B2(n_60),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_23),
.B(n_19),
.Y(n_133)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_27),
.B1(n_16),
.B2(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_61),
.B1(n_44),
.B2(n_33),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_79),
.B1(n_90),
.B2(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_37),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_106),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_23),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_130),
.B1(n_132),
.B2(n_112),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_71),
.B1(n_86),
.B2(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_128),
.B1(n_129),
.B2(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_86),
.B1(n_44),
.B2(n_33),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_85),
.B1(n_82),
.B2(n_78),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_29),
.B1(n_23),
.B2(n_19),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_99),
.B(n_114),
.Y(n_143)
);

OAI22x1_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_113),
.B1(n_98),
.B2(n_97),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_37),
.B1(n_29),
.B2(n_23),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_92),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_144),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_128),
.B1(n_139),
.B2(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_103),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_150),
.C(n_160),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_153),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_37),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_126),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_102),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_102),
.B(n_92),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_107),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_159),
.B1(n_126),
.B2(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_157),
.Y(n_182)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_95),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_116),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_176),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_188),
.B(n_162),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_115),
.B1(n_78),
.B2(n_0),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_138),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_179),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_160),
.C(n_143),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_119),
.C(n_120),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

AO21x2_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_134),
.B(n_121),
.Y(n_186)
);

OAI22x1_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_147),
.B1(n_155),
.B2(n_146),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_187),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_163),
.B(n_154),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_190),
.A2(n_197),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_193),
.CI(n_6),
.CON(n_226),
.SN(n_226)
);

OAI31xp33_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_169),
.A3(n_167),
.B(n_184),
.Y(n_219)
);

AOI22x1_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_144),
.B1(n_115),
.B2(n_19),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.Y(n_211)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_78),
.B1(n_1),
.B2(n_0),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_175),
.B(n_8),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_168),
.C(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_3),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_168),
.B1(n_188),
.B2(n_171),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_190),
.B1(n_197),
.B2(n_195),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_219),
.C(n_226),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_225),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_177),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_170),
.C(n_179),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.C(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_170),
.C(n_165),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_0),
.C(n_3),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_200),
.B1(n_207),
.B2(n_206),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_5),
.C(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

BUFx12_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_230),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_247)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_193),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_233),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_198),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_15),
.B(n_7),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_9),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_220),
.C(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_242),
.C(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_217),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_240),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_218),
.B1(n_7),
.B2(n_8),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_251),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_259),
.C(n_263),
.Y(n_266)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_233),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_249),
.B(n_239),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_244),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_232),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_270),
.C(n_247),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_247),
.C(n_253),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_263),
.B(n_262),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

AO21x2_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_276),
.B(n_230),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_275),
.C(n_277),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_279),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_239),
.B(n_228),
.C(n_230),
.D(n_12),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_282),
.A2(n_280),
.B(n_11),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_11),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_13),
.Y(n_285)
);


endmodule