module fake_aes_9082_n_1032 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1032);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1032;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_434;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1014;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_478;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_955;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_117), .Y(n_268) );
NOR2xp67_ASAP7_75t_L g269 ( .A(n_204), .B(n_259), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_121), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_95), .Y(n_271) );
CKINVDCx14_ASAP7_75t_R g272 ( .A(n_49), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_42), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_49), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_186), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_151), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_26), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_150), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_245), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_241), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_3), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_18), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_137), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_35), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_172), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_9), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_9), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_163), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_64), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_158), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_101), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_50), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_191), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g298 ( .A(n_224), .Y(n_298) );
CKINVDCx14_ASAP7_75t_R g299 ( .A(n_239), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_223), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_116), .Y(n_301) );
CKINVDCx14_ASAP7_75t_R g302 ( .A(n_66), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_61), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_168), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_112), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_22), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_213), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_91), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_258), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_160), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_155), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_79), .B(n_192), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_179), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_262), .Y(n_314) );
CKINVDCx14_ASAP7_75t_R g315 ( .A(n_228), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_231), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_139), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_5), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_124), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_45), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_29), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_225), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_247), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_6), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_13), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_244), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_8), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_85), .Y(n_328) );
BUFx10_ASAP7_75t_L g329 ( .A(n_185), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_243), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_202), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_161), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_44), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_138), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_38), .B(n_130), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_85), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_127), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_265), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_44), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_112), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_144), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_78), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_110), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_133), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_104), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_198), .Y(n_346) );
CKINVDCx16_ASAP7_75t_R g347 ( .A(n_1), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_36), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_36), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_6), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_235), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_40), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_255), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_193), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_227), .B(n_134), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_152), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_221), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_33), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_132), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_131), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_157), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_196), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_145), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_7), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_238), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_250), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_205), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_226), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_118), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_72), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_101), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_209), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_206), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_136), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_257), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_76), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_240), .Y(n_377) );
INVxp33_ASAP7_75t_SL g378 ( .A(n_249), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_178), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_98), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_167), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_208), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_99), .Y(n_383) );
BUFx10_ASAP7_75t_L g384 ( .A(n_97), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_135), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_38), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_115), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_207), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_216), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_254), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_100), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_105), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_113), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_69), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_13), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_190), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_251), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_80), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_181), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_149), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_212), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_129), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_218), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_166), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_222), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_30), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_73), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_47), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_68), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_68), .Y(n_410) );
BUFx10_ASAP7_75t_L g411 ( .A(n_153), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_187), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_200), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_108), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_102), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_23), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_263), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_253), .Y(n_418) );
BUFx12f_ASAP7_75t_L g419 ( .A(n_329), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_306), .B(n_0), .Y(n_420) );
INVx6_ASAP7_75t_L g421 ( .A(n_329), .Y(n_421) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_273), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_396), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_273), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_308), .B(n_0), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_396), .Y(n_427) );
BUFx12f_ASAP7_75t_L g428 ( .A(n_329), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_272), .B(n_2), .Y(n_429) );
INVx6_ASAP7_75t_L g430 ( .A(n_411), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_270), .A2(n_122), .B(n_120), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_283), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_270), .A2(n_125), .B(n_123), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_289), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_289), .Y(n_435) );
BUFx12f_ASAP7_75t_L g436 ( .A(n_411), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_285), .B(n_4), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_287), .B(n_4), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_295), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_295), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_302), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_302), .A2(n_10), .B1(n_5), .B2(n_7), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_318), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_274), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_311), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_288), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_347), .A2(n_14), .B1(n_11), .B2(n_12), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_318), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_361), .B(n_11), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_358), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_288), .Y(n_453) );
OAI21x1_ASAP7_75t_L g454 ( .A1(n_294), .A2(n_128), .B(n_126), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_294), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_313), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_311), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_448), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx8_ASAP7_75t_L g461 ( .A(n_419), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_448), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_448), .B(n_313), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_442), .B(n_299), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_422), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_419), .B(n_411), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_436), .B(n_358), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_453), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_420), .A2(n_296), .B1(n_301), .B2(n_286), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_453), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_455), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_455), .B(n_314), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_447), .Y(n_474) );
AND2x6_ASAP7_75t_L g475 ( .A(n_420), .B(n_316), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_455), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_456), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
BUFx10_ASAP7_75t_L g479 ( .A(n_421), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_422), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_446), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_456), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_422), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_456), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_431), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_436), .B(n_319), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_447), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_421), .B(n_314), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_430), .B(n_378), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_430), .Y(n_493) );
INVx8_ASAP7_75t_L g494 ( .A(n_461), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_492), .B(n_430), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_476), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_464), .B(n_430), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_464), .B(n_444), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_475), .A2(n_429), .B1(n_426), .B2(n_425), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_458), .A2(n_429), .B(n_454), .C(n_438), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_479), .B(n_428), .Y(n_502) );
OR2x6_ASAP7_75t_L g503 ( .A(n_461), .B(n_428), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_479), .B(n_437), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_461), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_486), .A2(n_454), .B(n_433), .Y(n_506) );
NOR2xp33_ASAP7_75t_SL g507 ( .A(n_461), .B(n_279), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_470), .A2(n_443), .B1(n_281), .B2(n_284), .Y(n_509) );
BUFx8_ASAP7_75t_L g510 ( .A(n_475), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_466), .B(n_451), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_467), .B(n_384), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_468), .B(n_378), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_491), .B(n_337), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_491), .B(n_337), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_462), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_467), .B(n_274), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_475), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_467), .B(n_449), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_475), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_467), .B(n_277), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_468), .B(n_377), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_477), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_475), .B(n_377), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_488), .B(n_423), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_493), .B(n_458), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_475), .B(n_412), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_477), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_481), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_479), .B(n_412), .Y(n_532) );
BUFx8_ASAP7_75t_L g533 ( .A(n_475), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_486), .A2(n_433), .B(n_431), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_493), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_458), .B(n_449), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_486), .B(n_425), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_469), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g539 ( .A(n_471), .B(n_355), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_477), .B(n_298), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_472), .B(n_315), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_463), .B(n_380), .C(n_320), .Y(n_542) );
NOR2xp33_ASAP7_75t_SL g543 ( .A(n_487), .B(n_298), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_487), .B(n_315), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_482), .B(n_384), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_487), .B(n_293), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_484), .B(n_432), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_463), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_489), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_473), .B(n_432), .Y(n_550) );
NAND2xp33_ASAP7_75t_L g551 ( .A(n_473), .B(n_300), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_485), .A2(n_435), .B1(n_440), .B2(n_434), .Y(n_552) );
OR2x6_ASAP7_75t_L g553 ( .A(n_489), .B(n_410), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_489), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_474), .B(n_435), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_474), .A2(n_450), .B1(n_452), .B2(n_445), .C(n_441), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_534), .A2(n_433), .B(n_431), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_534), .A2(n_433), .B(n_335), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_499), .A2(n_368), .B1(n_402), .B2(n_354), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_548), .B(n_277), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_536), .A2(n_406), .B1(n_407), .B2(n_364), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_545), .B(n_406), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_538), .A2(n_292), .B1(n_352), .B2(n_290), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_507), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_531), .Y(n_565) );
INVx3_ASAP7_75t_L g566 ( .A(n_494), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_538), .B(n_407), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_494), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_509), .A2(n_387), .B1(n_408), .B2(n_328), .C(n_336), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_519), .B(n_408), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_514), .B(n_268), .Y(n_571) );
INVx3_ASAP7_75t_SL g572 ( .A(n_503), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_523), .B(n_271), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_503), .Y(n_574) );
AOI33xp33_ASAP7_75t_L g575 ( .A1(n_552), .A2(n_452), .A3(n_348), .B1(n_339), .B2(n_370), .B3(n_369), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_506), .A2(n_276), .B(n_275), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_SL g577 ( .A1(n_546), .A2(n_278), .B(n_291), .C(n_280), .Y(n_577) );
CKINVDCx11_ASAP7_75t_R g578 ( .A(n_521), .Y(n_578) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_516), .B(n_343), .C(n_282), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_514), .B(n_303), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_542), .B(n_305), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_542), .B(n_321), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_506), .A2(n_323), .B(n_297), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_543), .A2(n_324), .B1(n_327), .B2(n_325), .Y(n_584) );
OA22x2_ASAP7_75t_L g585 ( .A1(n_516), .A2(n_395), .B1(n_349), .B2(n_350), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_512), .B(n_345), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_544), .A2(n_307), .B(n_304), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_501), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_541), .A2(n_310), .B(n_309), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
CKINVDCx6p67_ASAP7_75t_R g591 ( .A(n_505), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_515), .B(n_386), .Y(n_592) );
NOR2xp67_ASAP7_75t_L g593 ( .A(n_505), .B(n_12), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_517), .B(n_371), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_539), .B(n_474), .C(n_317), .Y(n_595) );
AOI21x1_ASAP7_75t_L g596 ( .A1(n_526), .A2(n_478), .B(n_460), .Y(n_596) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_513), .B(n_15), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_550), .Y(n_598) );
AOI21x1_ASAP7_75t_L g599 ( .A1(n_529), .A2(n_478), .B(n_460), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_527), .B(n_391), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_502), .B(n_392), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_552), .A2(n_394), .B1(n_409), .B2(n_393), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_415), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_510), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_528), .A2(n_306), .B(n_340), .C(n_333), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_497), .B(n_416), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g607 ( .A1(n_508), .A2(n_326), .B(n_322), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g608 ( .A1(n_528), .A2(n_342), .B(n_398), .C(n_340), .Y(n_608) );
OA22x2_ASAP7_75t_L g609 ( .A1(n_540), .A2(n_414), .B1(n_410), .B2(n_331), .Y(n_609) );
BUFx12f_ASAP7_75t_L g610 ( .A(n_533), .Y(n_610) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_522), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_495), .A2(n_332), .B(n_330), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_524), .A2(n_341), .B(n_338), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_511), .B(n_398), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_504), .A2(n_351), .B(n_346), .Y(n_615) );
AO21x2_ASAP7_75t_L g616 ( .A1(n_556), .A2(n_357), .B(n_356), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_518), .A2(n_360), .B(n_359), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_547), .B(n_414), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_496), .Y(n_619) );
BUFx2_ASAP7_75t_L g620 ( .A(n_553), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_551), .A2(n_363), .B(n_362), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_532), .A2(n_367), .B(n_365), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_SL g623 ( .A1(n_535), .A2(n_373), .B(n_374), .C(n_372), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_553), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_549), .A2(n_382), .B(n_379), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_553), .A2(n_312), .B1(n_389), .B2(n_388), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_L g628 ( .A1(n_525), .A2(n_399), .B(n_401), .C(n_397), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_530), .A2(n_405), .B(n_417), .C(n_403), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_554), .A2(n_385), .B(n_366), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_534), .A2(n_385), .B(n_366), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_534), .A2(n_404), .B(n_400), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_494), .Y(n_633) );
NOR2xp33_ASAP7_75t_SL g634 ( .A(n_494), .B(n_344), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_534), .A2(n_404), .B(n_400), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_536), .A2(n_383), .B1(n_376), .B2(n_447), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_534), .A2(n_483), .B(n_480), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_498), .B(n_334), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_548), .B(n_353), .Y(n_639) );
NOR2x1_ASAP7_75t_SL g640 ( .A(n_503), .B(n_316), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_548), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_548), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_548), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g644 ( .A(n_531), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_548), .B(n_375), .Y(n_645) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_494), .B(n_381), .Y(n_646) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_506), .A2(n_490), .B(n_269), .Y(n_647) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_534), .A2(n_474), .B(n_413), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_537), .A2(n_418), .B(n_390), .C(n_427), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_537), .A2(n_418), .B(n_390), .C(n_383), .Y(n_650) );
AO31x2_ASAP7_75t_L g651 ( .A1(n_558), .A2(n_457), .A3(n_447), .B(n_439), .Y(n_651) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_631), .A2(n_635), .A3(n_632), .B(n_648), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_568), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_598), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_588), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_637), .A2(n_465), .B(n_424), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_565), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_642), .B(n_383), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_583), .A2(n_465), .B(n_424), .Y(n_659) );
AO31x2_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_424), .A3(n_465), .B(n_18), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_587), .A2(n_424), .B(n_19), .C(n_16), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_561), .B(n_17), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_641), .B(n_17), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_573), .B(n_20), .C(n_21), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_644), .Y(n_665) );
INVx2_ASAP7_75t_SL g666 ( .A(n_572), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_643), .B(n_20), .Y(n_667) );
NAND2xp33_ASAP7_75t_R g668 ( .A(n_604), .B(n_22), .Y(n_668) );
AO31x2_ASAP7_75t_L g669 ( .A1(n_605), .A2(n_26), .A3(n_24), .B(n_25), .Y(n_669) );
OA21x2_ASAP7_75t_L g670 ( .A1(n_596), .A2(n_141), .B(n_140), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_570), .B(n_25), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_619), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_591), .B(n_27), .Y(n_673) );
NAND2x1_ASAP7_75t_L g674 ( .A(n_566), .B(n_142), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_569), .B(n_27), .Y(n_675) );
INVxp67_ASAP7_75t_SL g676 ( .A(n_559), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_566), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_578), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_613), .A2(n_146), .B(n_143), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_608), .A2(n_30), .B(n_28), .C(n_29), .Y(n_680) );
OAI21x1_ASAP7_75t_L g681 ( .A1(n_599), .A2(n_148), .B(n_147), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_610), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_636), .B(n_28), .C(n_31), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_620), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_594), .A2(n_156), .B(n_154), .Y(n_685) );
AO31x2_ASAP7_75t_L g686 ( .A1(n_649), .A2(n_40), .A3(n_37), .B(n_39), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_575), .B(n_37), .Y(n_687) );
AO31x2_ASAP7_75t_L g688 ( .A1(n_626), .A2(n_42), .A3(n_39), .B(n_41), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_592), .A2(n_162), .B(n_159), .Y(n_689) );
NOR2xp67_ASAP7_75t_SL g690 ( .A(n_633), .B(n_43), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_567), .B(n_560), .Y(n_691) );
AOI221x1_ASAP7_75t_L g692 ( .A1(n_626), .A2(n_46), .B1(n_47), .B2(n_48), .C(n_51), .Y(n_692) );
AO21x1_ASAP7_75t_L g693 ( .A1(n_630), .A2(n_165), .B(n_164), .Y(n_693) );
O2A1O1Ixp5_ASAP7_75t_SL g694 ( .A1(n_564), .A2(n_607), .B(n_602), .C(n_614), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_586), .B(n_51), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_612), .A2(n_52), .B(n_53), .C(n_54), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_624), .A2(n_52), .B1(n_53), .B2(n_54), .Y(n_697) );
OAI21x1_ASAP7_75t_L g698 ( .A1(n_625), .A2(n_170), .B(n_169), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_627), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_609), .A2(n_173), .B(n_171), .Y(n_700) );
NOR2xp67_ASAP7_75t_L g701 ( .A(n_595), .B(n_174), .Y(n_701) );
OAI21x1_ASAP7_75t_L g702 ( .A1(n_609), .A2(n_176), .B(n_175), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_571), .A2(n_180), .B(n_177), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_628), .A2(n_55), .B(n_56), .C(n_57), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_563), .B(n_56), .Y(n_705) );
AO21x2_ASAP7_75t_L g706 ( .A1(n_593), .A2(n_183), .B(n_182), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_580), .B(n_58), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_638), .B(n_58), .Y(n_708) );
NAND2xp33_ASAP7_75t_L g709 ( .A(n_590), .B(n_184), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_618), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_617), .A2(n_189), .B(n_188), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_616), .Y(n_712) );
OR2x6_ASAP7_75t_L g713 ( .A(n_574), .B(n_59), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_629), .A2(n_59), .B(n_60), .C(n_61), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_615), .A2(n_195), .B(n_194), .Y(n_715) );
AO31x2_ASAP7_75t_L g716 ( .A1(n_602), .A2(n_60), .A3(n_62), .B(n_63), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_621), .A2(n_622), .B(n_582), .Y(n_717) );
BUFx3_ASAP7_75t_L g718 ( .A(n_601), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_606), .Y(n_719) );
OA21x2_ASAP7_75t_L g720 ( .A1(n_600), .A2(n_199), .B(n_197), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g721 ( .A1(n_584), .A2(n_63), .B(n_64), .Y(n_721) );
AO31x2_ASAP7_75t_L g722 ( .A1(n_603), .A2(n_65), .A3(n_66), .B(n_67), .Y(n_722) );
OA21x2_ASAP7_75t_L g723 ( .A1(n_597), .A2(n_203), .B(n_201), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_562), .B(n_70), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_623), .Y(n_725) );
AO31x2_ASAP7_75t_L g726 ( .A1(n_640), .A2(n_71), .A3(n_72), .B(n_73), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_579), .A2(n_71), .B1(n_74), .B2(n_75), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_590), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_590), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_611), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_581), .B(n_74), .Y(n_731) );
AOI21xp5_ASAP7_75t_SL g732 ( .A1(n_611), .A2(n_211), .B(n_210), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_577), .A2(n_219), .B(n_266), .Y(n_733) );
AO31x2_ASAP7_75t_L g734 ( .A1(n_639), .A2(n_75), .A3(n_76), .B(n_77), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_585), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_585), .A2(n_215), .B(n_264), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_645), .B(n_77), .Y(n_737) );
AND3x4_ASAP7_75t_L g738 ( .A(n_634), .B(n_646), .C(n_81), .Y(n_738) );
AND2x4_ASAP7_75t_L g739 ( .A(n_634), .B(n_80), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_605), .A2(n_82), .B(n_83), .C(n_84), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_589), .A2(n_82), .B(n_83), .C(n_84), .Y(n_741) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_568), .Y(n_742) );
AOI31xp67_ASAP7_75t_L g743 ( .A1(n_609), .A2(n_220), .A3(n_261), .B(n_260), .Y(n_743) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_576), .A2(n_214), .B(n_256), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_570), .A2(n_86), .B(n_87), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_598), .Y(n_746) );
AOI21x1_ASAP7_75t_L g747 ( .A1(n_557), .A2(n_267), .B(n_252), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_598), .B(n_87), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_573), .B(n_88), .C(n_89), .Y(n_749) );
OA21x2_ASAP7_75t_L g750 ( .A1(n_576), .A2(n_248), .B(n_246), .Y(n_750) );
AOI31xp67_ASAP7_75t_L g751 ( .A1(n_609), .A2(n_242), .A3(n_237), .B(n_236), .Y(n_751) );
AOI21x1_ASAP7_75t_L g752 ( .A1(n_656), .A2(n_234), .B(n_233), .Y(n_752) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_657), .Y(n_753) );
AO31x2_ASAP7_75t_L g754 ( .A1(n_712), .A2(n_90), .A3(n_91), .B(n_92), .Y(n_754) );
BUFx2_ASAP7_75t_L g755 ( .A(n_665), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_719), .B(n_93), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_682), .Y(n_757) );
BUFx2_ASAP7_75t_L g758 ( .A(n_742), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_659), .A2(n_94), .B(n_96), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_699), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_678), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_655), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_668), .Y(n_763) );
OR2x2_ASAP7_75t_L g764 ( .A(n_718), .B(n_103), .Y(n_764) );
BUFx3_ASAP7_75t_L g765 ( .A(n_653), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_651), .Y(n_766) );
AO31x2_ASAP7_75t_L g767 ( .A1(n_693), .A2(n_106), .A3(n_107), .B(n_108), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_651), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_653), .B(n_107), .Y(n_769) );
OA21x2_ASAP7_75t_L g770 ( .A1(n_681), .A2(n_109), .B(n_110), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_710), .B(n_111), .Y(n_771) );
BUFx8_ASAP7_75t_L g772 ( .A(n_666), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_676), .B(n_113), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_748), .Y(n_774) );
AO21x2_ASAP7_75t_L g775 ( .A1(n_725), .A2(n_114), .B(n_115), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_672), .Y(n_776) );
INVx8_ASAP7_75t_L g777 ( .A(n_713), .Y(n_777) );
AO21x2_ASAP7_75t_L g778 ( .A1(n_725), .A2(n_119), .B(n_747), .Y(n_778) );
AOI21x1_ASAP7_75t_L g779 ( .A1(n_670), .A2(n_701), .B(n_720), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_662), .B(n_705), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_717), .A2(n_707), .B(n_695), .Y(n_781) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_739), .B(n_690), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_729), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_691), .B(n_724), .Y(n_784) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_687), .A2(n_675), .B(n_731), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_663), .Y(n_786) );
OA21x2_ASAP7_75t_L g787 ( .A1(n_700), .A2(n_702), .B(n_698), .Y(n_787) );
INVx4_ASAP7_75t_L g788 ( .A(n_729), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_673), .B(n_735), .Y(n_789) );
O2A1O1Ixp33_ASAP7_75t_L g790 ( .A1(n_741), .A2(n_696), .B(n_714), .C(n_661), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_729), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_671), .A2(n_737), .B(n_708), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_667), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_652), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_722), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_740), .A2(n_683), .B(n_689), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_727), .B(n_677), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_728), .A2(n_730), .B(n_674), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_722), .Y(n_799) );
AND2x4_ASAP7_75t_L g800 ( .A(n_736), .B(n_683), .Y(n_800) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_744), .A2(n_750), .B(n_703), .Y(n_801) );
A2O1A1Ixp33_ASAP7_75t_L g802 ( .A1(n_704), .A2(n_664), .B(n_749), .C(n_745), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_726), .B(n_658), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_722), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_716), .Y(n_805) );
OAI21x1_ASAP7_75t_L g806 ( .A1(n_723), .A2(n_685), .B(n_715), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_733), .A2(n_711), .B(n_679), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_684), .B(n_697), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_692), .A2(n_751), .B(n_743), .Y(n_809) );
OAI21x1_ASAP7_75t_L g810 ( .A1(n_732), .A2(n_706), .B(n_709), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_660), .A2(n_669), .B(n_686), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_716), .B(n_688), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_734), .B(n_688), .Y(n_813) );
BUFx3_ASAP7_75t_L g814 ( .A(n_734), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_654), .B(n_746), .Y(n_815) );
NOR2xp67_ASAP7_75t_L g816 ( .A(n_657), .B(n_610), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_654), .B(n_521), .Y(n_817) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_742), .Y(n_818) );
A2O1A1Ixp33_ASAP7_75t_L g819 ( .A1(n_721), .A2(n_680), .B(n_740), .C(n_704), .Y(n_819) );
INVx3_ASAP7_75t_L g820 ( .A(n_742), .Y(n_820) );
AO21x2_ASAP7_75t_L g821 ( .A1(n_712), .A2(n_576), .B(n_647), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_651), .Y(n_822) );
NAND2x1p5_ASAP7_75t_L g823 ( .A(n_742), .B(n_568), .Y(n_823) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_682), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_694), .A2(n_576), .B(n_500), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_654), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_651), .Y(n_827) );
OAI21xp5_ASAP7_75t_L g828 ( .A1(n_694), .A2(n_576), .B(n_500), .Y(n_828) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_656), .A2(n_557), .B(n_558), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_654), .B(n_746), .Y(n_830) );
BUFx2_ASAP7_75t_SL g831 ( .A(n_682), .Y(n_831) );
NAND2x1p5_ASAP7_75t_L g832 ( .A(n_742), .B(n_568), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_676), .A2(n_738), .B1(n_739), .B2(n_559), .Y(n_833) );
AO21x2_ASAP7_75t_L g834 ( .A1(n_811), .A2(n_829), .B(n_813), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g835 ( .A1(n_819), .A2(n_802), .B(n_792), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_815), .B(n_760), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_830), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_780), .B(n_817), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_815), .B(n_776), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_766), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_768), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_826), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_762), .Y(n_843) );
OA21x2_ASAP7_75t_L g844 ( .A1(n_801), .A2(n_812), .B(n_813), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_756), .Y(n_845) );
BUFx3_ASAP7_75t_L g846 ( .A(n_772), .Y(n_846) );
INVx3_ASAP7_75t_L g847 ( .A(n_788), .Y(n_847) );
BUFx2_ASAP7_75t_SL g848 ( .A(n_816), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_771), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_784), .B(n_764), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_822), .Y(n_851) );
INVxp67_ASAP7_75t_L g852 ( .A(n_831), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_827), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_769), .Y(n_854) );
AO21x2_ASAP7_75t_L g855 ( .A1(n_825), .A2(n_828), .B(n_812), .Y(n_855) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_819), .A2(n_802), .B(n_792), .Y(n_856) );
AND2x4_ASAP7_75t_L g857 ( .A(n_791), .B(n_788), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_769), .Y(n_858) );
INVx8_ASAP7_75t_L g859 ( .A(n_777), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_754), .Y(n_860) );
AND2x4_ASAP7_75t_L g861 ( .A(n_791), .B(n_818), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_754), .Y(n_862) );
AO21x2_ASAP7_75t_L g863 ( .A1(n_779), .A2(n_781), .B(n_804), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_808), .B(n_833), .Y(n_864) );
AND2x4_ASAP7_75t_L g865 ( .A(n_818), .B(n_820), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_783), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_785), .B(n_773), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_794), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_789), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_795), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_799), .Y(n_871) );
OA21x2_ASAP7_75t_L g872 ( .A1(n_781), .A2(n_805), .B(n_806), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_833), .B(n_774), .Y(n_873) );
AND2x4_ASAP7_75t_L g874 ( .A(n_818), .B(n_820), .Y(n_874) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_814), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_823), .Y(n_876) );
AOI21x1_ASAP7_75t_L g877 ( .A1(n_800), .A2(n_809), .B(n_810), .Y(n_877) );
INVx1_ASAP7_75t_SL g878 ( .A(n_755), .Y(n_878) );
INVx3_ASAP7_75t_L g879 ( .A(n_818), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_765), .B(n_797), .Y(n_880) );
INVx3_ASAP7_75t_L g881 ( .A(n_832), .Y(n_881) );
BUFx2_ASAP7_75t_L g882 ( .A(n_758), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_775), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_821), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_782), .Y(n_885) );
OR2x6_ASAP7_75t_L g886 ( .A(n_824), .B(n_757), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_786), .B(n_793), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_759), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_843), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_864), .B(n_767), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_839), .B(n_767), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_873), .B(n_767), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_835), .B(n_803), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_856), .B(n_800), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_870), .Y(n_895) );
HB1xp67_ASAP7_75t_L g896 ( .A(n_836), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_868), .Y(n_897) );
BUFx2_ASAP7_75t_L g898 ( .A(n_841), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_887), .Y(n_899) );
INVx2_ASAP7_75t_SL g900 ( .A(n_857), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_869), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_871), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_850), .B(n_763), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_867), .B(n_809), .Y(n_904) );
INVx5_ASAP7_75t_SL g905 ( .A(n_886), .Y(n_905) );
NAND2xp5_ASAP7_75t_SL g906 ( .A(n_847), .B(n_753), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_851), .B(n_778), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_842), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_838), .B(n_778), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_851), .B(n_770), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_875), .Y(n_911) );
BUFx2_ASAP7_75t_L g912 ( .A(n_875), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_837), .B(n_790), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_866), .B(n_796), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_836), .Y(n_915) );
NAND2xp5_ASAP7_75t_SL g916 ( .A(n_847), .B(n_761), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_840), .B(n_787), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_880), .B(n_798), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_882), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_878), .B(n_752), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_853), .B(n_807), .Y(n_921) );
NAND2x1_ASAP7_75t_L g922 ( .A(n_885), .B(n_879), .Y(n_922) );
INVx2_ASAP7_75t_SL g923 ( .A(n_857), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_884), .Y(n_924) );
A2O1A1Ixp33_ASAP7_75t_SL g925 ( .A1(n_847), .A2(n_852), .B(n_883), .C(n_854), .Y(n_925) );
BUFx3_ASAP7_75t_L g926 ( .A(n_846), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_855), .B(n_860), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_862), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_928), .Y(n_929) );
INVx3_ASAP7_75t_R g930 ( .A(n_898), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_924), .Y(n_931) );
AND2x4_ASAP7_75t_L g932 ( .A(n_894), .B(n_834), .Y(n_932) );
BUFx2_ASAP7_75t_L g933 ( .A(n_898), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_899), .B(n_845), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_911), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_904), .B(n_855), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_893), .B(n_844), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_893), .B(n_844), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_891), .B(n_844), .Y(n_939) );
INVx2_ASAP7_75t_SL g940 ( .A(n_912), .Y(n_940) );
AND2x4_ASAP7_75t_L g941 ( .A(n_918), .B(n_877), .Y(n_941) );
BUFx3_ASAP7_75t_L g942 ( .A(n_900), .Y(n_942) );
NAND2x1_ASAP7_75t_L g943 ( .A(n_918), .B(n_885), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_895), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_919), .Y(n_945) );
INVx5_ASAP7_75t_L g946 ( .A(n_905), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_896), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_902), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_890), .B(n_863), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_901), .B(n_849), .Y(n_950) );
NAND2x1p5_ASAP7_75t_L g951 ( .A(n_922), .B(n_858), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_914), .B(n_888), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_890), .B(n_863), .Y(n_953) );
INVxp67_ASAP7_75t_L g954 ( .A(n_926), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_927), .B(n_872), .Y(n_955) );
INVx2_ASAP7_75t_SL g956 ( .A(n_923), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_929), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_937), .B(n_938), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_929), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_944), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_944), .Y(n_961) );
AND2x2_ASAP7_75t_L g962 ( .A(n_938), .B(n_907), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_945), .B(n_954), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_948), .Y(n_964) );
AND2x2_ASAP7_75t_L g965 ( .A(n_936), .B(n_910), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_933), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_948), .Y(n_967) );
NAND2xp33_ASAP7_75t_SL g968 ( .A(n_930), .B(n_915), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_934), .B(n_889), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_949), .B(n_917), .Y(n_970) );
INVx2_ASAP7_75t_L g971 ( .A(n_931), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_950), .Y(n_972) );
AND2x2_ASAP7_75t_L g973 ( .A(n_953), .B(n_917), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_933), .Y(n_974) );
AND2x4_ASAP7_75t_L g975 ( .A(n_941), .B(n_921), .Y(n_975) );
AND2x4_ASAP7_75t_L g976 ( .A(n_941), .B(n_897), .Y(n_976) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_966), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_957), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_957), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_971), .Y(n_980) );
INVxp67_ASAP7_75t_L g981 ( .A(n_963), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_959), .Y(n_982) );
INVx3_ASAP7_75t_L g983 ( .A(n_976), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_959), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_971), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_972), .B(n_955), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_960), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_958), .B(n_939), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_961), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_965), .B(n_947), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_964), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_958), .B(n_939), .Y(n_992) );
INVx2_ASAP7_75t_L g993 ( .A(n_967), .Y(n_993) );
BUFx2_ASAP7_75t_L g994 ( .A(n_968), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_970), .B(n_932), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_970), .B(n_932), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_973), .B(n_932), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_980), .Y(n_998) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_977), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_991), .B(n_973), .Y(n_1000) );
O2A1O1Ixp33_ASAP7_75t_L g1001 ( .A1(n_981), .A2(n_886), .B(n_916), .C(n_925), .Y(n_1001) );
OAI21xp33_ASAP7_75t_L g1002 ( .A1(n_986), .A2(n_974), .B(n_962), .Y(n_1002) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_994), .A2(n_906), .B(n_943), .Y(n_1003) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_983), .B(n_975), .Y(n_1004) );
NAND2x1_ASAP7_75t_L g1005 ( .A(n_983), .B(n_935), .Y(n_1005) );
INVxp67_ASAP7_75t_L g1006 ( .A(n_990), .Y(n_1006) );
AOI21xp33_ASAP7_75t_L g1007 ( .A1(n_1001), .A2(n_920), .B(n_903), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_1002), .A2(n_969), .B1(n_996), .B2(n_995), .C(n_997), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1009 ( .A1(n_1006), .A2(n_987), .B1(n_988), .B2(n_992), .C(n_989), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1010 ( .A1(n_1005), .A2(n_942), .B1(n_956), .B2(n_946), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_1003), .A2(n_940), .B(n_993), .Y(n_1011) );
INVxp67_ASAP7_75t_L g1012 ( .A(n_999), .Y(n_1012) );
AOI21xp5_ASAP7_75t_L g1013 ( .A1(n_1011), .A2(n_1004), .B(n_1000), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1012), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1009), .B(n_998), .Y(n_1015) );
O2A1O1Ixp33_ASAP7_75t_L g1016 ( .A1(n_1014), .A2(n_1007), .B(n_1010), .C(n_1008), .Y(n_1016) );
NOR2x1_ASAP7_75t_L g1017 ( .A(n_1013), .B(n_848), .Y(n_1017) );
O2A1O1Ixp5_ASAP7_75t_L g1018 ( .A1(n_1015), .A2(n_985), .B(n_913), .C(n_941), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_1017), .B(n_859), .Y(n_1019) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_1016), .B(n_978), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_1018), .A2(n_951), .B(n_909), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1020), .B(n_1019), .Y(n_1022) );
A2O1A1Ixp33_ASAP7_75t_L g1023 ( .A1(n_1021), .A2(n_946), .B(n_942), .C(n_908), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1022), .Y(n_1024) );
INVx2_ASAP7_75t_SL g1025 ( .A(n_1023), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1024), .Y(n_1026) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_1026), .A2(n_1025), .B(n_951), .Y(n_1027) );
NAND3xp33_ASAP7_75t_SL g1028 ( .A(n_1027), .B(n_892), .C(n_952), .Y(n_1028) );
AOI21xp5_ASAP7_75t_L g1029 ( .A1(n_1028), .A2(n_876), .B(n_984), .Y(n_1029) );
OAI21xp5_ASAP7_75t_L g1030 ( .A1(n_1029), .A2(n_861), .B(n_881), .Y(n_1030) );
OAI21xp5_ASAP7_75t_L g1031 ( .A1(n_1030), .A2(n_865), .B(n_874), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_1031), .A2(n_984), .B1(n_982), .B2(n_979), .Y(n_1032) );
endmodule