module fake_ariane_2385_n_191 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_191);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_191;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_128;
wire n_105;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_146;
wire n_80;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_2),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_R g70 ( 
.A(n_38),
.B(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_37),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_9),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g74 ( 
.A(n_32),
.B(n_10),
.CON(n_74),
.SN(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_46),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_53),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_43),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_52),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

AOI221xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.C(n_44),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_56),
.B(n_57),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_65),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_71),
.B1(n_74),
.B2(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_65),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_56),
.B(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_72),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_73),
.B(n_58),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_91),
.B(n_89),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_81),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_74),
.B1(n_81),
.B2(n_82),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

AOI222xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_74),
.B1(n_81),
.B2(n_82),
.C1(n_103),
.C2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_79),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_98),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_110),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OR2x6_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NOR2x1p5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_110),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_116),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_114),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_117),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_104),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_118),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_71),
.Y(n_136)
);

AOI211xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_35),
.B(n_40),
.C(n_36),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_106),
.B1(n_109),
.B2(n_107),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_94),
.B(n_106),
.Y(n_139)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_38),
.B1(n_42),
.B2(n_49),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_109),
.B1(n_107),
.B2(n_92),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_58),
.C(n_70),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_133),
.B1(n_131),
.B2(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_131),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_50),
.B1(n_51),
.B2(n_98),
.C(n_91),
.Y(n_146)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_124),
.Y(n_147)
);

AOI211xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_75),
.B(n_87),
.C(n_86),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_75),
.B1(n_132),
.B2(n_87),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_75),
.B1(n_87),
.B2(n_85),
.C(n_86),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_132),
.B1(n_127),
.B2(n_125),
.Y(n_151)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_59),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_66),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_59),
.C(n_62),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_89),
.C(n_85),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_99),
.B(n_93),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_127),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_11),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_68),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_65),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

NOR2xp67_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_105),
.Y(n_164)
);

NOR4xp25_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_146),
.C(n_66),
.D(n_68),
.Y(n_165)
);

NOR2x1p5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_64),
.Y(n_166)
);

NOR4xp75_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_167)
);

OAI221xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_64),
.B1(n_95),
.B2(n_100),
.C(n_80),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

OAI221xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_64),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_159),
.A3(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_95),
.B1(n_77),
.B2(n_90),
.C(n_18),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_12),
.A3(n_19),
.B1(n_100),
.B2(n_99),
.C1(n_93),
.C2(n_80),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_99),
.A3(n_80),
.B1(n_90),
.B2(n_77),
.C1(n_94),
.C2(n_27),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_80),
.A3(n_22),
.B1(n_23),
.B2(n_25),
.C1(n_26),
.C2(n_30),
.Y(n_176)
);

OAI221xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_162),
.B1(n_168),
.B2(n_164),
.C(n_166),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_173),
.B1(n_164),
.B2(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_175),
.B(n_105),
.C(n_20),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_171),
.A2(n_105),
.B1(n_92),
.B2(n_63),
.Y(n_182)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_105),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_105),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_L g190 ( 
.A(n_188),
.B(n_184),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B1(n_185),
.B2(n_186),
.C(n_189),
.Y(n_191)
);


endmodule