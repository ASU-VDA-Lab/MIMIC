module real_aes_8424_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_329;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_316;
wire n_746;
wire n_532;
wire n_656;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_0), .A2(n_239), .B1(n_400), .B2(n_402), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_1), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_2), .A2(n_222), .B1(n_731), .B2(n_764), .Y(n_763) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_3), .B(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_4), .A2(n_175), .B1(n_466), .B2(n_469), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_5), .A2(n_55), .B1(n_460), .B2(n_582), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_6), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_7), .A2(n_244), .B1(n_332), .B2(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_8), .Y(n_570) );
INVx1_ASAP7_75t_L g717 ( .A(n_9), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g813 ( .A1(n_10), .A2(n_27), .B1(n_232), .B2(n_428), .C1(n_698), .C2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_11), .A2(n_121), .B1(n_358), .B2(n_473), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_12), .A2(n_171), .B1(n_412), .B2(n_567), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_13), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_14), .B(n_584), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_15), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_16), .A2(n_70), .B1(n_511), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_17), .A2(n_152), .B1(n_539), .B2(n_564), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_18), .A2(n_205), .B1(n_397), .B2(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_19), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_20), .A2(n_389), .B1(n_441), .B2(n_442), .Y(n_388) );
INVx1_ASAP7_75t_L g441 ( .A(n_20), .Y(n_441) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_21), .B(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_22), .A2(n_72), .B1(n_355), .B2(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g681 ( .A(n_23), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_24), .A2(n_85), .B1(n_464), .B2(n_814), .Y(n_846) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_25), .A2(n_77), .B1(n_308), .B2(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g832 ( .A(n_25), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_26), .A2(n_148), .B1(n_401), .B2(n_415), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_28), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g621 ( .A1(n_29), .A2(n_194), .B1(n_593), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g547 ( .A(n_30), .Y(n_547) );
AOI222xp33_ASAP7_75t_L g569 ( .A1(n_31), .A2(n_83), .B1(n_259), .B2(n_326), .C1(n_338), .C2(n_539), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_32), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_33), .A2(n_183), .B1(n_338), .B2(n_683), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_34), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_35), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_36), .A2(n_48), .B1(n_671), .B2(n_672), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_37), .A2(n_38), .B1(n_582), .B2(n_584), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_39), .A2(n_215), .B1(n_377), .B2(n_567), .Y(n_664) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_40), .A2(n_79), .B1(n_308), .B2(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g833 ( .A(n_40), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_41), .A2(n_127), .B1(n_730), .B2(n_731), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_42), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_43), .A2(n_69), .B1(n_473), .B2(n_549), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_44), .A2(n_46), .B1(n_653), .B2(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_45), .A2(n_111), .B1(n_511), .B2(n_706), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g842 ( .A1(n_47), .A2(n_271), .B1(n_425), .B2(n_698), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_49), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g384 ( .A(n_50), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_51), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_52), .A2(n_84), .B1(n_411), .B2(n_413), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_53), .A2(n_238), .B1(n_408), .B2(n_453), .Y(n_659) );
AOI22xp5_ASAP7_75t_SL g665 ( .A1(n_54), .A2(n_266), .B1(n_666), .B2(n_668), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_56), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_57), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_58), .A2(n_203), .B1(n_402), .B2(n_452), .Y(n_849) );
AOI222xp33_ASAP7_75t_L g876 ( .A1(n_59), .A2(n_192), .B1(n_258), .B2(n_601), .C1(n_698), .C2(n_750), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_60), .A2(n_262), .B1(n_425), .B2(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_61), .B(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_62), .A2(n_237), .B1(n_652), .B2(n_674), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_63), .A2(n_261), .B1(n_640), .B2(n_648), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_64), .A2(n_270), .B1(n_338), .B2(n_478), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_65), .B(n_537), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_66), .A2(n_214), .B1(n_362), .B2(n_412), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_67), .A2(n_182), .B1(n_408), .B2(n_655), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_68), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_71), .A2(n_184), .B1(n_355), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_73), .A2(n_153), .B1(n_371), .B2(n_375), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_74), .A2(n_145), .B1(n_432), .B2(n_468), .Y(n_579) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_75), .A2(n_118), .B1(n_539), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_76), .A2(n_273), .B1(n_457), .B2(n_462), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_78), .A2(n_140), .B1(n_362), .B2(n_365), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_80), .A2(n_268), .B1(n_450), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_81), .A2(n_220), .B1(n_401), .B2(n_507), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_82), .A2(n_212), .B1(n_448), .B2(n_674), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_86), .Y(n_864) );
INVx1_ASAP7_75t_L g294 ( .A(n_87), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_88), .B(n_643), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_89), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_90), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_91), .B(n_495), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_92), .A2(n_186), .B1(n_397), .B2(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g290 ( .A(n_93), .Y(n_290) );
INVx1_ASAP7_75t_L g684 ( .A(n_94), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_95), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_96), .A2(n_207), .B1(n_413), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_97), .A2(n_142), .B1(n_375), .B2(n_507), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_98), .A2(n_240), .B1(n_365), .B2(n_567), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_99), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_100), .A2(n_170), .B1(n_373), .B2(n_412), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_101), .A2(n_193), .B1(n_617), .B2(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_102), .A2(n_113), .B1(n_397), .B2(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_103), .A2(n_157), .B1(n_539), .B2(n_648), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_104), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_105), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_106), .Y(n_302) );
INVx1_ASAP7_75t_L g550 ( .A(n_107), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_108), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_109), .A2(n_161), .B1(n_332), .B2(n_338), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_110), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_112), .A2(n_126), .B1(n_379), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_114), .A2(n_123), .B1(n_332), .B2(n_564), .Y(n_804) );
INVx1_ASAP7_75t_L g542 ( .A(n_115), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_116), .A2(n_225), .B1(n_413), .B2(n_766), .Y(n_765) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_117), .A2(n_741), .B1(n_742), .B2(n_768), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_117), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_119), .A2(n_255), .B1(n_411), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_120), .B(n_496), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_122), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_124), .A2(n_276), .B1(n_507), .B2(n_593), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_125), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_128), .A2(n_130), .B1(n_355), .B2(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g545 ( .A(n_129), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_131), .A2(n_202), .B1(n_362), .B2(n_365), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_132), .A2(n_167), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_133), .A2(n_181), .B1(n_188), .B2(n_327), .C1(n_332), .C2(n_496), .Y(n_552) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_134), .A2(n_169), .B1(n_216), .B2(n_327), .C1(n_478), .C2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_135), .A2(n_254), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_136), .A2(n_198), .B1(n_624), .B2(n_655), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_137), .A2(n_243), .B1(n_400), .B2(n_668), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_138), .A2(n_201), .B1(n_624), .B2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_139), .A2(n_281), .B1(n_456), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_141), .A2(n_260), .B1(n_528), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_143), .Y(n_426) );
AND2x2_ASAP7_75t_L g293 ( .A(n_144), .B(n_294), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_146), .A2(n_211), .B1(n_530), .B2(n_619), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_147), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_149), .A2(n_245), .B1(n_432), .B2(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_150), .Y(n_752) );
AOI222xp33_ASAP7_75t_L g795 ( .A1(n_151), .A2(n_162), .B1(n_226), .B2(n_327), .C1(n_683), .C2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_154), .A2(n_246), .B1(n_464), .B2(n_468), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_155), .A2(n_229), .B1(n_476), .B2(n_530), .Y(n_658) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_156), .A2(n_284), .B1(n_452), .B2(n_708), .Y(n_707) );
AND2x6_ASAP7_75t_L g289 ( .A(n_158), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_158), .Y(n_826) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_159), .A2(n_236), .B1(n_308), .B2(n_312), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_160), .A2(n_269), .B1(n_453), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_163), .A2(n_204), .B1(n_476), .B2(n_549), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_164), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_165), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_166), .A2(n_235), .B1(n_379), .B2(n_381), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_168), .Y(n_498) );
INVx1_ASAP7_75t_L g594 ( .A(n_172), .Y(n_594) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_173), .B(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_174), .A2(n_176), .B1(n_613), .B2(n_615), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_177), .A2(n_275), .B1(n_472), .B2(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g533 ( .A(n_178), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_179), .A2(n_688), .B1(n_689), .B2(n_712), .Y(n_687) );
CKINVDCx14_ASAP7_75t_R g712 ( .A(n_179), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_180), .Y(n_435) );
INVx1_ASAP7_75t_L g553 ( .A(n_185), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_187), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_189), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_190), .A2(n_233), .B1(n_511), .B2(n_560), .Y(n_589) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_191), .A2(n_247), .B1(n_308), .B2(n_309), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g725 ( .A1(n_195), .A2(n_251), .B1(n_381), .B2(n_472), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_196), .B(n_460), .Y(n_844) );
XOR2x2_ASAP7_75t_L g444 ( .A(n_197), .B(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g726 ( .A1(n_199), .A2(n_206), .B1(n_362), .B2(n_560), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_200), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_208), .A2(n_256), .B1(n_464), .B2(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g346 ( .A(n_209), .Y(n_346) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_210), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_213), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_217), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_218), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_219), .A2(n_481), .B1(n_514), .B2(n_515), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_219), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_221), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_223), .B(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g585 ( .A1(n_224), .A2(n_279), .B1(n_466), .B2(n_478), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_227), .A2(n_274), .B1(n_415), .B2(n_854), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_228), .A2(n_253), .B1(n_362), .B2(n_365), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_230), .A2(n_836), .B1(n_837), .B2(n_855), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_230), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_231), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_234), .A2(n_278), .B1(n_400), .B2(n_402), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_236), .B(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_241), .A2(n_257), .B1(n_582), .B2(n_584), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_242), .A2(n_250), .B1(n_475), .B2(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g829 ( .A(n_247), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_248), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_249), .A2(n_280), .B1(n_456), .B2(n_460), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_252), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_263), .A2(n_265), .B1(n_373), .B2(n_375), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_264), .Y(n_841) );
INVx1_ASAP7_75t_L g308 ( .A(n_267), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_272), .A2(n_287), .B(n_295), .C(n_834), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_277), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_282), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_283), .B(n_457), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_285), .A2(n_771), .B1(n_797), .B2(n_798), .Y(n_770) );
CKINVDCx16_ASAP7_75t_R g797 ( .A(n_285), .Y(n_797) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
HB1xp67_ASAP7_75t_L g825 ( .A(n_290), .Y(n_825) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_291), .A2(n_824), .B(n_863), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_629), .B1(n_819), .B2(n_820), .C(n_821), .Y(n_295) );
INVx1_ASAP7_75t_L g819 ( .A(n_296), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_521), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_385), .B1(n_519), .B2(n_520), .Y(n_297) );
INVx2_ASAP7_75t_SL g519 ( .A(n_298), .Y(n_519) );
XOR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_384), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_352), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_323), .C(n_341), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_318), .B2(n_319), .Y(n_301) );
BUFx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g420 ( .A(n_304), .Y(n_420) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_304), .Y(n_791) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_313), .Y(n_304) );
INVx2_ASAP7_75t_L g374 ( .A(n_305), .Y(n_374) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_311), .Y(n_305) );
AND2x2_ASAP7_75t_L g322 ( .A(n_306), .B(n_311), .Y(n_322) );
AND2x2_ASAP7_75t_L g357 ( .A(n_306), .B(n_336), .Y(n_357) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g328 ( .A(n_307), .B(n_311), .Y(n_328) );
AND2x2_ASAP7_75t_L g337 ( .A(n_307), .B(n_317), .Y(n_337) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_310), .Y(n_312) );
INVx2_ASAP7_75t_L g336 ( .A(n_311), .Y(n_336) );
INVx1_ASAP7_75t_L g367 ( .A(n_311), .Y(n_367) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_314), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g380 ( .A(n_314), .B(n_357), .Y(n_380) );
AND2x4_ASAP7_75t_L g459 ( .A(n_314), .B(n_374), .Y(n_459) );
AND2x6_ASAP7_75t_L g462 ( .A(n_314), .B(n_322), .Y(n_462) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g330 ( .A(n_315), .Y(n_330) );
INVx1_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_315), .B(n_317), .Y(n_368) );
AND2x2_ASAP7_75t_L g329 ( .A(n_316), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g360 ( .A(n_317), .B(n_351), .Y(n_360) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g422 ( .A(n_320), .Y(n_422) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g488 ( .A(n_321), .Y(n_488) );
AND2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_360), .Y(n_364) );
AND2x4_ASAP7_75t_L g377 ( .A(n_322), .B(n_329), .Y(n_377) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B(n_331), .Y(n_323) );
OAI21xp5_ASAP7_75t_SL g716 ( .A1(n_325), .A2(n_717), .B(n_718), .Y(n_716) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_327), .Y(n_428) );
INVx2_ASAP7_75t_L g577 ( .A(n_327), .Y(n_577) );
INVx2_ASAP7_75t_SL g635 ( .A(n_327), .Y(n_635) );
INVx4_ASAP7_75t_L g680 ( .A(n_327), .Y(n_680) );
AND2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g348 ( .A(n_328), .Y(n_348) );
AND2x4_ASAP7_75t_L g469 ( .A(n_328), .B(n_350), .Y(n_469) );
AND2x2_ASAP7_75t_L g356 ( .A(n_329), .B(n_357), .Y(n_356) );
AND2x6_ASAP7_75t_L g373 ( .A(n_329), .B(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_332), .Y(n_425) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx4f_ASAP7_75t_SL g478 ( .A(n_333), .Y(n_478) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_333), .Y(n_601) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_333), .Y(n_647) );
BUFx2_ASAP7_75t_L g683 ( .A(n_333), .Y(n_683) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g340 ( .A(n_335), .Y(n_340) );
INVx1_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
AND2x4_ASAP7_75t_L g339 ( .A(n_337), .B(n_340), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_337), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g466 ( .A(n_337), .B(n_467), .Y(n_466) );
BUFx4f_ASAP7_75t_SL g479 ( .A(n_338), .Y(n_479) );
INVx2_ASAP7_75t_L g699 ( .A(n_338), .Y(n_699) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_339), .Y(n_432) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_339), .Y(n_496) );
INVx1_ASAP7_75t_L g603 ( .A(n_339), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_346), .B2(n_347), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_343), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
BUFx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx4_ASAP7_75t_L g437 ( .A(n_344), .Y(n_437) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_344), .Y(n_499) );
AND2x2_ASAP7_75t_L g560 ( .A(n_345), .B(n_383), .Y(n_560) );
CKINVDCx16_ASAP7_75t_R g440 ( .A(n_347), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_347), .A2(n_499), .B1(n_701), .B2(n_702), .Y(n_700) );
OR2x6_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_369), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_361), .Y(n_353) );
BUFx2_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_356), .Y(n_412) );
INVx2_ASAP7_75t_L g656 ( .A(n_356), .Y(n_656) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_356), .Y(n_706) );
AND2x2_ASAP7_75t_L g359 ( .A(n_357), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g382 ( .A(n_357), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_357), .B(n_360), .Y(n_394) );
BUFx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx3_ASAP7_75t_L g472 ( .A(n_359), .Y(n_472) );
BUFx3_ASAP7_75t_L g567 ( .A(n_359), .Y(n_567) );
BUFx3_ASAP7_75t_L g653 ( .A(n_359), .Y(n_653) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx5_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
BUFx3_ASAP7_75t_L g531 ( .A(n_363), .Y(n_531) );
INVx4_ASAP7_75t_L g667 ( .A(n_363), .Y(n_667) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
BUFx2_ASAP7_75t_L g453 ( .A(n_365), .Y(n_453) );
BUFx2_ASAP7_75t_L g668 ( .A(n_365), .Y(n_668) );
BUFx2_ASAP7_75t_L g708 ( .A(n_365), .Y(n_708) );
INVx6_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g619 ( .A(n_366), .Y(n_619) );
OR2x6_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g467 ( .A(n_367), .Y(n_467) );
INVx1_ASAP7_75t_L g383 ( .A(n_368), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_378), .Y(n_369) );
INVx1_ASAP7_75t_SL g404 ( .A(n_371), .Y(n_404) );
INVx4_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g475 ( .A(n_372), .Y(n_475) );
INVx2_ASAP7_75t_SL g617 ( .A(n_372), .Y(n_617) );
INVx2_ASAP7_75t_L g672 ( .A(n_372), .Y(n_672) );
INVx5_ASAP7_75t_SL g787 ( .A(n_372), .Y(n_787) );
INVx11_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx11_ASAP7_75t_L g508 ( .A(n_373), .Y(n_508) );
INVx1_ASAP7_75t_L g551 ( .A(n_375), .Y(n_551) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g476 ( .A(n_376), .Y(n_476) );
INVx2_ASAP7_75t_L g776 ( .A(n_376), .Y(n_776) );
INVx6_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
BUFx3_ASAP7_75t_L g593 ( .A(n_377), .Y(n_593) );
INVxp67_ASAP7_75t_L g782 ( .A(n_379), .Y(n_782) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
INVx2_ASAP7_75t_L g512 ( .A(n_380), .Y(n_512) );
BUFx3_ASAP7_75t_L g731 ( .A(n_380), .Y(n_731) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g397 ( .A(n_382), .Y(n_397) );
BUFx3_ASAP7_75t_L g473 ( .A(n_382), .Y(n_473) );
BUFx3_ASAP7_75t_L g624 ( .A(n_382), .Y(n_624) );
BUFx2_ASAP7_75t_SL g674 ( .A(n_382), .Y(n_674) );
INVx1_ASAP7_75t_L g809 ( .A(n_382), .Y(n_809) );
BUFx2_ASAP7_75t_SL g852 ( .A(n_382), .Y(n_852) );
INVx1_ASAP7_75t_L g520 ( .A(n_385), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_443), .B2(n_518), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_416), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_403), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_395), .B1(n_396), .B2(n_398), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g543 ( .A(n_393), .Y(n_543) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_401), .Y(n_452) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B1(n_406), .B2(n_409), .C(n_410), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g614 ( .A(n_412), .Y(n_614) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_412), .Y(n_671) );
BUFx3_ASAP7_75t_L g764 ( .A(n_412), .Y(n_764) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_423), .C(n_434), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_421), .B2(n_422), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_419), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g693 ( .A(n_420), .Y(n_693) );
INVx1_ASAP7_75t_SL g746 ( .A(n_420), .Y(n_746) );
OAI222xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_429), .C1(n_430), .C2(n_433), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g748 ( .A1(n_424), .A2(n_749), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_748) );
INVx2_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_SL g490 ( .A(n_428), .Y(n_490) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g796 ( .A(n_432), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_438), .B2(n_439), .Y(n_434) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_439), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_497) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g757 ( .A(n_440), .Y(n_757) );
INVx3_ASAP7_75t_L g518 ( .A(n_443), .Y(n_518) );
OA22x2_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_480), .B1(n_516), .B2(n_517), .Y(n_443) );
INVx1_ASAP7_75t_L g517 ( .A(n_444), .Y(n_517) );
NAND4xp75_ASAP7_75t_L g445 ( .A(n_446), .B(n_454), .C(n_470), .D(n_477), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .Y(n_446) );
INVx4_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx3_ASAP7_75t_L g528 ( .A(n_449), .Y(n_528) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_SL g454 ( .A(n_455), .B(n_463), .Y(n_454) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_457), .Y(n_643) );
INVx5_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g537 ( .A(n_458), .Y(n_537) );
INVx2_ASAP7_75t_L g582 ( .A(n_458), .Y(n_582) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g609 ( .A(n_461), .Y(n_609) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_462), .Y(n_584) );
BUFx2_ASAP7_75t_L g645 ( .A(n_462), .Y(n_645) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g564 ( .A(n_466), .Y(n_564) );
BUFx2_ASAP7_75t_L g607 ( .A(n_466), .Y(n_607) );
BUFx2_ASAP7_75t_L g648 ( .A(n_466), .Y(n_648) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_469), .Y(n_640) );
BUFx2_ASAP7_75t_SL g814 ( .A(n_469), .Y(n_814) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g505 ( .A(n_472), .Y(n_505) );
BUFx2_ASAP7_75t_L g622 ( .A(n_472), .Y(n_622) );
INVxp67_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
INVx1_ASAP7_75t_L g492 ( .A(n_478), .Y(n_492) );
INVx1_ASAP7_75t_L g516 ( .A(n_480), .Y(n_516) );
INVx2_ASAP7_75t_L g515 ( .A(n_481), .Y(n_515) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_501), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_489), .C(n_497), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_486), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
OAI221xp5_ASAP7_75t_SL g790 ( .A1(n_486), .A2(n_791), .B1(n_792), .B2(n_793), .C(n_794), .Y(n_790) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx3_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B1(n_492), .B2(n_493), .C(n_494), .Y(n_489) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_490), .A2(n_599), .B1(n_600), .B2(n_602), .C1(n_603), .C2(n_604), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g840 ( .A1(n_490), .A2(n_841), .B(n_842), .Y(n_840) );
BUFx4f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g549 ( .A(n_508), .Y(n_549) );
INVx2_ASAP7_75t_SL g854 ( .A(n_508), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_554), .B2(n_628), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
XOR2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_553), .Y(n_524) );
NAND4xp75_ASAP7_75t_L g525 ( .A(n_526), .B(n_532), .C(n_540), .D(n_552), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OA211x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .C(n_538), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_534), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_691) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_546), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_543), .A2(n_774), .B1(n_775), .B2(n_777), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_550), .B2(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g628 ( .A(n_554), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_571), .B1(n_626), .B2(n_627), .Y(n_554) );
INVx2_ASAP7_75t_SL g626 ( .A(n_555), .Y(n_626) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_570), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g556 ( .A(n_557), .B(n_561), .C(n_565), .D(n_569), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g767 ( .A(n_567), .Y(n_767) );
INVx2_ASAP7_75t_L g627 ( .A(n_571), .Y(n_627) );
OA22x2_ASAP7_75t_SL g571 ( .A1(n_572), .A2(n_573), .B1(n_595), .B2(n_625), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
XOR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_594), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_575), .B(n_586), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
OAI21xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_578), .B(n_579), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .C(n_585), .Y(n_580) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g625 ( .A(n_595), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_610), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_605), .Y(n_597) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_620), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_618), .Y(n_611) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g820 ( .A(n_629), .Y(n_820) );
AOI22xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_738), .B1(n_817), .B2(n_818), .Y(n_629) );
INVx1_ASAP7_75t_L g817 ( .A(n_630), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_660), .B1(n_736), .B2(n_737), .Y(n_630) );
INVx2_ASAP7_75t_L g736 ( .A(n_631), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_633), .B(n_649), .Y(n_632) );
NOR2xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_641), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_636), .B(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .C(n_646), .Y(n_641) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_657), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
BUFx4f_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g730 ( .A(n_656), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g737 ( .A(n_660), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_685), .B1(n_686), .B2(n_735), .Y(n_660) );
INVx2_ASAP7_75t_SL g735 ( .A(n_661), .Y(n_735) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_684), .Y(n_661) );
NOR4xp75_ASAP7_75t_L g662 ( .A(n_663), .B(n_669), .C(n_675), .D(n_678), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_665), .Y(n_663) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_SL g780 ( .A(n_671), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_676), .B(n_677), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_681), .B(n_682), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_679), .A2(n_696), .B(n_697), .Y(n_695) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx4_ASAP7_75t_L g750 ( .A(n_680), .Y(n_750) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
AO22x1_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_713), .B1(n_733), .B2(n_734), .Y(n_686) );
INVx1_ASAP7_75t_L g734 ( .A(n_687), .Y(n_734) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_703), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_695), .C(n_700), .Y(n_690) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_709), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx3_ASAP7_75t_SL g733 ( .A(n_713), .Y(n_733) );
XOR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_732), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_723), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .C(n_722), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g818 ( .A(n_738), .Y(n_818) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_769), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_758), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .C(n_754), .Y(n_743) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_765), .Y(n_762) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_799), .B1(n_815), .B2(n_816), .Y(n_769) );
INVx1_ASAP7_75t_L g815 ( .A(n_770), .Y(n_815) );
INVx2_ASAP7_75t_SL g798 ( .A(n_771), .Y(n_798) );
AND4x1_ASAP7_75t_L g771 ( .A(n_772), .B(n_783), .C(n_789), .D(n_795), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_778), .Y(n_772) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B1(n_781), .B2(n_782), .Y(n_778) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_788), .Y(n_783) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_L g816 ( .A(n_799), .Y(n_816) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .C(n_810), .D(n_813), .Y(n_801) );
AND2x2_ASAP7_75t_SL g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_SL g821 ( .A(n_822), .Y(n_821) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_827), .Y(n_822) );
OR2x2_ASAP7_75t_SL g879 ( .A(n_823), .B(n_828), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_826), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_825), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_825), .B(n_860), .Y(n_863) );
CKINVDCx16_ASAP7_75t_R g860 ( .A(n_826), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
OAI322xp33_ASAP7_75t_L g834 ( .A1(n_835), .A2(n_856), .A3(n_857), .B1(n_861), .B2(n_864), .C1(n_865), .C2(n_877), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_837), .Y(n_836) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_847), .C(n_850), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .C(n_846), .Y(n_843) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_853), .Y(n_850) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
HB1xp67_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
CKINVDCx16_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
XOR2x2_ASAP7_75t_L g865 ( .A(n_864), .B(n_866), .Y(n_865) );
NAND4xp75_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .C(n_873), .D(n_876), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
AND2x2_ASAP7_75t_SL g870 ( .A(n_871), .B(n_872), .Y(n_870) );
AND2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_879), .Y(n_878) );
endmodule