module fake_jpeg_29764_n_410 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_410);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_47),
.B(n_50),
.Y(n_134)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_14),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_61),
.Y(n_101)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_71),
.Y(n_104)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_69),
.Y(n_96)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_18),
.B(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_22),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_81),
.Y(n_116)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_25),
.Y(n_113)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_1),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_33),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_113),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_39),
.B1(n_41),
.B2(n_30),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_124),
.B(n_64),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_100),
.B(n_120),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_56),
.B1(n_30),
.B2(n_34),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_119),
.B1(n_125),
.B2(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_42),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_42),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_44),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_71),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_40),
.B(n_38),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_32),
.B1(n_40),
.B2(n_43),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_16),
.B1(n_35),
.B2(n_33),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_11),
.B1(n_12),
.B2(n_129),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_45),
.A2(n_32),
.B1(n_43),
.B2(n_35),
.Y(n_129)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_84),
.B1(n_83),
.B2(n_49),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_137),
.A2(n_159),
.B1(n_164),
.B2(n_93),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_138),
.B(n_163),
.Y(n_203)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_103),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_86),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_68),
.B1(n_81),
.B2(n_78),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_153),
.B1(n_155),
.B2(n_168),
.Y(n_216)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_22),
.B(n_38),
.C(n_58),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_119),
.B(n_128),
.C(n_95),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_148),
.B(n_166),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_149),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_73),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_59),
.B1(n_75),
.B2(n_63),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_3),
.B(n_4),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_132),
.B(n_95),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_52),
.B1(n_82),
.B2(n_51),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_106),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_174),
.B1(n_180),
.B2(n_112),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_109),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_111),
.A2(n_132),
.B1(n_127),
.B2(n_112),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_167),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_6),
.B1(n_8),
.B2(n_11),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_176),
.Y(n_182)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_175),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_11),
.C(n_12),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_123),
.C(n_128),
.Y(n_195)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_102),
.A2(n_11),
.B1(n_12),
.B2(n_122),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_179),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_121),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_203),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_186),
.A2(n_193),
.B(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_200),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_180),
.B1(n_149),
.B2(n_127),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_201),
.B1(n_209),
.B2(n_148),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_136),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_205),
.B1(n_212),
.B2(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_123),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_110),
.B1(n_122),
.B2(n_88),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_110),
.B1(n_94),
.B2(n_105),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_202),
.B(n_158),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_93),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_213),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_105),
.B1(n_178),
.B2(n_151),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_163),
.A2(n_146),
.B1(n_142),
.B2(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_142),
.B(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_197),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_140),
.A2(n_143),
.B1(n_158),
.B2(n_152),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_222),
.A2(n_230),
.B(n_217),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_183),
.Y(n_225)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_185),
.A2(n_187),
.B(n_200),
.C(n_204),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_250),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_233),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_172),
.B(n_139),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_207),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_237),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_170),
.B1(n_156),
.B2(n_173),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_238),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_169),
.B1(n_145),
.B2(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_245),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_139),
.B1(n_202),
.B2(n_216),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_240),
.A2(n_241),
.B1(n_181),
.B2(n_228),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_194),
.B1(n_212),
.B2(n_202),
.Y(n_241)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_206),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_249),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_196),
.B(n_192),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_185),
.B1(n_184),
.B2(n_186),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_248),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_182),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_195),
.B(n_182),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_210),
.C(n_182),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_217),
.C(n_192),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_191),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_247),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_190),
.B(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_235),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_211),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_257),
.A2(n_269),
.B(n_279),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_265),
.B(n_237),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_267),
.Y(n_292)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_263),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_196),
.B(n_191),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_268),
.B(n_230),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_252),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_271),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_242),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_243),
.C(n_279),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_222),
.A2(n_181),
.B(n_251),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_286),
.B1(n_232),
.B2(n_233),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_271),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_285),
.Y(n_287)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_250),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_297),
.C(n_300),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_221),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_228),
.B1(n_241),
.B2(n_234),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_281),
.B1(n_270),
.B2(n_267),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_223),
.B(n_224),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_305),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_221),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_298),
.B(n_299),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_236),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_225),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_262),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_283),
.B(n_226),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_303),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_227),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_262),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_277),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_257),
.A2(n_255),
.B1(n_243),
.B2(n_229),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_272),
.B1(n_265),
.B2(n_256),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_260),
.C(n_275),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_310),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_313),
.A2(n_306),
.B1(n_272),
.B2(n_288),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_335),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_276),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_302),
.Y(n_349)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_325),
.Y(n_350)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

XOR2x1_ASAP7_75t_SL g327 ( 
.A(n_289),
.B(n_257),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_332),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_277),
.Y(n_329)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_329),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_291),
.A2(n_275),
.B(n_256),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_295),
.B(n_299),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_296),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_333),
.B(n_334),
.C(n_297),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_282),
.C(n_261),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_327),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_341),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_337),
.A2(n_325),
.B1(n_295),
.B2(n_321),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_319),
.A2(n_309),
.B(n_305),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_339),
.A2(n_314),
.B(n_330),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_320),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_344),
.C(n_345),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_347),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_303),
.C(n_300),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_298),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_352),
.C(n_316),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_305),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_348),
.A2(n_328),
.B(n_317),
.Y(n_362)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_316),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_310),
.C(n_273),
.Y(n_352)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_343),
.Y(n_356)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_357),
.A2(n_368),
.B(n_348),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_347),
.A2(n_313),
.B1(n_335),
.B2(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_360),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_325),
.B1(n_319),
.B2(n_326),
.Y(n_361)
);

OAI321xp33_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_366),
.A3(n_341),
.B1(n_338),
.B2(n_337),
.C(n_307),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_364),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_322),
.C(n_328),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_340),
.C(n_345),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_315),
.B1(n_280),
.B2(n_266),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_353),
.A2(n_315),
.B(n_307),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_342),
.B(n_264),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_369),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_356),
.A2(n_350),
.B1(n_336),
.B2(n_354),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_363),
.B(n_338),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_350),
.B(n_336),
.Y(n_372)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_355),
.C(n_360),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_377),
.A2(n_358),
.B1(n_367),
.B2(n_362),
.Y(n_385)
);

NOR2x1_ASAP7_75t_SL g378 ( 
.A(n_368),
.B(n_352),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_372),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_355),
.C(n_365),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_381),
.B(n_382),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_364),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_385),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_374),
.Y(n_392)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_346),
.C(n_357),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_379),
.B(n_363),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_370),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_391),
.B(n_392),
.Y(n_401)
);

AOI322xp5_ASAP7_75t_L g395 ( 
.A1(n_384),
.A2(n_388),
.A3(n_380),
.B1(n_374),
.B2(n_284),
.C1(n_273),
.C2(n_266),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_349),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_391),
.C(n_396),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_381),
.C(n_384),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_400),
.B(n_402),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_373),
.C(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_284),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_404),
.B(n_266),
.C(n_322),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_392),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_401),
.B(n_273),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_407),
.B(n_403),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_263),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_263),
.Y(n_410)
);


endmodule