module fake_jpeg_24304_n_31 (n_3, n_2, n_1, n_0, n_4, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_2),
.Y(n_5)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_10),
.B(n_11),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_5),
.B1(n_7),
.B2(n_6),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_5),
.C(n_7),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_10),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_12),
.B1(n_2),
.B2(n_1),
.Y(n_21)
);

AO22x1_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_11),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_1),
.C(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_15),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_15),
.B(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_20),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI321xp33_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_1),
.A3(n_16),
.B1(n_18),
.B2(n_27),
.C(n_28),
.Y(n_31)
);


endmodule