module fake_jpeg_3258_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_83),
.Y(n_94)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_1),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.B(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_57),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_91),
.B(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_69),
.B1(n_66),
.B2(n_56),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_98),
.B1(n_57),
.B2(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_66),
.B1(n_55),
.B2(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_82),
.B1(n_79),
.B2(n_74),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_101),
.B1(n_71),
.B2(n_59),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_82),
.B1(n_74),
.B2(n_72),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_56),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_65),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_96),
.B1(n_86),
.B2(n_73),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_84),
.B(n_58),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_104),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_117),
.A2(n_102),
.B1(n_113),
.B2(n_108),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_129),
.B(n_71),
.C(n_21),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_125),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_58),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_64),
.C(n_61),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_10),
.C(n_11),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_58),
.B1(n_63),
.B2(n_59),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_71),
.A3(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_2),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_138),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_3),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_6),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_119),
.B1(n_30),
.B2(n_37),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_7),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_8),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_158),
.B1(n_120),
.B2(n_129),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_24),
.B1(n_50),
.B2(n_49),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_12),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_155),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_22),
.B1(n_46),
.B2(n_44),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_12),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_13),
.B(n_14),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_16),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_14),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_166),
.B1(n_171),
.B2(n_176),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_119),
.C(n_29),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_153),
.Y(n_185)
);

INVxp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_180),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_20),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_28),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_157),
.B1(n_148),
.B2(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_189),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_16),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_145),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_199),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_169),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_165),
.B(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_203),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_193),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_200),
.B(n_195),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_192),
.B(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_174),
.C(n_145),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_206),
.A2(n_207),
.B1(n_178),
.B2(n_39),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_208),
.A2(n_201),
.B(n_164),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_210),
.B(n_19),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_42),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_43),
.B(n_51),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_17),
.Y(n_214)
);


endmodule