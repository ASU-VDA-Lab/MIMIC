module fake_jpeg_3493_n_636 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_636);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_636;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_0),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_61),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_64),
.Y(n_144)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_72),
.Y(n_164)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_73),
.Y(n_179)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_76),
.B(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_78),
.Y(n_175)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_84),
.B(n_86),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_91),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_92),
.Y(n_178)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_94),
.Y(n_212)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_95),
.Y(n_213)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_32),
.B(n_0),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_98),
.B(n_105),
.Y(n_183)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_104),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_36),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_114),
.B(n_117),
.Y(n_197)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_45),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_45),
.Y(n_125)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_51),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_128),
.B(n_43),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_65),
.A2(n_20),
.B1(n_56),
.B2(n_53),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_133),
.A2(n_165),
.B1(n_23),
.B2(n_27),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_135),
.B(n_143),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_52),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_138),
.B(n_159),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_124),
.B1(n_72),
.B2(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_140),
.A2(n_158),
.B1(n_207),
.B2(n_218),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_76),
.B(n_20),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_151),
.B(n_173),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_50),
.B1(n_30),
.B2(n_29),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_156),
.B(n_168),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_91),
.A2(n_50),
.B1(n_30),
.B2(n_29),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_64),
.B(n_19),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_75),
.A2(n_19),
.B1(n_56),
.B2(n_53),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_120),
.B(n_52),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_68),
.B(n_57),
.C(n_23),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_174),
.B(n_5),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_21),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_SL g242 ( 
.A(n_187),
.B(n_200),
.C(n_209),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_77),
.B(n_21),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_63),
.Y(n_203)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_107),
.A2(n_30),
.B1(n_50),
.B2(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_78),
.B(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_69),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_79),
.Y(n_214)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_82),
.Y(n_217)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_89),
.A2(n_29),
.B1(n_28),
.B2(n_35),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_85),
.Y(n_219)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_28),
.B1(n_43),
.B2(n_41),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_220),
.A2(n_244),
.B1(n_270),
.B2(n_274),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_226),
.A2(n_261),
.B1(n_178),
.B2(n_212),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_148),
.B(n_130),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_228),
.B(n_233),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_27),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_237),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_232),
.B(n_241),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g233 ( 
.A(n_131),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_211),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_236),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_144),
.A2(n_41),
.B(n_35),
.C(n_2),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_235),
.A2(n_15),
.B(n_212),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_112),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_103),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_176),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_238),
.B(n_258),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_100),
.B(n_94),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_239),
.A2(n_256),
.B(n_290),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_166),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_153),
.A2(n_92),
.B1(n_90),
.B2(n_88),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_166),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_248),
.B(n_252),
.Y(n_328)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_150),
.Y(n_250)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_196),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_251),
.B(n_272),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_168),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_144),
.B(n_87),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_254),
.B(n_281),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_255),
.A2(n_154),
.B1(n_175),
.B2(n_189),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_133),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_164),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_257),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_180),
.B(n_3),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_162),
.Y(n_259)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_156),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_260),
.B(n_145),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_199),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_152),
.Y(n_262)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_279),
.Y(n_338)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_142),
.Y(n_267)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

CKINVDCx12_ASAP7_75t_R g268 ( 
.A(n_157),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_268),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_161),
.A2(n_193),
.B1(n_149),
.B2(n_179),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_179),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_155),
.B(n_15),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_289),
.C(n_175),
.Y(n_341)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_167),
.Y(n_276)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx3_ASAP7_75t_SL g277 ( 
.A(n_196),
.Y(n_277)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_213),
.B(n_7),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_140),
.Y(n_280)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_129),
.B(n_8),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_155),
.Y(n_282)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_147),
.Y(n_283)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_191),
.Y(n_285)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_147),
.Y(n_286)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_134),
.Y(n_287)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_287),
.Y(n_349)
);

HAxp5_ASAP7_75t_SL g288 ( 
.A(n_156),
.B(n_8),
.CON(n_288),
.SN(n_288)
);

OR2x2_ASAP7_75t_SL g350 ( 
.A(n_288),
.B(n_216),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_155),
.B(n_163),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_158),
.A2(n_9),
.B(n_10),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_201),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_296),
.B1(n_171),
.B2(n_139),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_207),
.B(n_141),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_181),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_154),
.Y(n_293)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_177),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_294),
.B(n_295),
.Y(n_342)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_137),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g297 ( 
.A(n_162),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_251),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_242),
.B(n_202),
.CI(n_206),
.CON(n_306),
.SN(n_306)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_306),
.B(n_319),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_307),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_309),
.A2(n_320),
.B1(n_337),
.B2(n_345),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_280),
.A2(n_215),
.B1(n_205),
.B2(n_182),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_316),
.A2(n_318),
.B1(n_323),
.B2(n_257),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_269),
.A2(n_230),
.B1(n_292),
.B2(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_237),
.B(n_141),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_322),
.B(n_336),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_230),
.A2(n_162),
.B1(n_190),
.B2(n_184),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_331),
.B(n_350),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_254),
.B(n_145),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_332),
.B(n_294),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_231),
.B(n_146),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_333),
.B(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_230),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_226),
.A2(n_146),
.B1(n_198),
.B2(n_181),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_341),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_198),
.B1(n_189),
.B2(n_190),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_229),
.B(n_184),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_246),
.B(n_216),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_303),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_239),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_353),
.B(n_297),
.Y(n_392)
);

NAND2x1_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_277),
.Y(n_373)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_345),
.A2(n_288),
.B1(n_272),
.B2(n_256),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_379),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_221),
.B(n_235),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_358),
.A2(n_373),
.B(n_377),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_324),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_359),
.B(n_361),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_353),
.A2(n_224),
.B1(n_261),
.B2(n_275),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_360),
.A2(n_363),
.B1(n_368),
.B2(n_380),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_306),
.B(n_289),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_320),
.A2(n_275),
.B1(n_283),
.B2(n_286),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_324),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_366),
.B(n_375),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_336),
.A2(n_240),
.B1(n_249),
.B2(n_247),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_327),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_372),
.B(n_314),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_355),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_334),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_L g427 ( 
.A1(n_376),
.A2(n_378),
.B(n_392),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_282),
.B(n_257),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_298),
.A2(n_263),
.B(n_262),
.C(n_250),
.Y(n_378)
);

AO22x1_ASAP7_75t_SL g379 ( 
.A1(n_312),
.A2(n_240),
.B1(n_249),
.B2(n_247),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_302),
.A2(n_222),
.B1(n_293),
.B2(n_267),
.Y(n_380)
);

OA22x2_ASAP7_75t_L g381 ( 
.A1(n_339),
.A2(n_266),
.B1(n_295),
.B2(n_287),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_322),
.A2(n_227),
.B1(n_253),
.B2(n_243),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_383),
.A2(n_369),
.B1(n_382),
.B2(n_387),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_312),
.A2(n_266),
.B(n_259),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

INVx13_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_385),
.Y(n_440)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_300),
.A2(n_285),
.B(n_278),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_332),
.A2(n_243),
.B1(n_273),
.B2(n_225),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_399),
.B1(n_401),
.B2(n_356),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_305),
.B(n_223),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_396),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_342),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_394),
.B(n_310),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_313),
.A2(n_328),
.B1(n_350),
.B2(n_325),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_398),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_302),
.B(n_298),
.Y(n_396)
);

NAND2x1p5_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_245),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_341),
.A2(n_265),
.B1(n_271),
.B2(n_313),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_338),
.A2(n_271),
.B1(n_306),
.B2(n_346),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_414),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_363),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_364),
.A2(n_326),
.B1(n_346),
.B2(n_354),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_412),
.A2(n_430),
.B1(n_357),
.B2(n_386),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_364),
.A2(n_326),
.B1(n_354),
.B2(n_349),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_308),
.C(n_327),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_428),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_420),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_308),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_393),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_422),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_376),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_424),
.B(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_344),
.C(n_314),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_344),
.C(n_299),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_398),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_369),
.A2(n_391),
.B1(n_360),
.B2(n_401),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_391),
.A2(n_343),
.B1(n_301),
.B2(n_317),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_436),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_365),
.A2(n_317),
.B1(n_315),
.B2(n_311),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_384),
.B1(n_388),
.B2(n_373),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_373),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_375),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_299),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_439),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_441),
.Y(n_485)
);

INVx4_ASAP7_75t_SL g444 ( 
.A(n_440),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_444),
.B(n_456),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_420),
.B(n_397),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_445),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_377),
.B(n_391),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_446),
.B(n_453),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_437),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_473),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_417),
.C(n_418),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_397),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_451),
.B(n_454),
.Y(n_476)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_419),
.A2(n_370),
.B(n_392),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_383),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_455),
.A2(n_470),
.B1(n_432),
.B2(n_361),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_436),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_425),
.Y(n_459)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_460),
.Y(n_488)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_461),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_368),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_462),
.B(n_468),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_413),
.A2(n_358),
.B(n_395),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_464),
.B(n_413),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_390),
.Y(n_465)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_465),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_410),
.B(n_378),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_467),
.B(n_472),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_428),
.B(n_370),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_366),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_469),
.B(n_471),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_359),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_416),
.A2(n_398),
.B(n_399),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_474),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_405),
.B1(n_407),
.B2(n_404),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g479 ( 
.A(n_457),
.Y(n_479)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

NOR3xp33_ASAP7_75t_SL g482 ( 
.A(n_443),
.B(n_423),
.C(n_408),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_482),
.B(n_498),
.Y(n_518)
);

AOI32xp33_ASAP7_75t_L g483 ( 
.A1(n_441),
.A2(n_408),
.A3(n_403),
.B1(n_426),
.B2(n_430),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_483),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_403),
.Y(n_484)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_448),
.C(n_453),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_489),
.A2(n_493),
.B1(n_495),
.B2(n_503),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_471),
.Y(n_492)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_475),
.A2(n_416),
.B1(n_427),
.B2(n_426),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_455),
.A2(n_442),
.B1(n_463),
.B2(n_456),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_496),
.A2(n_453),
.B1(n_455),
.B2(n_463),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_429),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_442),
.A2(n_404),
.B1(n_416),
.B2(n_426),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_450),
.B1(n_461),
.B2(n_411),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_451),
.B(n_412),
.Y(n_503)
);

AO21x1_ASAP7_75t_L g509 ( 
.A1(n_504),
.A2(n_464),
.B(n_446),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_448),
.B(n_380),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_505),
.B(n_493),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_445),
.B(n_411),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_507),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_468),
.B(n_352),
.Y(n_508)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_508),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_511),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_466),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_510),
.B(n_515),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_466),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_449),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_512),
.B(n_516),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_514),
.A2(n_504),
.B1(n_532),
.B2(n_533),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_465),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_474),
.C(n_473),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_529),
.C(n_531),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_362),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_519),
.B(n_433),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_490),
.B(n_444),
.Y(n_521)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_521),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_489),
.A2(n_454),
.B1(n_462),
.B2(n_444),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_522),
.A2(n_530),
.B1(n_492),
.B2(n_500),
.Y(n_549)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_472),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_527),
.B(n_501),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_485),
.B(n_459),
.C(n_458),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_495),
.A2(n_450),
.B1(n_452),
.B2(n_460),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_483),
.B(n_469),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_533),
.A2(n_524),
.B1(n_526),
.B2(n_501),
.Y(n_554)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_478),
.Y(n_535)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_535),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_485),
.B(n_321),
.C(n_433),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_536),
.B(n_440),
.C(n_494),
.Y(n_557)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_537),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_521),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_538),
.B(n_560),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_532),
.A2(n_486),
.B(n_491),
.Y(n_539)
);

OAI21x1_ASAP7_75t_SL g561 ( 
.A1(n_539),
.A2(n_542),
.B(n_551),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_529),
.B(n_491),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_530),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_476),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_SL g573 ( 
.A(n_546),
.B(n_513),
.C(n_534),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_549),
.A2(n_523),
.B1(n_528),
.B2(n_522),
.Y(n_574)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_550),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_514),
.A2(n_486),
.B(n_502),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_553),
.B(n_557),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_554),
.A2(n_503),
.B1(n_499),
.B2(n_517),
.Y(n_578)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_537),
.Y(n_555)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_555),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_531),
.A2(n_486),
.B(n_502),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_556),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_511),
.B(n_494),
.C(n_481),
.Y(n_560)
);

INVx13_ASAP7_75t_L g562 ( 
.A(n_559),
.Y(n_562)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

XNOR2x1_ASAP7_75t_L g580 ( 
.A(n_564),
.B(n_573),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_542),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_566),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_520),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_558),
.C(n_544),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_568),
.B(n_575),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_544),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_571),
.B(n_577),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_574),
.A2(n_499),
.B1(n_476),
.B2(n_527),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_552),
.B(n_516),
.C(n_512),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_548),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_579),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_509),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_578),
.A2(n_556),
.B1(n_549),
.B2(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_581),
.A2(n_591),
.B1(n_592),
.B2(n_593),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_557),
.C(n_540),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_583),
.B(n_585),
.C(n_590),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_540),
.C(n_547),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_545),
.Y(n_587)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_587),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_551),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_589),
.B(n_573),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_536),
.C(n_541),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_518),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_578),
.A2(n_541),
.B1(n_482),
.B2(n_555),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_488),
.C(n_480),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_595),
.B(n_569),
.C(n_567),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_582),
.A2(n_572),
.B1(n_574),
.B2(n_566),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_598),
.B(n_601),
.Y(n_609)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_600),
.Y(n_615)
);

BUFx24_ASAP7_75t_SL g601 ( 
.A(n_594),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_583),
.A2(n_561),
.B(n_585),
.Y(n_602)
);

AOI31xp67_ASAP7_75t_L g613 ( 
.A1(n_602),
.A2(n_604),
.A3(n_607),
.B(n_608),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_570),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_603),
.B(n_606),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_584),
.A2(n_564),
.B(n_562),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_605),
.B(n_580),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_588),
.A2(n_543),
.B1(n_488),
.B2(n_481),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_584),
.A2(n_543),
.B(n_480),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_593),
.A2(n_402),
.B(n_381),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_597),
.A2(n_580),
.B(n_595),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_610),
.A2(n_614),
.B(n_616),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_617),
.Y(n_625)
);

OA21x2_ASAP7_75t_SL g614 ( 
.A1(n_599),
.A2(n_586),
.B(n_589),
.Y(n_614)
);

AOI31xp67_ASAP7_75t_L g616 ( 
.A1(n_596),
.A2(n_357),
.A3(n_379),
.B(n_311),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_605),
.A2(n_330),
.B(n_343),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_597),
.B(n_301),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_618),
.B(n_381),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_600),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_619),
.B(n_622),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g620 ( 
.A1(n_609),
.A2(n_310),
.B1(n_340),
.B2(n_330),
.C(n_357),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_620),
.A2(n_621),
.B1(n_624),
.B2(n_321),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_381),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_381),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_623),
.A2(n_613),
.B(n_616),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_626),
.A2(n_629),
.B1(n_621),
.B2(n_385),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_627),
.Y(n_631)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_625),
.A2(n_385),
.B(n_340),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_630),
.B(n_631),
.C(n_628),
.Y(n_632)
);

BUFx24_ASAP7_75t_SL g633 ( 
.A(n_632),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_633),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_634),
.B(n_379),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_379),
.B(n_352),
.Y(n_636)
);


endmodule