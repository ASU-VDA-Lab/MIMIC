module fake_jpeg_26771_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_51),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_16),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_30),
.B(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_29),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_68),
.Y(n_114)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_43),
.B1(n_44),
.B2(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_100),
.B1(n_29),
.B2(n_32),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_71),
.Y(n_112)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_96),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_50),
.B(n_56),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_36),
.C(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_26),
.B1(n_44),
.B2(n_39),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_91),
.B1(n_21),
.B2(n_22),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_26),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_87),
.Y(n_135)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_44),
.B1(n_39),
.B2(n_36),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_50),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_28),
.B1(n_40),
.B2(n_45),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_45),
.B(n_42),
.C(n_37),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g109 ( 
.A1(n_77),
.A2(n_25),
.B1(n_45),
.B2(n_37),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_124),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_34),
.B(n_22),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_83),
.B1(n_92),
.B2(n_31),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_45),
.C(n_40),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_132),
.B1(n_134),
.B2(n_72),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_80),
.A2(n_45),
.B1(n_42),
.B2(n_37),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_45),
.B1(n_42),
.B2(n_20),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_106),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_137),
.B(n_146),
.C(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_143),
.Y(n_169)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_147),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_144),
.B(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_145),
.B(n_154),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_9),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_67),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_89),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_158),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_123),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_12),
.C(n_15),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_125),
.B1(n_156),
.B2(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_119),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_155),
.B1(n_84),
.B2(n_102),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_93),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_83),
.B1(n_66),
.B2(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_156),
.B(n_161),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_34),
.B(n_31),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_34),
.B(n_30),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_79),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_98),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_160),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_21),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_21),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_164),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_108),
.B1(n_118),
.B2(n_105),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_191),
.B1(n_195),
.B2(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_127),
.B1(n_110),
.B2(n_128),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_175),
.B1(n_155),
.B2(n_154),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_107),
.C(n_110),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_176),
.C(n_188),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_128),
.A3(n_107),
.B1(n_120),
.B2(n_20),
.Y(n_170)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_171),
.B(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_187),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_139),
.A2(n_108),
.B1(n_117),
.B2(n_120),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_90),
.C(n_117),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_28),
.B(n_31),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_180),
.B(n_17),
.Y(n_204)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_27),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_90),
.C(n_112),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_143),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_28),
.Y(n_228)
);

NAND2x1_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_125),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_193),
.A2(n_157),
.B(n_146),
.C(n_147),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_118),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_27),
.C(n_103),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_14),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_169),
.B(n_138),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_207),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_199),
.A2(n_201),
.B1(n_205),
.B2(n_213),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_203),
.B(n_224),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_186),
.B1(n_193),
.B2(n_167),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_219),
.B(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_177),
.A2(n_164),
.B1(n_147),
.B2(n_163),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_169),
.B(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_182),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_151),
.B1(n_141),
.B2(n_112),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_180),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_73),
.C(n_42),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_165),
.C(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_17),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_30),
.B(n_20),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_17),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_222),
.Y(n_251)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_193),
.A2(n_113),
.B1(n_133),
.B2(n_27),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_27),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_227),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_133),
.B(n_28),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_28),
.B(n_133),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_228),
.B(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_195),
.A2(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_196),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_194),
.B1(n_197),
.B2(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_234),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_171),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_214),
.C(n_213),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_242),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_179),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_243),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_170),
.B1(n_168),
.B2(n_190),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_202),
.B1(n_205),
.B2(n_227),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_181),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_181),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_262),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_268),
.C(n_200),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_211),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_230),
.B(n_201),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_226),
.C(n_200),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_237),
.C(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_251),
.B1(n_267),
.B2(n_245),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_199),
.B1(n_253),
.B2(n_248),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_248),
.B1(n_241),
.B2(n_249),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_242),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_282),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_279),
.A2(n_283),
.B1(n_262),
.B2(n_256),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_250),
.B(n_200),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_280),
.A2(n_285),
.B(n_259),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_R g281 ( 
.A(n_270),
.B(n_232),
.C(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_250),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_222),
.B1(n_253),
.B2(n_235),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_200),
.B(n_245),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_239),
.B1(n_234),
.B2(n_251),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_283),
.B1(n_291),
.B2(n_292),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_261),
.B1(n_273),
.B2(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_257),
.B(n_225),
.C(n_219),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_254),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

OAI321xp33_ASAP7_75t_L g310 ( 
.A1(n_296),
.A2(n_298),
.A3(n_307),
.B1(n_293),
.B2(n_302),
.C(n_295),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_0),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_264),
.B(n_263),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_306),
.B1(n_13),
.B2(n_12),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_9),
.B(n_5),
.Y(n_316)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_305),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_260),
.C(n_265),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_275),
.B(n_278),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_SL g305 ( 
.A1(n_285),
.A2(n_265),
.A3(n_256),
.B1(n_204),
.B2(n_225),
.C1(n_258),
.C2(n_272),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_0),
.B(n_3),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_282),
.C(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_277),
.C(n_14),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_13),
.C(n_12),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_296),
.B(n_9),
.CI(n_4),
.CON(n_314),
.SN(n_314)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_318),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_294),
.B1(n_298),
.B2(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_307),
.Y(n_323)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_323),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_0),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_330),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_312),
.B1(n_308),
.B2(n_311),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_322),
.B1(n_320),
.B2(n_7),
.Y(n_333)
);

NAND4xp25_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_321),
.C(n_320),
.D(n_325),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_5),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_331),
.B1(n_334),
.B2(n_329),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_332),
.B(n_6),
.C(n_7),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_5),
.C(n_6),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_6),
.Y(n_341)
);


endmodule