module fake_aes_11211_n_833 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_833);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_833;
wire n_663;
wire n_791;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_818;
wire n_725;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_243;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_409;
wire n_315;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_28), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_214), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_113), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_152), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_51), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_52), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_14), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_125), .B(n_93), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_104), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_60), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_82), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_136), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_118), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_202), .Y(n_252) );
INVx1_ASAP7_75t_SL g253 ( .A(n_138), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_190), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_130), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_227), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_126), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_135), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_32), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_219), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_158), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_66), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_124), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_228), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_64), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_54), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_218), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_44), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_87), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_204), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_123), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_15), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_216), .B(n_115), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_211), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_102), .Y(n_275) );
BUFx5_ASAP7_75t_L g276 ( .A(n_173), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_112), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_231), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_22), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_29), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_75), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_88), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_197), .Y(n_284) );
BUFx10_ASAP7_75t_L g285 ( .A(n_176), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_58), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_175), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_148), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_12), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_30), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_157), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_139), .Y(n_292) );
BUFx2_ASAP7_75t_SL g293 ( .A(n_95), .Y(n_293) );
CKINVDCx14_ASAP7_75t_R g294 ( .A(n_213), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_90), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_223), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_16), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_169), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_132), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_39), .Y(n_300) );
BUFx10_ASAP7_75t_L g301 ( .A(n_206), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_106), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_147), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_114), .B(n_186), .Y(n_304) );
BUFx10_ASAP7_75t_L g305 ( .A(n_99), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_72), .B(n_33), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_188), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_184), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_154), .Y(n_310) );
BUFx2_ASAP7_75t_SL g311 ( .A(n_181), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_162), .Y(n_312) );
CKINVDCx14_ASAP7_75t_R g313 ( .A(n_6), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_55), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_196), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_78), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_222), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_221), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_111), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_155), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_215), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_53), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_182), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_27), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_34), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_49), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_107), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_24), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_127), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_131), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_191), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_224), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_146), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_183), .B(n_220), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_69), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_47), .B(n_16), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_25), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_199), .Y(n_338) );
BUFx10_ASAP7_75t_L g339 ( .A(n_109), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_98), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_165), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_38), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_57), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_67), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_3), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_45), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_8), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_42), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_85), .Y(n_349) );
BUFx10_ASAP7_75t_L g350 ( .A(n_18), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_56), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_159), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_12), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_41), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_233), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_17), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_120), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_92), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_229), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_128), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_37), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_174), .Y(n_362) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_84), .Y(n_363) );
BUFx5_ASAP7_75t_L g364 ( .A(n_6), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_166), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_43), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_278), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_310), .B(n_0), .Y(n_368) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_251), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_251), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_350), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_313), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_279), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_303), .Y(n_374) );
OAI22x1_ASAP7_75t_SL g375 ( .A1(n_345), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_244), .B(n_1), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_272), .B(n_2), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_289), .B(n_3), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_361), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_364), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_297), .B(n_4), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_350), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_251), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_302), .B(n_4), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_242), .A2(n_26), .B(n_23), .Y(n_385) );
AND2x6_ASAP7_75t_L g386 ( .A(n_246), .B(n_237), .Y(n_386) );
BUFx8_ASAP7_75t_SL g387 ( .A(n_267), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_325), .B(n_5), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_364), .B(n_5), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_353), .B(n_7), .Y(n_390) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_256), .Y(n_391) );
INVx6_ASAP7_75t_L g392 ( .A(n_285), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_364), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_331), .B(n_7), .Y(n_394) );
INVx4_ASAP7_75t_L g395 ( .A(n_238), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_356), .B(n_8), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_276), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_376), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_376), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_377), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_392), .B(n_277), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_380), .B(n_249), .C(n_247), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_397), .Y(n_403) );
OR2x6_ASAP7_75t_L g404 ( .A(n_372), .B(n_293), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_393), .B(n_395), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_396), .A2(n_347), .B1(n_363), .B2(n_270), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_367), .B(n_294), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
INVx6_ASAP7_75t_L g414 ( .A(n_392), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_371), .B(n_301), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_392), .B(n_341), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_371), .B(n_301), .Y(n_418) );
AND2x6_ASAP7_75t_L g419 ( .A(n_381), .B(n_252), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_373), .B(n_240), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_387), .Y(n_423) );
INVx5_ASAP7_75t_L g424 ( .A(n_419), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_415), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_410), .B(n_374), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_419), .A2(n_390), .B1(n_368), .B2(n_394), .Y(n_427) );
BUFx10_ASAP7_75t_L g428 ( .A(n_404), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_415), .B(n_379), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_405), .B(n_382), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_405), .B(n_382), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_402), .B(n_368), .C(n_384), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_400), .B(n_388), .Y(n_436) );
INVx8_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_411), .B(n_388), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_412), .B(n_389), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_414), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_402), .B(n_389), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_419), .B(n_386), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_419), .A2(n_386), .B1(n_312), .B2(n_333), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_364), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_422), .B(n_239), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_416), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_401), .B(n_417), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_407), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_418), .B(n_386), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_414), .B(n_268), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_409), .B(n_243), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_409), .B(n_248), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_423), .B(n_305), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_425), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_424), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_426), .A2(n_255), .B(n_261), .C(n_259), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_444), .A2(n_385), .B(n_263), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_441), .B(n_357), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_452), .B(n_305), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_453), .A2(n_262), .B(n_266), .C(n_264), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_424), .B(n_250), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_443), .A2(n_269), .B(n_282), .C(n_271), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_443), .A2(n_283), .B(n_287), .C(n_284), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_436), .B(n_254), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_440), .B(n_439), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_424), .B(n_257), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_445), .B(n_258), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_432), .B(n_288), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_452), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_433), .B(n_260), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_428), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g475 ( .A1(n_438), .A2(n_332), .A3(n_291), .B1(n_295), .B2(n_296), .B3(n_366), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_451), .A2(n_309), .B(n_298), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_449), .B(n_375), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_428), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_446), .B(n_265), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_435), .A2(n_321), .B(n_323), .C(n_315), .Y(n_480) );
NAND2x1_ASAP7_75t_L g481 ( .A(n_429), .B(n_256), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_448), .B(n_324), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_431), .A2(n_328), .B(n_326), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_454), .A2(n_335), .B(n_337), .C(n_329), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_434), .B(n_275), .Y(n_485) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_455), .A2(n_420), .B(n_413), .Y(n_486) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_427), .B(n_286), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_430), .B(n_290), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_447), .A2(n_342), .B(n_338), .Y(n_491) );
AOI21x1_ASAP7_75t_L g492 ( .A1(n_450), .A2(n_421), .B(n_304), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_460), .A2(n_437), .B(n_445), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_468), .B(n_437), .Y(n_494) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_458), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_461), .A2(n_245), .B1(n_334), .B2(n_273), .Y(n_496) );
CKINVDCx11_ASAP7_75t_R g497 ( .A(n_488), .Y(n_497) );
OAI21x1_ASAP7_75t_SL g498 ( .A1(n_471), .A2(n_355), .B(n_346), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_457), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_476), .A2(n_471), .B(n_473), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_475), .B(n_477), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_467), .A2(n_359), .B(n_358), .Y(n_502) );
OAI21x1_ASAP7_75t_L g503 ( .A1(n_486), .A2(n_362), .B(n_360), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_487), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_487), .B(n_292), .Y(n_505) );
AO21x1_ASAP7_75t_L g506 ( .A1(n_492), .A2(n_365), .B(n_336), .Y(n_506) );
AO22x1_ASAP7_75t_L g507 ( .A1(n_487), .A2(n_456), .B1(n_354), .B2(n_318), .Y(n_507) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_465), .A2(n_466), .A3(n_480), .B(n_483), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_459), .A2(n_281), .B(n_241), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_482), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_491), .A2(n_349), .B(n_306), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_489), .B(n_299), .Y(n_512) );
OAI21x1_ASAP7_75t_L g513 ( .A1(n_481), .A2(n_352), .B(n_307), .Y(n_513) );
OAI21xp5_ASAP7_75t_SL g514 ( .A1(n_472), .A2(n_316), .B(n_253), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_470), .B(n_300), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g516 ( .A1(n_485), .A2(n_351), .B(n_276), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_462), .B(n_339), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_458), .B(n_308), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_490), .B(n_314), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_463), .B(n_274), .C(n_256), .Y(n_520) );
AO21x1_ASAP7_75t_L g521 ( .A1(n_484), .A2(n_276), .B(n_311), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_479), .A2(n_469), .B(n_464), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_458), .A2(n_319), .B(n_317), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_474), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_478), .A2(n_322), .B(n_320), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_460), .A2(n_330), .B(n_327), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_468), .B(n_343), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_457), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_500), .A2(n_348), .B(n_344), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_501), .A2(n_339), .B1(n_276), .B2(n_340), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_528), .Y(n_531) );
NOR2xp67_ASAP7_75t_SL g532 ( .A(n_495), .B(n_280), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_495), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_499), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_497), .Y(n_535) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_514), .B(n_383), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_510), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_503), .A2(n_391), .B(n_383), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_504), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_495), .Y(n_541) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_513), .A2(n_35), .B(n_31), .Y(n_542) );
AO31x2_ASAP7_75t_L g543 ( .A1(n_506), .A2(n_9), .A3(n_10), .B(n_11), .Y(n_543) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_498), .A2(n_40), .B(n_36), .Y(n_544) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_527), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_496), .B(n_9), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_517), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_547) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_493), .A2(n_144), .B(n_235), .Y(n_548) );
INVx2_ASAP7_75t_SL g549 ( .A(n_524), .Y(n_549) );
OAI21x1_ASAP7_75t_L g550 ( .A1(n_526), .A2(n_143), .B(n_234), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_502), .A2(n_17), .B(n_18), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_507), .B(n_19), .Y(n_552) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_521), .A2(n_149), .B(n_230), .Y(n_553) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_522), .A2(n_145), .B(n_226), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_508), .Y(n_555) );
BUFx8_ASAP7_75t_L g556 ( .A(n_505), .Y(n_556) );
NOR2xp33_ASAP7_75t_SL g557 ( .A(n_516), .B(n_20), .Y(n_557) );
INVx4_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_508), .B(n_21), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_523), .B(n_46), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_508), .Y(n_561) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_512), .A2(n_48), .A3(n_50), .B(n_59), .Y(n_562) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_511), .A2(n_61), .B(n_62), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_509), .B(n_63), .Y(n_565) );
OAI21x1_ASAP7_75t_SL g566 ( .A1(n_525), .A2(n_519), .B(n_515), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_494), .B(n_65), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_500), .A2(n_68), .B(n_70), .C(n_71), .Y(n_568) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_495), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_494), .B(n_73), .Y(n_570) );
AO21x1_ASAP7_75t_L g571 ( .A1(n_493), .A2(n_74), .B(n_76), .Y(n_571) );
OAI222xp33_ASAP7_75t_L g572 ( .A1(n_501), .A2(n_77), .B1(n_79), .B2(n_80), .C1(n_81), .C2(n_83), .Y(n_572) );
AO21x1_ASAP7_75t_L g573 ( .A1(n_493), .A2(n_86), .B(n_89), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_501), .A2(n_91), .B1(n_94), .B2(n_96), .Y(n_574) );
OR2x6_ASAP7_75t_L g575 ( .A(n_494), .B(n_97), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_534), .B(n_100), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_537), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_575), .Y(n_578) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_559), .A2(n_101), .B(n_103), .Y(n_579) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_536), .B(n_105), .Y(n_580) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_533), .Y(n_581) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_555), .A2(n_108), .B(n_110), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_538), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_555), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_561), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_540), .B(n_236), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_561), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_543), .Y(n_589) );
INVxp67_ASAP7_75t_SL g590 ( .A(n_533), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_543), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_570), .B(n_116), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_545), .A2(n_117), .B1(n_119), .B2(n_121), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_556), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_122), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_552), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_558), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_551), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_549), .B(n_129), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_556), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_535), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_557), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_133), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_566), .A2(n_134), .B(n_137), .C(n_140), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_547), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_542), .Y(n_609) );
OAI21x1_ASAP7_75t_L g610 ( .A1(n_539), .A2(n_141), .B(n_142), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_529), .B(n_150), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_567), .A2(n_151), .B1(n_153), .B2(n_156), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_565), .B(n_161), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_548), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_553), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_560), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_530), .B(n_163), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_571), .B(n_164), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_564), .Y(n_620) );
OR2x6_ASAP7_75t_L g621 ( .A(n_550), .B(n_167), .Y(n_621) );
AO21x2_ASAP7_75t_L g622 ( .A1(n_573), .A2(n_168), .B(n_171), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_554), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_563), .Y(n_624) );
OR2x6_ASAP7_75t_L g625 ( .A(n_568), .B(n_172), .Y(n_625) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_553), .A2(n_177), .B(n_178), .Y(n_626) );
AO21x2_ASAP7_75t_L g627 ( .A1(n_572), .A2(n_564), .B(n_532), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_532), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_574), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_534), .Y(n_630) );
OA21x2_ASAP7_75t_L g631 ( .A1(n_555), .A2(n_179), .B(n_180), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_538), .B(n_185), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_534), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_531), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_534), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_534), .B(n_225), .Y(n_636) );
AOI211xp5_ASAP7_75t_SL g637 ( .A1(n_572), .A2(n_187), .B(n_189), .C(n_192), .Y(n_637) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_533), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_538), .B(n_193), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_534), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_534), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_597), .B(n_194), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_583), .B(n_195), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_630), .B(n_198), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_605), .Y(n_646) );
AND2x4_ASAP7_75t_L g647 ( .A(n_578), .B(n_200), .Y(n_647) );
INVx3_ASAP7_75t_L g648 ( .A(n_593), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_633), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_602), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_578), .B(n_201), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_635), .Y(n_652) );
INVx4_ASAP7_75t_R g653 ( .A(n_595), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_640), .B(n_203), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_590), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_600), .B(n_205), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_642), .B(n_207), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_577), .B(n_208), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_634), .B(n_209), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_599), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
INVx4_ASAP7_75t_L g663 ( .A(n_593), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_581), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_585), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_588), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_598), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_598), .B(n_210), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_591), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_576), .Y(n_670) );
NOR2x1_ASAP7_75t_SL g671 ( .A(n_606), .B(n_212), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_587), .Y(n_672) );
INVx3_ASAP7_75t_L g673 ( .A(n_581), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_589), .B(n_217), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_636), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_620), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_638), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_632), .B(n_639), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_617), .B(n_620), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_586), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_620), .Y(n_682) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_617), .B(n_601), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_592), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_596), .B(n_608), .Y(n_685) );
BUFx6f_ASAP7_75t_L g686 ( .A(n_628), .Y(n_686) );
INVxp67_ASAP7_75t_L g687 ( .A(n_580), .Y(n_687) );
BUFx3_ASAP7_75t_L g688 ( .A(n_603), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_618), .B(n_614), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_579), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_627), .B(n_612), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_580), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_582), .B(n_631), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_611), .B(n_629), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_610), .Y(n_695) );
INVx5_ASAP7_75t_L g696 ( .A(n_621), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_594), .B(n_629), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_604), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_637), .B(n_613), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_615), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_625), .B(n_621), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_625), .A2(n_621), .B1(n_622), .B2(n_616), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_625), .B(n_622), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_607), .B(n_619), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_607), .Y(n_705) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_624), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_699), .A2(n_623), .B1(n_609), .B2(n_626), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_649), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_652), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_655), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_696), .B(n_701), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_667), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_696), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_662), .B(n_665), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_666), .B(n_684), .Y(n_715) );
INVx5_ASAP7_75t_L g716 ( .A(n_696), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_706), .B(n_672), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_706), .B(n_672), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_661), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_698), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_646), .B(n_656), .Y(n_721) );
AND2x4_ASAP7_75t_L g722 ( .A(n_696), .B(n_691), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_669), .B(n_700), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_685), .B(n_681), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_677), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_700), .B(n_703), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_670), .B(n_676), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_648), .B(n_663), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_686), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_682), .B(n_686), .Y(n_730) );
BUFx3_ASAP7_75t_L g731 ( .A(n_674), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_682), .B(n_694), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_663), .B(n_679), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_688), .B(n_680), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_689), .B(n_697), .Y(n_735) );
INVx4_ASAP7_75t_L g736 ( .A(n_668), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_643), .B(n_683), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_675), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_650), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_675), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_702), .B(n_705), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_647), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_668), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_643), .B(n_658), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_690), .B(n_704), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_650), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_664), .B(n_678), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_647), .Y(n_748) );
INVxp67_ASAP7_75t_L g749 ( .A(n_651), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_673), .B(n_692), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_687), .B(n_693), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_653), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_711), .B(n_695), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_719), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_736), .B(n_695), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_708), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_733), .B(n_683), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_735), .B(n_659), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_739), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_711), .B(n_671), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_724), .B(n_654), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_709), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_710), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_746), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_732), .B(n_645), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_720), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_727), .B(n_644), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_715), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_712), .B(n_660), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_715), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_714), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_714), .Y(n_772) );
INVx4_ASAP7_75t_L g773 ( .A(n_736), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_749), .B(n_657), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_711), .B(n_653), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_742), .B(n_748), .Y(n_776) );
AND2x4_ASAP7_75t_L g777 ( .A(n_722), .B(n_751), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_726), .B(n_730), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_754), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_759), .Y(n_780) );
NAND3x1_ASAP7_75t_L g781 ( .A(n_757), .B(n_752), .C(n_713), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_768), .B(n_741), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_773), .B(n_721), .Y(n_783) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_764), .B(n_734), .Y(n_784) );
NAND2xp67_ASAP7_75t_SL g785 ( .A(n_769), .B(n_721), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_770), .B(n_723), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_766), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_773), .B(n_751), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_771), .B(n_741), .Y(n_789) );
OR2x6_ASAP7_75t_L g790 ( .A(n_775), .B(n_743), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_778), .B(n_777), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_772), .B(n_777), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_756), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_762), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_763), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_782), .B(n_717), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_795), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_795), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_789), .B(n_718), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_779), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_791), .B(n_777), .Y(n_801) );
OAI21xp33_ASAP7_75t_L g802 ( .A1(n_780), .A2(n_774), .B(n_776), .Y(n_802) );
AOI32xp33_ASAP7_75t_L g803 ( .A1(n_783), .A2(n_737), .A3(n_760), .B1(n_765), .B2(n_774), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_781), .A2(n_755), .B(n_760), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_784), .B(n_776), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_787), .B(n_717), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_797), .Y(n_807) );
INVxp67_ASAP7_75t_L g808 ( .A(n_800), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_798), .Y(n_809) );
INVx1_ASAP7_75t_SL g810 ( .A(n_801), .Y(n_810) );
OAI21xp5_ASAP7_75t_SL g811 ( .A1(n_804), .A2(n_788), .B(n_785), .Y(n_811) );
INVx1_ASAP7_75t_SL g812 ( .A(n_806), .Y(n_812) );
OAI322xp33_ASAP7_75t_L g813 ( .A1(n_805), .A2(n_794), .A3(n_793), .B1(n_761), .B2(n_767), .C1(n_758), .C2(n_792), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_813), .A2(n_802), .B1(n_803), .B2(n_799), .C(n_796), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g815 ( .A(n_811), .B(n_802), .C(n_728), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_813), .A2(n_790), .B(n_716), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_808), .A2(n_716), .B(n_744), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_810), .A2(n_786), .B1(n_716), .B2(n_713), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_814), .B(n_812), .Y(n_819) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_816), .B(n_807), .Y(n_820) );
NOR3xp33_ASAP7_75t_SL g821 ( .A(n_818), .B(n_809), .C(n_740), .Y(n_821) );
OAI21xp33_ASAP7_75t_L g822 ( .A1(n_819), .A2(n_815), .B(n_817), .Y(n_822) );
NAND5xp2_ASAP7_75t_L g823 ( .A(n_821), .B(n_707), .C(n_745), .D(n_738), .E(n_750), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_822), .B(n_820), .Y(n_824) );
NOR2xp67_ASAP7_75t_L g825 ( .A(n_824), .B(n_823), .Y(n_825) );
INVx2_ASAP7_75t_SL g826 ( .A(n_825), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_826), .A2(n_716), .B1(n_713), .B2(n_731), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_827), .A2(n_716), .B(n_745), .Y(n_828) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_828), .B(n_731), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_829), .A2(n_725), .B(n_747), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_830), .B(n_729), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_831), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_832), .B(n_753), .Y(n_833) );
endmodule