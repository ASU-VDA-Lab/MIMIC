module real_jpeg_28119_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_302, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_302;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_221;
wire n_288;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_295;
wire n_128;
wire n_244;
wire n_179;
wire n_167;
wire n_133;
wire n_202;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_0),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_0),
.A2(n_32),
.B1(n_34),
.B2(n_53),
.Y(n_227)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_32),
.B1(n_34),
.B2(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_72),
.B1(n_73),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_32),
.B1(n_34),
.B2(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_121),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_121),
.Y(n_240)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_45),
.B1(n_72),
.B2(n_73),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_5),
.A2(n_32),
.B1(n_34),
.B2(n_45),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_6),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_75),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_32),
.B1(n_34),
.B2(n_75),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_75),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_26),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_25),
.B(n_26),
.C(n_134),
.D(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_47),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_10),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_83),
.B(n_151),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_43),
.B(n_46),
.C(n_184),
.D(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_10),
.B(n_43),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_68),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_70),
.B(n_73),
.C(n_229),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_10),
.A2(n_72),
.B1(n_73),
.B2(n_166),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_11),
.A2(n_72),
.B1(n_73),
.B2(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_11),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_98),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_32),
.B1(n_34),
.B2(n_98),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_98),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_12),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_12),
.A2(n_32),
.B1(n_34),
.B2(n_146),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_12),
.A2(n_72),
.B1(n_73),
.B2(n_146),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_13),
.A2(n_26),
.B(n_28),
.C(n_31),
.Y(n_25)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_32),
.Y(n_135)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_16),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_99),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_80),
.B2(n_81),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_54),
.B1(n_55),
.B2(n_79),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_23),
.A2(n_24),
.B(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_25),
.A2(n_31),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_25),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_25),
.A2(n_31),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_26),
.A2(n_44),
.A3(n_184),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_27),
.A2(n_30),
.A3(n_34),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_27),
.B(n_196),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_32),
.B(n_84),
.Y(n_83)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_34),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_42),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_43),
.A2(n_69),
.B(n_166),
.Y(n_229)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_47),
.B1(n_52),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_46),
.B(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_46),
.A2(n_47),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_78),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_61),
.A2(n_62),
.B1(n_93),
.B2(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_61),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_61),
.A2(n_62),
.B1(n_113),
.B2(n_243),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_62),
.B(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_62),
.A2(n_145),
.B(n_147),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_62),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_62),
.A2(n_147),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_66),
.A2(n_119),
.B(n_122),
.Y(n_118)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_67),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_67),
.A2(n_68),
.B1(n_120),
.B2(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_97),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_76),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_76),
.A2(n_96),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B(n_94),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_94),
.B1(n_95),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_103),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_88),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_83),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_83),
.B(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_83),
.A2(n_87),
.B1(n_193),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_83),
.A2(n_87),
.B1(n_110),
.B2(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_85),
.A2(n_158),
.B(n_168),
.Y(n_167)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_86),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_169),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_86),
.A2(n_159),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_106),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_289)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_106),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.C(n_118),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_107),
.A2(n_108),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_109),
.B(n_112),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_114),
.B(n_118),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_115),
.A2(n_253),
.B(n_254),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_116),
.A2(n_117),
.B(n_205),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_117),
.B(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_117),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_281),
.A3(n_290),
.B1(n_295),
.B2(n_300),
.C(n_302),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_245),
.C(n_277),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_219),
.B(n_244),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_199),
.B(n_218),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_179),
.B(n_198),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_154),
.B(n_178),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_139),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_144),
.C(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_163),
.B(n_177),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_170),
.B(n_176),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_181),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_190),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_187),
.C(n_190),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_194),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_214),
.C(n_215),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_208),
.C(n_211),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_232),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_224),
.C(n_232),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_238),
.C(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_246),
.A2(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_247),
.B(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.C(n_263),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_251),
.C(n_258),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_258),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_263),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_273),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_273),
.C(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_288),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.C(n_287),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_296),
.B(n_299),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_293),
.Y(n_299)
);


endmodule