module fake_ariane_2223_n_756 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_756);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_756;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_699;
wire n_727;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_52),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_0),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_9),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_47),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_11),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_53),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_85),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_128),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_49),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_L g178 ( 
.A(n_73),
.B(n_123),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_36),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_25),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_21),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_28),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_113),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_90),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_82),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_39),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_42),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_10),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_156),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_27),
.B(n_2),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_0),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_3),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

AOI22x1_ASAP7_75t_SL g225 ( 
.A1(n_164),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_6),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_7),
.Y(n_236)
);

OAI22x1_ASAP7_75t_SL g237 ( 
.A1(n_159),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_237)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_171),
.B(n_12),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_12),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_159),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_194),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_16),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_187),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_197),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

NAND2xp33_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_162),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_182),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_209),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_183),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_252),
.B(n_161),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_165),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_242),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_215),
.B(n_184),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_220),
.A2(n_213),
.B(n_212),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_188),
.B1(n_207),
.B2(n_206),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_238),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g285 ( 
.A1(n_248),
.A2(n_198),
.B(n_200),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_238),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_217),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_199),
.B1(n_176),
.B2(n_178),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_234),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_228),
.B(n_169),
.Y(n_293)
);

CKINVDCx6p67_ASAP7_75t_R g294 ( 
.A(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_215),
.B(n_172),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_231),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g297 ( 
.A(n_214),
.B(n_210),
.C(n_205),
.Y(n_297)
);

OR2x6_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_16),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_217),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_174),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_247),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_261),
.B(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_235),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_221),
.C(n_233),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_257),
.A2(n_228),
.B(n_243),
.C(n_236),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_239),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_236),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_240),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_240),
.B1(n_243),
.B2(n_256),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_223),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_223),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_291),
.A2(n_237),
.B1(n_245),
.B2(n_180),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_223),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_259),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_226),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_226),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_287),
.B(n_177),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_293),
.B(n_226),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_253),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_239),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_259),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_287),
.B(n_190),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_269),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_274),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g344 ( 
.A(n_266),
.B(n_232),
.C(n_225),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

BUFx6f_ASAP7_75t_SL g346 ( 
.A(n_298),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_253),
.Y(n_348)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_259),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_286),
.B(n_241),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_259),
.A2(n_192),
.B1(n_196),
.B2(n_201),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_268),
.B(n_255),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_260),
.B(n_255),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_241),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_297),
.B(n_255),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_255),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_294),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_258),
.B(n_255),
.Y(n_361)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_258),
.A2(n_305),
.B(n_301),
.C(n_299),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_298),
.A2(n_225),
.B1(n_227),
.B2(n_224),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_280),
.B(n_218),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_280),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_218),
.Y(n_368)
);

OR2x6_ASAP7_75t_SL g369 ( 
.A(n_298),
.B(n_17),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_285),
.B(n_218),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_305),
.B(n_301),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_313),
.A2(n_299),
.B(n_290),
.C(n_288),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_311),
.A2(n_259),
.B(n_288),
.C(n_284),
.Y(n_373)
);

INVx11_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_259),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_320),
.A2(n_290),
.B(n_284),
.C(n_279),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_279),
.B1(n_275),
.B2(n_273),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_SL g378 ( 
.A(n_312),
.B(n_17),
.C(n_18),
.Y(n_378)
);

NAND2x1_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_273),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_275),
.B(n_269),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_327),
.B(n_323),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_319),
.A2(n_269),
.B(n_227),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_331),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

OAI321xp33_ASAP7_75t_L g386 ( 
.A1(n_363),
.A2(n_227),
.A3(n_224),
.B1(n_269),
.B2(n_18),
.C(n_19),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_310),
.B(n_224),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_333),
.A2(n_227),
.B(n_224),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_224),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_346),
.A2(n_227),
.B1(n_19),
.B2(n_22),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_348),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_20),
.B(n_23),
.C(n_24),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_26),
.B(n_29),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_308),
.A2(n_30),
.B(n_31),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_345),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_332),
.B(n_32),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_308),
.A2(n_33),
.B(n_34),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_343),
.B(n_157),
.Y(n_400)
);

NAND2x1p5_ASAP7_75t_L g401 ( 
.A(n_307),
.B(n_329),
.Y(n_401)
);

CKINVDCx6p67_ASAP7_75t_R g402 ( 
.A(n_360),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_35),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_155),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_309),
.A2(n_37),
.B(n_38),
.C(n_40),
.Y(n_407)
);

O2A1O1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_326),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_339),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_309),
.A2(n_314),
.B(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_338),
.B(n_152),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_352),
.B(n_54),
.Y(n_414)
);

NOR2x1p5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_149),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_335),
.B(n_55),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_349),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_351),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_351),
.B(n_148),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_356),
.A2(n_64),
.B(n_66),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_337),
.A2(n_67),
.B(n_68),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_69),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_147),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_359),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_426)
);

O2A1O1Ixp33_ASAP7_75t_L g427 ( 
.A1(n_358),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_359),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_315),
.A2(n_86),
.B(n_87),
.Y(n_429)
);

BUFx4f_ASAP7_75t_L g430 ( 
.A(n_360),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_316),
.B(n_88),
.C(n_92),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_328),
.B(n_94),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_322),
.B(n_98),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_355),
.B(n_146),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_99),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_145),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_370),
.B(n_100),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_143),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_325),
.B(n_101),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_L g441 ( 
.A(n_342),
.B(n_103),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_362),
.B(n_344),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_410),
.A2(n_365),
.B(n_367),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_364),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_347),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_390),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_371),
.A2(n_361),
.B(n_347),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_375),
.A2(n_347),
.B(n_342),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_379),
.A2(n_106),
.B(n_107),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_392),
.B(n_109),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_390),
.B(n_112),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

AO31x2_ASAP7_75t_L g454 ( 
.A1(n_438),
.A2(n_114),
.A3(n_117),
.B(n_118),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_383),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_385),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_373),
.A2(n_124),
.B(n_125),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_430),
.B(n_127),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_417),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_140),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_129),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_416),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_462)
);

CKINVDCx6p67_ASAP7_75t_R g463 ( 
.A(n_433),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_134),
.B(n_135),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_396),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_437),
.A2(n_136),
.B(n_137),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_417),
.B(n_138),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_139),
.B(n_421),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_413),
.A2(n_380),
.B(n_394),
.Y(n_471)
);

AO31x2_ASAP7_75t_L g472 ( 
.A1(n_376),
.A2(n_428),
.A3(n_425),
.B(n_405),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_381),
.A2(n_389),
.B(n_372),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_374),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_435),
.A2(n_434),
.B(n_440),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_397),
.A2(n_400),
.B(n_388),
.Y(n_476)
);

OAI21x1_ASAP7_75t_SL g477 ( 
.A1(n_391),
.A2(n_409),
.B(n_408),
.Y(n_477)
);

OAI21xp33_ASAP7_75t_L g478 ( 
.A1(n_378),
.A2(n_424),
.B(n_391),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_382),
.A2(n_414),
.B(n_387),
.Y(n_479)
);

AO21x1_ASAP7_75t_L g480 ( 
.A1(n_418),
.A2(n_423),
.B(n_420),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_426),
.A2(n_431),
.B1(n_399),
.B2(n_412),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_401),
.B(n_431),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_395),
.A2(n_422),
.B(n_398),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_407),
.A2(n_393),
.B(n_377),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_431),
.A2(n_430),
.B1(n_415),
.B2(n_386),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_432),
.B(n_429),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_441),
.A2(n_410),
.B(n_371),
.Y(n_487)
);

NAND2x1_ASAP7_75t_L g488 ( 
.A(n_390),
.B(n_417),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_390),
.B(n_327),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_416),
.A2(n_313),
.B(n_257),
.C(n_424),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_419),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_410),
.A2(n_375),
.B(n_373),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_410),
.A2(n_371),
.B(n_366),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_410),
.A2(n_371),
.B(n_366),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_384),
.B(n_385),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_471),
.A2(n_492),
.B(n_493),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_495),
.A2(n_487),
.B(n_476),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_483),
.A2(n_475),
.B(n_448),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_478),
.A2(n_467),
.B1(n_461),
.B2(n_465),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_490),
.B(n_444),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_446),
.Y(n_503)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_457),
.A2(n_484),
.B(n_486),
.Y(n_504)
);

O2A1O1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_478),
.A2(n_477),
.B(n_456),
.C(n_485),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_461),
.Y(n_506)
);

AOI222xp33_ASAP7_75t_L g507 ( 
.A1(n_458),
.A2(n_494),
.B1(n_464),
.B2(n_443),
.C1(n_453),
.C2(n_484),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_445),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_496),
.B1(n_443),
.B2(n_453),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_479),
.A2(n_449),
.B(n_473),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_482),
.B(n_442),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_462),
.A2(n_466),
.B(n_468),
.C(n_450),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_480),
.B(n_481),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_474),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_474),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_451),
.A2(n_489),
.B1(n_442),
.B2(n_470),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_452),
.A2(n_455),
.B(n_488),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_SL g518 ( 
.A1(n_472),
.A2(n_447),
.B(n_459),
.C(n_470),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

AOI221xp5_ASAP7_75t_L g520 ( 
.A1(n_469),
.A2(n_311),
.B1(n_257),
.B2(n_281),
.C(n_478),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_454),
.Y(n_521)
);

AO21x2_ASAP7_75t_L g522 ( 
.A1(n_472),
.A2(n_492),
.B(n_477),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_472),
.B(n_458),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_461),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_471),
.A2(n_492),
.B(n_493),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_490),
.A2(n_492),
.B(n_491),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_471),
.A2(n_492),
.B(n_493),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_461),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_478),
.A2(n_490),
.B(n_313),
.C(n_386),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_458),
.B(n_491),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_490),
.A2(n_492),
.B(n_491),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_464),
.Y(n_532)
);

AO32x2_ASAP7_75t_L g533 ( 
.A1(n_485),
.A2(n_481),
.A3(n_428),
.B1(n_409),
.B2(n_418),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_491),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_478),
.B(n_490),
.C(n_257),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_474),
.B(n_461),
.Y(n_536)
);

NAND2x1p5_ASAP7_75t_L g537 ( 
.A(n_442),
.B(n_458),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_458),
.B(n_491),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_491),
.B(n_467),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_471),
.A2(n_492),
.B(n_493),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_505),
.A2(n_529),
.B(n_535),
.C(n_513),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_526),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_532),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_520),
.B(n_513),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_538),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_528),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_514),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_522),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

O2A1O1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_534),
.B(n_538),
.C(n_530),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_499),
.A2(n_498),
.B(n_527),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_539),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_511),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_504),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_530),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_502),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_534),
.B(n_536),
.Y(n_565)
);

A2O1A1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_501),
.A2(n_509),
.B(n_516),
.C(n_512),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_504),
.A2(n_507),
.B(n_512),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_524),
.Y(n_571)
);

AO21x2_ASAP7_75t_L g572 ( 
.A1(n_518),
.A2(n_540),
.B(n_527),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_551),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_537),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_537),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_558),
.B(n_533),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_543),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_552),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_551),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_533),
.Y(n_583)
);

BUFx12f_ASAP7_75t_L g584 ( 
.A(n_550),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_533),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_533),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_569),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_536),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_542),
.B(n_536),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_543),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_547),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_545),
.B(n_499),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_553),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_545),
.B(n_510),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_519),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_553),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_544),
.B(n_500),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_550),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_500),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_546),
.B(n_517),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_543),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_515),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_517),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_549),
.B(n_565),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_562),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_561),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_571),
.B(n_550),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_571),
.B(n_560),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_567),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_606),
.B(n_559),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_556),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_576),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_607),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_579),
.B(n_568),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_602),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_581),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_602),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_608),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_607),
.B(n_568),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_610),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_576),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_579),
.B(n_567),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_587),
.B(n_570),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_583),
.B(n_585),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_591),
.B(n_555),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_591),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_588),
.B(n_589),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_584),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_587),
.B(n_575),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_582),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_589),
.B(n_541),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_585),
.B(n_570),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_600),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_574),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_600),
.B(n_572),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_609),
.B(n_573),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_597),
.B(n_599),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_597),
.B(n_572),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_598),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_604),
.B(n_566),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_635),
.B(n_594),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_635),
.B(n_594),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_615),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_617),
.B(n_605),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_633),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_622),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_614),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_614),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_628),
.B(n_605),
.Y(n_651)
);

NAND2x1_ASAP7_75t_L g652 ( 
.A(n_641),
.B(n_601),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_626),
.B(n_611),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_639),
.B(n_592),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_619),
.B(n_626),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_623),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_639),
.B(n_592),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_634),
.B(n_604),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_629),
.B(n_611),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_632),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_634),
.B(n_603),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_627),
.A2(n_603),
.B(n_595),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_636),
.B(n_593),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_620),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_621),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_624),
.Y(n_667)
);

AOI32xp33_ASAP7_75t_L g668 ( 
.A1(n_642),
.A2(n_578),
.A3(n_595),
.B1(n_609),
.B2(n_598),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_612),
.B(n_598),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_636),
.B(n_596),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_632),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_625),
.B(n_596),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_647),
.B(n_645),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_667),
.B(n_637),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_666),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_669),
.B(n_618),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_672),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_667),
.B(n_630),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_649),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_650),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_653),
.B(n_625),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_653),
.B(n_631),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_643),
.B(n_637),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_652),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_654),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_643),
.B(n_640),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_651),
.A2(n_642),
.B(n_631),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_665),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_656),
.A2(n_613),
.B1(n_578),
.B2(n_577),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_651),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_682),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_684),
.B(n_644),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_685),
.B(n_668),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_680),
.Y(n_695)
);

NOR2x1_ASAP7_75t_L g696 ( 
.A(n_685),
.B(n_672),
.Y(n_696)
);

OAI322xp33_ASAP7_75t_L g697 ( 
.A1(n_678),
.A2(n_660),
.A3(n_646),
.B1(n_671),
.B2(n_657),
.C1(n_661),
.C2(n_670),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_676),
.B(n_630),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_644),
.Y(n_699)
);

AO22x1_ASAP7_75t_L g700 ( 
.A1(n_691),
.A2(n_630),
.B1(n_648),
.B2(n_663),
.Y(n_700)
);

NAND2x1p5_ASAP7_75t_L g701 ( 
.A(n_678),
.B(n_641),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_680),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_695),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_673),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_SL g705 ( 
.A1(n_694),
.A2(n_688),
.B(n_679),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_698),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_698),
.B(n_683),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_693),
.B(n_674),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_700),
.B(n_674),
.Y(n_709)
);

OAI211xp5_ASAP7_75t_SL g710 ( 
.A1(n_705),
.A2(n_696),
.B(n_702),
.C(n_686),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_709),
.A2(n_697),
.B1(n_690),
.B2(n_681),
.C(n_686),
.Y(n_711)
);

NAND4xp25_ASAP7_75t_L g712 ( 
.A(n_703),
.B(n_681),
.C(n_666),
.D(n_699),
.Y(n_712)
);

AOI211xp5_ASAP7_75t_L g713 ( 
.A1(n_707),
.A2(n_697),
.B(n_683),
.C(n_662),
.Y(n_713)
);

OA22x2_ASAP7_75t_L g714 ( 
.A1(n_706),
.A2(n_684),
.B1(n_687),
.B2(n_662),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_714),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_711),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_712),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_713),
.A2(n_710),
.B1(n_704),
.B2(n_708),
.C(n_687),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_714),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_716),
.Y(n_720)
);

NAND4xp25_ASAP7_75t_L g721 ( 
.A(n_717),
.B(n_666),
.C(n_621),
.D(n_655),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_719),
.B(n_548),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_720),
.B(n_715),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_721),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_722),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_718),
.C(n_548),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

XNOR2x1_ASAP7_75t_L g728 ( 
.A(n_724),
.B(n_701),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_726),
.B(n_675),
.Y(n_729)
);

XNOR2x1_ASAP7_75t_L g730 ( 
.A(n_725),
.B(n_577),
.Y(n_730)
);

XNOR2xp5_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_595),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_725),
.B(n_555),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_727),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_731),
.A2(n_730),
.B1(n_728),
.B2(n_732),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_731),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_729),
.A2(n_584),
.B1(n_595),
.B2(n_677),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_727),
.B(n_548),
.C(n_670),
.Y(n_737)
);

AOI22x1_ASAP7_75t_L g738 ( 
.A1(n_727),
.A2(n_548),
.B1(n_658),
.B2(n_655),
.Y(n_738)
);

AO22x2_ASAP7_75t_L g739 ( 
.A1(n_727),
.A2(n_689),
.B1(n_677),
.B2(n_580),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_733),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_739),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_738),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_734),
.B(n_638),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_658),
.Y(n_744)
);

OA21x2_ASAP7_75t_L g745 ( 
.A1(n_740),
.A2(n_735),
.B(n_736),
.Y(n_745)
);

OAI22x1_ASAP7_75t_L g746 ( 
.A1(n_742),
.A2(n_741),
.B1(n_743),
.B2(n_744),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_659),
.Y(n_748)
);

OA21x2_ASAP7_75t_L g749 ( 
.A1(n_740),
.A2(n_689),
.B(n_557),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_659),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_746),
.A2(n_555),
.B(n_590),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_750),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_748),
.B1(n_745),
.B2(n_749),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_753),
.B(n_555),
.Y(n_754)
);

OR2x6_ASAP7_75t_L g755 ( 
.A(n_754),
.B(n_752),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_755),
.A2(n_584),
.B1(n_555),
.B2(n_664),
.Y(n_756)
);


endmodule