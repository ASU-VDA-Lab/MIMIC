module fake_jpeg_24327_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_44),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_35),
.B1(n_23),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_51),
.B1(n_69),
.B2(n_30),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_35),
.B1(n_23),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_35),
.B1(n_23),
.B2(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_55),
.B(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_34),
.B1(n_33),
.B2(n_18),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_61),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_67),
.B1(n_68),
.B2(n_20),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_64),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_25),
.B1(n_18),
.B2(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_71),
.B(n_78),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_84),
.Y(n_111)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_32),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_38),
.B(n_41),
.C(n_45),
.Y(n_81)
);

OAI21x1_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_87),
.B(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_29),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_29),
.B(n_28),
.C(n_17),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_93),
.B1(n_96),
.B2(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_102),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_19),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_22),
.Y(n_95)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_97),
.Y(n_112)
);

NOR4xp25_ASAP7_75t_SL g98 ( 
.A(n_50),
.B(n_15),
.C(n_16),
.D(n_14),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_107),
.C(n_53),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_41),
.B(n_27),
.C(n_21),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_106),
.B1(n_70),
.B2(n_59),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_50),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_45),
.B1(n_44),
.B2(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_40),
.B1(n_36),
.B2(n_21),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_44),
.B1(n_40),
.B2(n_36),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_21),
.B(n_17),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_108),
.A2(n_115),
.B1(n_44),
.B2(n_104),
.Y(n_163)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_123),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_70),
.B1(n_45),
.B2(n_17),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_103),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_77),
.B1(n_79),
.B2(n_102),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_94),
.B(n_101),
.Y(n_152)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_133),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_11),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_130),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_40),
.B1(n_36),
.B2(n_92),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_12),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_40),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_80),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_86),
.B1(n_81),
.B2(n_75),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_138),
.A2(n_31),
.B1(n_26),
.B2(n_22),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_139),
.A2(n_150),
.B1(n_163),
.B2(n_168),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_105),
.B(n_81),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_151),
.B(n_40),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_125),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_154),
.Y(n_192)
);

AOI22x1_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_87),
.B1(n_99),
.B2(n_107),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_125),
.B1(n_134),
.B2(n_36),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_159),
.B(n_160),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_98),
.B1(n_88),
.B2(n_100),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_122),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_36),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_157),
.B1(n_162),
.B2(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_90),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_118),
.B(n_83),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_129),
.C(n_118),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_169),
.B(n_170),
.C(n_179),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_129),
.C(n_117),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_132),
.B1(n_130),
.B2(n_127),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_194),
.B1(n_143),
.B2(n_144),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_147),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_176),
.A2(n_183),
.B(n_196),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_112),
.C(n_114),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_188),
.C(n_26),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_187),
.Y(n_221)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_186),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_31),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_134),
.B1(n_112),
.B2(n_31),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_166),
.B1(n_165),
.B2(n_141),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_26),
.B1(n_31),
.B2(n_97),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_0),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_148),
.A2(n_10),
.B(n_16),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_9),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_22),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_196),
.B1(n_183),
.B2(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_214),
.B1(n_223),
.B2(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_206),
.B(n_208),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_138),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_222),
.B(n_228),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_178),
.B(n_164),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_227),
.B1(n_195),
.B2(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_182),
.C(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_175),
.B(n_8),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_221),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_235),
.C(n_242),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_170),
.C(n_188),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_227),
.B1(n_220),
.B2(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_176),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_240),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_222),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_196),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_216),
.B(n_208),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_186),
.C(n_171),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_201),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_213),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_172),
.C(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_248),
.C(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_173),
.C(n_195),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_263),
.C(n_230),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_241),
.A2(n_216),
.B(n_219),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_241),
.B(n_233),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_202),
.C(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_262),
.C(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_265),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_206),
.B1(n_225),
.B2(n_213),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_212),
.C(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_267),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_238),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_276),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_9),
.B(n_10),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_274),
.C(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_234),
.C(n_242),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_229),
.C(n_248),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_246),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_236),
.CI(n_215),
.CON(n_279),
.SN(n_279)
);

A2O1A1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_260),
.B(n_268),
.C(n_261),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_283),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_177),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_284),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_256),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_177),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_252),
.B(n_251),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_292),
.B(n_296),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_228),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_279),
.Y(n_299)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_120),
.B(n_6),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_272),
.C(n_274),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_304),
.C(n_5),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_291),
.A2(n_279),
.B(n_282),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_120),
.B(n_191),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_310),
.B(n_4),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_285),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_308),
.A3(n_12),
.B1(n_14),
.B2(n_13),
.C1(n_3),
.C2(n_0),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_285),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_285),
.B1(n_292),
.B2(n_6),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_312),
.C(n_4),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_5),
.B(n_14),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_305),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_314),
.A3(n_315),
.B1(n_316),
.B2(n_308),
.C1(n_311),
.C2(n_13),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_22),
.C2(n_304),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_1),
.B(n_2),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_1),
.Y(n_321)
);


endmodule