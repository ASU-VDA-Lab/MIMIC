module fake_jpeg_12495_n_92 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_37),
.C(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_36),
.B1(n_30),
.B2(n_29),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_49),
.C(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_37),
.B1(n_38),
.B2(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_4),
.Y(n_73)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_5),
.B(n_10),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_20),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_16),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_75),
.B1(n_77),
.B2(n_83),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_86),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_88),
.B(n_80),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_85),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_74),
.Y(n_92)
);


endmodule