module fake_jpeg_17308_n_357 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_357);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_271;
wire n_67;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_58),
.Y(n_71)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_28),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_78),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_28),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_20),
.B(n_41),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_37),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_81),
.B1(n_64),
.B2(n_58),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_41),
.B1(n_42),
.B2(n_35),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_101),
.B1(n_106),
.B2(n_118),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_114),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_104),
.B1(n_107),
.B2(n_116),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_56),
.B1(n_41),
.B2(n_36),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_75),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_36),
.B1(n_23),
.B2(n_37),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_37),
.B1(n_36),
.B2(n_42),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_108),
.B(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_83),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_120),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_61),
.B(n_35),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_34),
.B1(n_26),
.B2(n_31),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_40),
.B1(n_29),
.B2(n_27),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_87),
.B1(n_84),
.B2(n_31),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_123),
.B1(n_70),
.B2(n_66),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_0),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_94),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_40),
.B1(n_26),
.B2(n_30),
.Y(n_123)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_129),
.Y(n_163)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_138),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_137),
.B1(n_149),
.B2(n_153),
.Y(n_172)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_71),
.CI(n_33),
.CON(n_135),
.SN(n_135)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_135),
.B(n_141),
.Y(n_177)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_25),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_21),
.C(n_32),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_95),
.C(n_101),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_21),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_77),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_151),
.Y(n_169)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_170),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_165),
.B(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_110),
.B1(n_95),
.B2(n_120),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_171),
.B1(n_135),
.B2(n_154),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_119),
.B(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_96),
.C(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_173),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_126),
.B1(n_130),
.B2(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_118),
.Y(n_173)
);

NOR2x1p5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_123),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_123),
.B1(n_113),
.B2(n_117),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_111),
.C(n_76),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_123),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_183),
.B1(n_184),
.B2(n_199),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_179),
.B(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_198),
.Y(n_209)
);

AO21x2_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_130),
.B(n_97),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_154),
.B1(n_124),
.B2(n_141),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_186),
.B(n_167),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_146),
.C(n_125),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.C(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_124),
.B1(n_128),
.B2(n_117),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_189),
.A2(n_165),
.B1(n_128),
.B2(n_104),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_123),
.C(n_129),
.Y(n_192)
);

NOR4xp25_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_159),
.C(n_177),
.D(n_156),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

BUFx4f_ASAP7_75t_SL g194 ( 
.A(n_158),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_194),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_149),
.B1(n_127),
.B2(n_153),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_196),
.B(n_162),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_150),
.B(n_40),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_92),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_92),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_175),
.B1(n_171),
.B2(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_222),
.B1(n_199),
.B2(n_100),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_205),
.B(n_182),
.Y(n_232)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_210),
.Y(n_226)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_160),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_160),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_219),
.Y(n_230)
);

OR2x4_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_177),
.Y(n_217)
);

NOR4xp25_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_199),
.C(n_106),
.D(n_121),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_92),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_186),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_176),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_224),
.B(n_191),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_98),
.B1(n_136),
.B2(n_139),
.Y(n_222)
);

INVx2_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_223),
.Y(n_231)
);

NAND2x1_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_176),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_182),
.C(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_234),
.C(n_239),
.Y(n_252)
);

O2A1O1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_245),
.B(n_244),
.C(n_228),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_148),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_187),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_236),
.B(n_216),
.Y(n_260)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_199),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_144),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_243),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_194),
.C(n_164),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_201),
.C(n_200),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_208),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_200),
.B1(n_210),
.B2(n_223),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_218),
.B1(n_204),
.B2(n_224),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_157),
.B1(n_100),
.B2(n_111),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_157),
.B(n_121),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_221),
.B1(n_223),
.B2(n_217),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_256),
.B1(n_263),
.B2(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_216),
.B1(n_212),
.B2(n_207),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_220),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_267),
.C(n_231),
.Y(n_279)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_212),
.B1(n_222),
.B2(n_164),
.Y(n_263)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_248),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_76),
.C(n_111),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_229),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_113),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_233),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_65),
.B1(n_80),
.B2(n_66),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_225),
.B1(n_241),
.B2(n_249),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_82),
.B1(n_90),
.B2(n_73),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_239),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_285),
.C(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_281),
.B(n_287),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_283),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_253),
.B(n_234),
.CI(n_232),
.CON(n_283),
.SN(n_283)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_268),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_251),
.A2(n_243),
.B1(n_230),
.B2(n_246),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_269),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_266),
.B1(n_265),
.B2(n_270),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_259),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_257),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_283),
.C(n_275),
.Y(n_309)
);

HAxp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_264),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_256),
.Y(n_294)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_252),
.C(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_30),
.C(n_21),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_263),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_277),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_303),
.B(n_0),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_21),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_288),
.B1(n_73),
.B2(n_278),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_307),
.B(n_308),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_297),
.A2(n_274),
.B1(n_281),
.B2(n_283),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_312),
.C(n_313),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_82),
.B1(n_12),
.B2(n_2),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_319),
.C(n_30),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_77),
.C(n_67),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_67),
.C(n_32),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_10),
.B(n_18),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_9),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_306),
.B1(n_300),
.B2(n_292),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_315),
.A2(n_318),
.B1(n_10),
.B2(n_17),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_32),
.C(n_30),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_30),
.C(n_1),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_305),
.B(n_295),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_7),
.B(n_16),
.Y(n_338)
);

HAxp5_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_305),
.CON(n_322),
.SN(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_326),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_303),
.B(n_9),
.C(n_2),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_330),
.B(n_318),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_329),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_0),
.B(n_1),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_312),
.B(n_8),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_331),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_324),
.B(n_319),
.CI(n_313),
.CON(n_334),
.SN(n_334)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_334),
.B(n_340),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_322),
.A2(n_316),
.B(n_12),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_336),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_323),
.A2(n_7),
.B(n_17),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_339),
.B(n_3),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_342),
.B(n_344),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_325),
.B(n_328),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_325),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_4),
.B(n_5),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_337),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_349),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_5),
.C(n_6),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_341),
.C(n_12),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_347),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_352),
.B1(n_13),
.B2(n_15),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_6),
.C(n_15),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_16),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_18),
.B(n_353),
.Y(n_357)
);


endmodule