module fake_jpeg_29243_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_15),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_37),
.Y(n_62)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_25),
.B1(n_20),
.B2(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_61),
.B1(n_16),
.B2(n_18),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_69),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_36),
.B(n_27),
.C(n_18),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_33),
.B(n_19),
.C(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_24),
.B1(n_20),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_32),
.B1(n_23),
.B2(n_22),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_23),
.B1(n_22),
.B2(n_32),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_21),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_44),
.B1(n_38),
.B2(n_46),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_70),
.A2(n_106),
.B1(n_23),
.B2(n_36),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_88),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_33),
.B1(n_51),
.B2(n_31),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_77),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_56),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_39),
.C(n_33),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_92),
.C(n_24),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_41),
.B1(n_47),
.B2(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_98),
.B1(n_85),
.B2(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_85),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_94),
.Y(n_111)
);

OA22x2_ASAP7_75t_SL g82 ( 
.A1(n_67),
.A2(n_59),
.B1(n_55),
.B2(n_63),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_83),
.Y(n_110)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_29),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_48),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_16),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_107),
.B1(n_108),
.B2(n_16),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_96),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_35),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_52),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_35),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_121),
.C(n_136),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_118),
.B1(n_134),
.B2(n_137),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_117),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_68),
.B1(n_18),
.B2(n_36),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_49),
.C(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_75),
.B1(n_80),
.B2(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_82),
.B1(n_77),
.B2(n_78),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_34),
.C(n_28),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_76),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_140),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_15),
.B1(n_5),
.B2(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_73),
.B1(n_88),
.B2(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_86),
.B1(n_93),
.B2(n_71),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_131),
.B1(n_128),
.B2(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_86),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_102),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_27),
.B(n_96),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_125),
.B(n_124),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_74),
.B(n_95),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_135),
.B(n_133),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_89),
.B1(n_101),
.B2(n_91),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_159),
.B1(n_136),
.B2(n_110),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_84),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_7),
.B1(n_14),
.B2(n_12),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_10),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_148),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_155),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_156),
.C(n_112),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_172),
.C(n_176),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_173),
.B1(n_185),
.B2(n_139),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_140),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_121),
.C(n_109),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_180),
.B(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_178),
.B(n_190),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_133),
.B1(n_115),
.B2(n_125),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_146),
.B1(n_142),
.B2(n_141),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_135),
.B(n_119),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_119),
.B1(n_115),
.B2(n_110),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_110),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_1),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_1),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_6),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_192),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_172),
.B1(n_167),
.B2(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_165),
.B1(n_168),
.B2(n_177),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_211),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_203),
.A2(n_215),
.B(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_210),
.B1(n_167),
.B2(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_185),
.B1(n_186),
.B2(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_3),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_1),
.B(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_226),
.B1(n_228),
.B2(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_210),
.B1(n_199),
.B2(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_176),
.C(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_231),
.C(n_215),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_192),
.B1(n_182),
.B2(n_184),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_191),
.C(n_174),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_207),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_194),
.C(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_252),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_SL g241 ( 
.A(n_225),
.B(n_203),
.C(n_198),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_231),
.B(n_220),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_247),
.B1(n_248),
.B2(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_226),
.C(n_218),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_213),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_251),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_246),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_214),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_212),
.B1(n_206),
.B2(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_224),
.B1(n_218),
.B2(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_235),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_233),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_255),
.B(n_259),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_261),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_243),
.C(n_238),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_228),
.C(n_237),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_266),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_220),
.B(n_202),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_244),
.C(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_174),
.C(n_4),
.Y(n_270)
);

NAND2x1_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_8),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_12),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_259),
.C(n_256),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_254),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_266),
.B1(n_262),
.B2(n_257),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

HAxp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_265),
.CON(n_281),
.SN(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_268),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_264),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_289),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_276),
.B(n_271),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_284),
.B(n_279),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_285),
.C(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.C(n_280),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.B(n_285),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_283),
.B1(n_278),
.B2(n_8),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_8),
.B(n_9),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_12),
.B(n_1),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_2),
.C(n_283),
.Y(n_300)
);


endmodule