module fake_jpeg_19049_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_27),
.C(n_16),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_50),
.C(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_8),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_24),
.B(n_20),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_16),
.B1(n_31),
.B2(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_24),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_14),
.B(n_19),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_53),
.B(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_58),
.Y(n_82)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_37),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_60),
.B(n_68),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_20),
.B1(n_13),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_67),
.B1(n_51),
.B2(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_18),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_23),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_17),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_22),
.B(n_8),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_81),
.Y(n_87)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_80),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_57),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_43),
.Y(n_78)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_52),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_43),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_94),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_53),
.B(n_59),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_89),
.B(n_93),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_61),
.B(n_69),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_57),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_80),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_64),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_71),
.C(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_105),
.C(n_97),
.Y(n_108)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_106),
.B(n_98),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_79),
.C(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_58),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_109),
.C(n_112),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_92),
.C(n_87),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_78),
.A3(n_85),
.B1(n_42),
.B2(n_79),
.C(n_44),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_55),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_43),
.C(n_44),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_101),
.B(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_3),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_3),
.B(n_4),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_122),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_4),
.B(n_5),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_121),
.A2(n_10),
.B(n_12),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_10),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_5),
.B(n_49),
.C(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_12),
.Y(n_125)
);

AO221x1_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_5),
.B1(n_52),
.B2(n_49),
.C(n_117),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_49),
.Y(n_129)
);


endmodule