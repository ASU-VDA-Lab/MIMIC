module fake_jpeg_25376_n_199 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_49),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_42),
.B1(n_50),
.B2(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_30),
.C(n_22),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_51),
.C(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_12),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_18),
.B1(n_13),
.B2(n_20),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_18),
.B(n_13),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_12),
.B1(n_17),
.B2(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_66),
.B(n_67),
.C(n_70),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_27),
.B1(n_54),
.B2(n_52),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_73),
.B1(n_23),
.B2(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_17),
.B1(n_12),
.B2(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_72),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_20),
.B1(n_18),
.B2(n_13),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_37),
.B1(n_23),
.B2(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_40),
.C(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_30),
.C(n_25),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_73),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_42),
.B1(n_39),
.B2(n_25),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_91),
.B1(n_83),
.B2(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_15),
.B(n_21),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_19),
.B(n_1),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_30),
.C(n_22),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_14),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_113),
.B1(n_114),
.B2(n_0),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_58),
.B1(n_81),
.B2(n_77),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_111),
.B1(n_6),
.B2(n_2),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_106),
.B(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_108),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_88),
.B(n_74),
.C(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_57),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_116),
.B(n_0),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_56),
.B1(n_65),
.B2(n_63),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_39),
.B1(n_22),
.B2(n_15),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_16),
.B1(n_19),
.B2(n_14),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

XOR2x1_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_19),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_122),
.B1(n_95),
.B2(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_9),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_135),
.C(n_127),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_127),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_2),
.B(n_4),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_7),
.C(n_4),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_95),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_2),
.B(n_4),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_6),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_149),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_151),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_104),
.C(n_102),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_121),
.C(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_129),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_143),
.Y(n_165)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_123),
.B1(n_134),
.B2(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_159),
.B1(n_151),
.B2(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_112),
.B1(n_98),
.B2(n_119),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_98),
.B(n_131),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_94),
.C(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_135),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_171),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_144),
.B1(n_148),
.B2(n_108),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_139),
.C(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_165),
.C(n_166),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_140),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_156),
.B(n_162),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_156),
.B(n_160),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_185),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_171),
.B1(n_157),
.B2(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_173),
.B(n_177),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_190),
.B(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_158),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_195),
.A3(n_122),
.B1(n_159),
.B2(n_117),
.C1(n_130),
.C2(n_114),
.Y(n_197)
);

AO21x1_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_6),
.B(n_2),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_5),
.Y(n_199)
);


endmodule