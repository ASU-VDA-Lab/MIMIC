module fake_jpeg_8772_n_88 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_7),
.B(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_2),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_47),
.B(n_50),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_2),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_5),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_53),
.B(n_56),
.C(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_9),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_14),
.B1(n_40),
.B2(n_41),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_43),
.B(n_34),
.C(n_32),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_36),
.B1(n_27),
.B2(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_62),
.B1(n_49),
.B2(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_35),
.C(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_39),
.B1(n_43),
.B2(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_67),
.B(n_60),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_68),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_74),
.B(n_64),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_58),
.B1(n_51),
.B2(n_57),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_80),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_71),
.C(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_59),
.C(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_84),
.B(n_85),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_82),
.A2(n_55),
.B(n_37),
.C(n_64),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_69),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);


endmodule