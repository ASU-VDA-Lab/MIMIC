module fake_jpeg_12754_n_381 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_381);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_381;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_64),
.Y(n_113)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_69),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_78),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_20),
.B1(n_36),
.B2(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_111),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_64),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_22),
.C(n_33),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_33),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_23),
.B1(n_37),
.B2(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_102),
.B1(n_107),
.B2(n_117),
.Y(n_143)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_27),
.CON(n_97),
.SN(n_97)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_28),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_39),
.B1(n_42),
.B2(n_40),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_99),
.A2(n_116),
.B1(n_117),
.B2(n_123),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_57),
.A2(n_37),
.B1(n_31),
.B2(n_35),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_62),
.A2(n_35),
.B1(n_31),
.B2(n_18),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_71),
.B1(n_26),
.B2(n_59),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_60),
.B(n_20),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_50),
.A2(n_24),
.B1(n_42),
.B2(n_40),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_24),
.B1(n_42),
.B2(n_40),
.Y(n_117)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_53),
.A2(n_24),
.B1(n_42),
.B2(n_40),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_35),
.B1(n_26),
.B2(n_28),
.Y(n_142)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_77),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_2),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_54),
.B1(n_26),
.B2(n_35),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_136),
.A2(n_147),
.B1(n_158),
.B2(n_163),
.Y(n_192)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_140),
.B(n_151),
.Y(n_181)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_109),
.B1(n_115),
.B2(n_105),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_38),
.C(n_36),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_150),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_28),
.B1(n_97),
.B2(n_18),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_34),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_89),
.B(n_43),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_34),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_156),
.B(n_165),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_1),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_86),
.A2(n_43),
.B1(n_46),
.B2(n_75),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_161),
.Y(n_201)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_100),
.B(n_72),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_162),
.A2(n_121),
.B(n_118),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_98),
.A2(n_43),
.B1(n_46),
.B2(n_75),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_92),
.A2(n_72),
.B(n_60),
.C(n_13),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_12),
.B(n_11),
.C(n_124),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_43),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_43),
.B1(n_52),
.B2(n_41),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_41),
.B1(n_16),
.B2(n_14),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_95),
.B1(n_115),
.B2(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_168),
.B(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_93),
.B(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_172),
.A2(n_175),
.B1(n_180),
.B2(n_182),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_130),
.A2(n_93),
.B(n_95),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_153),
.B(n_152),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_149),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_103),
.B1(n_88),
.B2(n_90),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_103),
.B1(n_88),
.B2(n_90),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_124),
.B1(n_118),
.B2(n_122),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_183),
.A2(n_199),
.B1(n_207),
.B2(n_173),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_158),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_146),
.B(n_2),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_5),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_127),
.B1(n_139),
.B2(n_135),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_3),
.B(n_4),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_193),
.B(n_203),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_236),
.B1(n_183),
.B2(n_225),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_233),
.Y(n_246)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_138),
.B(n_129),
.C(n_144),
.D(n_136),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_211),
.A2(n_238),
.B(n_191),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_129),
.B1(n_168),
.B2(n_155),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_216),
.B1(n_236),
.B2(n_199),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_160),
.B1(n_131),
.B2(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_141),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_226),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_232),
.B(n_184),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_134),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_128),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_145),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_131),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_235),
.Y(n_263)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_133),
.C(n_154),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_133),
.B(n_149),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g235 ( 
.A1(n_182),
.A2(n_5),
.B1(n_180),
.B2(n_196),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_196),
.B1(n_177),
.B2(n_175),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_186),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_SL g240 ( 
.A(n_173),
.B(n_196),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_242),
.A2(n_243),
.B(n_245),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_260),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_203),
.B(n_201),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_207),
.B1(n_194),
.B2(n_197),
.Y(n_247)
);

OAI22x1_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_257),
.B1(n_237),
.B2(n_210),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_234),
.A2(n_216),
.B1(n_226),
.B2(n_230),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_211),
.B(n_238),
.Y(n_289)
);

INVx3_ASAP7_75t_SL g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_197),
.B1(n_188),
.B2(n_191),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_186),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_217),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_200),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_222),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_285),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_240),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_275),
.C(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_228),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_280),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_219),
.B1(n_232),
.B2(n_235),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_254),
.B1(n_264),
.B2(n_256),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_260),
.C(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_223),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_246),
.B(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_283),
.Y(n_310)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_252),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_241),
.B(n_248),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_290),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_200),
.B(n_206),
.Y(n_312)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_221),
.A3(n_231),
.B1(n_213),
.B2(n_237),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_195),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_281),
.A2(n_244),
.B(n_247),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_305),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_256),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_297),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_259),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_303),
.C(n_311),
.Y(n_328)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_289),
.A2(n_254),
.B(n_251),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_251),
.B(n_262),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_270),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_289),
.A2(n_262),
.B1(n_213),
.B2(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_308),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_195),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_291),
.Y(n_329)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_316),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_295),
.B1(n_311),
.B2(n_301),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_318),
.B(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_300),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_321),
.B1(n_322),
.B2(n_325),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_304),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_293),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_272),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_301),
.B1(n_312),
.B2(n_305),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_298),
.C(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_339),
.C(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_297),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_334),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_303),
.CI(n_309),
.CON(n_335),
.SN(n_335)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_321),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_342),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_296),
.C(n_307),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_294),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_326),
.A2(n_284),
.B1(n_295),
.B2(n_278),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_329),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_351),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_339),
.A2(n_316),
.B(n_322),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_345),
.A2(n_347),
.B(n_352),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_325),
.C(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_350),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_317),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_315),
.B(n_313),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_292),
.C(n_282),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_353),
.B(n_338),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_337),
.C(n_338),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_358),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_341),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_348),
.B(n_343),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_360),
.B(n_362),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_285),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_346),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_349),
.C(n_353),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_330),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_365),
.A2(n_368),
.B(n_370),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_359),
.B(n_351),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_366),
.B(n_357),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_361),
.Y(n_374)
);

OAI21x1_ASAP7_75t_SL g370 ( 
.A1(n_356),
.A2(n_269),
.B(n_335),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_372),
.A2(n_373),
.B(n_374),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

A2O1A1O1Ixp25_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_367),
.B(n_369),
.C(n_349),
.D(n_290),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_375),
.B(n_286),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_376),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_379),
.B(n_277),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_277),
.B(n_206),
.Y(n_381)
);


endmodule