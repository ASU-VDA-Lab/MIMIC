module fake_jpeg_22116_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_6),
.B(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_37),
.Y(n_74)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_72),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_77),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_70),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_25),
.B1(n_36),
.B2(n_27),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_92),
.B1(n_17),
.B2(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_26),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_97),
.B(n_26),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_39),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_93),
.B1(n_63),
.B2(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_49),
.B(n_46),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_27),
.B1(n_60),
.B2(n_94),
.Y(n_103)
);

OR2x4_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_26),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_38),
.B1(n_41),
.B2(n_22),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_112),
.B1(n_121),
.B2(n_69),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_97),
.A2(n_38),
.B(n_41),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_103),
.B1(n_122),
.B2(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_109),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_48),
.B1(n_37),
.B2(n_24),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_48),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_47),
.C(n_24),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_90),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_94),
.B1(n_24),
.B2(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_84),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_130),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_8),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_20),
.Y(n_185)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_133),
.Y(n_173)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_138),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_37),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_150),
.B(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_145),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_37),
.B1(n_98),
.B2(n_83),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_154),
.B1(n_145),
.B2(n_146),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_67),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_0),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_85),
.B1(n_21),
.B2(n_17),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_156),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_166),
.B(n_187),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_99),
.B1(n_123),
.B2(n_114),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_123),
.B1(n_108),
.B2(n_125),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_136),
.B1(n_148),
.B2(n_134),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_29),
.B(n_17),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_171),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_181),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_142),
.A2(n_108),
.B1(n_104),
.B2(n_119),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_120),
.B1(n_132),
.B2(n_133),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_126),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_141),
.C(n_140),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_179),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_155),
.A2(n_107),
.B1(n_138),
.B2(n_153),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_150),
.B(n_131),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_129),
.B1(n_21),
.B2(n_104),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_28),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_143),
.C(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_129),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_167),
.C(n_170),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_204),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_210),
.B(n_218),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_126),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_201),
.B(n_203),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_132),
.B1(n_157),
.B2(n_98),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_127),
.C(n_75),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_208),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_29),
.B(n_33),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_220),
.B1(n_177),
.B2(n_163),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_70),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_43),
.C(n_40),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_34),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_169),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_174),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_31),
.B(n_30),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_28),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_219),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_199),
.Y(n_252)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_183),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_R g235 ( 
.A(n_199),
.B(n_166),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_209),
.B1(n_193),
.B2(n_195),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_206),
.A2(n_185),
.B(n_158),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_18),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_18),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_246),
.Y(n_255)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_196),
.A2(n_34),
.A3(n_32),
.B1(n_18),
.B2(n_28),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_34),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_189),
.C(n_216),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_249),
.C(n_253),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_228),
.C(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_205),
.C(n_210),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_200),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_209),
.B1(n_213),
.B2(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_217),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_221),
.C(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_28),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_28),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_32),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_13),
.B(n_16),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_226),
.B1(n_43),
.B2(n_40),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_234),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_227),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_274),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_235),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_226),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_277),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_225),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_241),
.C(n_245),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_251),
.A2(n_239),
.B1(n_242),
.B2(n_236),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_251),
.B1(n_253),
.B2(n_259),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_287),
.A2(n_297),
.B1(n_23),
.B2(n_30),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_247),
.B(n_256),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_289),
.B(n_1),
.Y(n_308)
);

BUFx12f_ASAP7_75t_SL g289 ( 
.A(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_293),
.Y(n_307)
);

XOR2x1_ASAP7_75t_SL g291 ( 
.A(n_274),
.B(n_261),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_275),
.C(n_285),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_262),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_270),
.A2(n_230),
.B1(n_250),
.B2(n_243),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_276),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_230),
.B1(n_223),
.B2(n_240),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_279),
.C(n_285),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_279),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_309),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.C(n_310),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_275),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_305),
.A2(n_8),
.B(n_15),
.C(n_3),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_282),
.B1(n_272),
.B2(n_31),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_292),
.B1(n_304),
.B2(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_32),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_291),
.B(n_299),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_10),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_313),
.B(n_16),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_8),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_303),
.C(n_305),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_320),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_23),
.C(n_10),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_11),
.C(n_15),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_316),
.B(n_10),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_11),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_314),
.A2(n_7),
.B(n_14),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_325),
.A2(n_326),
.B(n_327),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_7),
.B(n_12),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_331),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_321),
.B(n_313),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_319),
.B(n_7),
.C(n_4),
.D(n_6),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_329),
.B1(n_330),
.B2(n_12),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_333),
.B(n_12),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_14),
.C(n_1),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_1),
.B(n_2),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_2),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_339),
.B(n_2),
.Y(n_340)
);


endmodule