module real_jpeg_9043_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_20),
.B1(n_21),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_3),
.A2(n_55),
.B(n_57),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_3),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_3),
.B(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_3),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_22),
.B1(n_29),
.B2(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_46),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_36),
.B(n_38),
.C(n_39),
.D(n_44),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_43),
.Y(n_68)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_20),
.B(n_24),
.C(n_78),
.D(n_79),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_10),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_58),
.B(n_71),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_74),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_73),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_62),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_62),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_50),
.B2(n_61),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B1(n_32),
.B2(n_34),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_19),
.A2(n_34),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_20),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_25),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_25),
.B(n_31),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_27),
.A2(n_29),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_59),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_31),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_34),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_59),
.A2(n_91),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_99),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.C(n_69),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_70),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_87),
.B(n_108),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_80),
.B1(n_81),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_96),
.B(n_107),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_94),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_102),
.B(n_106),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);


endmodule