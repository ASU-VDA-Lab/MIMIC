module real_aes_475_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_0), .B(n_152), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_1), .A2(n_161), .B(n_166), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_2), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_3), .B(n_152), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_4), .B(n_168), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_5), .B(n_168), .Y(n_206) );
INVx1_ASAP7_75t_L g159 ( .A(n_6), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_7), .B(n_168), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_8), .Y(n_109) );
NAND2xp33_ASAP7_75t_L g195 ( .A(n_9), .B(n_170), .Y(n_195) );
AND2x2_ASAP7_75t_L g505 ( .A(n_10), .B(n_189), .Y(n_505) );
AND2x2_ASAP7_75t_L g513 ( .A(n_11), .B(n_146), .Y(n_513) );
INVx2_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
AOI221x1_ASAP7_75t_L g241 ( .A1(n_13), .A2(n_24), .B1(n_152), .B2(n_161), .C(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_14), .B(n_168), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_16), .B(n_152), .Y(n_191) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_17), .A2(n_189), .B(n_190), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_18), .B(n_172), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_19), .B(n_168), .Y(n_182) );
AO21x1_ASAP7_75t_L g201 ( .A1(n_20), .A2(n_152), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_21), .B(n_152), .Y(n_486) );
INVx1_ASAP7_75t_L g106 ( .A(n_22), .Y(n_106) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_23), .A2(n_90), .B1(n_152), .B2(n_521), .Y(n_520) );
NAND2x1_ASAP7_75t_L g214 ( .A(n_25), .B(n_168), .Y(n_214) );
NAND2x1_ASAP7_75t_L g233 ( .A(n_26), .B(n_170), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g781 ( .A1(n_27), .A2(n_63), .B1(n_782), .B2(n_783), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_27), .Y(n_782) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_28), .A2(n_87), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g174 ( .A(n_28), .B(n_87), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_29), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_30), .B(n_168), .Y(n_194) );
AO21x2_ASAP7_75t_L g460 ( .A1(n_31), .A2(n_146), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_32), .B(n_170), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_33), .A2(n_161), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_34), .B(n_168), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_35), .A2(n_161), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g158 ( .A(n_36), .B(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g162 ( .A(n_36), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g529 ( .A(n_36), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_37), .B(n_108), .C(n_110), .Y(n_107) );
OR2x6_ASAP7_75t_L g124 ( .A(n_37), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_38), .B(n_152), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_39), .B(n_152), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_40), .B(n_168), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_41), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_42), .B(n_170), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_43), .B(n_152), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_44), .A2(n_161), .B(n_509), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_45), .A2(n_161), .B(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_46), .B(n_170), .Y(n_552) );
INVxp33_ASAP7_75t_L g788 ( .A(n_47), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_48), .A2(n_52), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_48), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_49), .B(n_170), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_50), .B(n_152), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_51), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_52), .Y(n_130) );
INVx1_ASAP7_75t_L g155 ( .A(n_53), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_53), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_54), .B(n_168), .Y(n_511) );
AND2x2_ASAP7_75t_L g477 ( .A(n_55), .B(n_172), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_56), .B(n_170), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_57), .B(n_168), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_58), .B(n_170), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_59), .A2(n_161), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_60), .B(n_152), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_61), .B(n_152), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_62), .A2(n_161), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_63), .Y(n_783) );
AO21x1_ASAP7_75t_L g203 ( .A1(n_64), .A2(n_161), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g492 ( .A(n_65), .B(n_173), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_66), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_67), .B(n_170), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_68), .B(n_152), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_69), .B(n_170), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_70), .A2(n_95), .B1(n_161), .B2(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g226 ( .A(n_71), .B(n_173), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_72), .B(n_168), .Y(n_489) );
INVx1_ASAP7_75t_L g157 ( .A(n_73), .Y(n_157) );
INVx1_ASAP7_75t_L g163 ( .A(n_73), .Y(n_163) );
AND2x2_ASAP7_75t_L g237 ( .A(n_74), .B(n_146), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_75), .B(n_170), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_76), .A2(n_161), .B(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_77), .A2(n_161), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_78), .A2(n_161), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g474 ( .A(n_79), .B(n_173), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_80), .B(n_172), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_81), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
AND2x2_ASAP7_75t_L g145 ( .A(n_82), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_83), .B(n_152), .Y(n_184) );
AND2x2_ASAP7_75t_L g553 ( .A(n_84), .B(n_189), .Y(n_553) );
AND2x2_ASAP7_75t_L g202 ( .A(n_85), .B(n_178), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_86), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_170), .Y(n_183) );
AND2x2_ASAP7_75t_L g218 ( .A(n_89), .B(n_146), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_91), .B(n_168), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_92), .A2(n_161), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_93), .B(n_170), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_94), .A2(n_161), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_96), .B(n_168), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_97), .B(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g491 ( .A(n_98), .Y(n_491) );
BUFx2_ASAP7_75t_L g115 ( .A(n_99), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_100), .A2(n_161), .B(n_193), .Y(n_192) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_111), .B(n_787), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g790 ( .A(n_103), .Y(n_790) );
INVx3_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_107), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_106), .B(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_110), .B(n_123), .Y(n_122) );
OR2x6_ASAP7_75t_SL g136 ( .A(n_110), .B(n_123), .Y(n_136) );
AND2x6_ASAP7_75t_SL g766 ( .A(n_110), .B(n_124), .Y(n_766) );
OR2x2_ASAP7_75t_L g775 ( .A(n_110), .B(n_124), .Y(n_775) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_128), .B(n_776), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_115), .Y(n_777) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_117), .A2(n_779), .B(n_784), .Y(n_778) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_127), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g786 ( .A(n_122), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_767), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_129), .A2(n_768), .B(n_772), .Y(n_767) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B1(n_454), .B2(n_763), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g771 ( .A(n_135), .Y(n_771) );
CKINVDCx11_ASAP7_75t_R g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g770 ( .A(n_137), .Y(n_770) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_363), .Y(n_137) );
NOR4xp25_ASAP7_75t_L g138 ( .A(n_139), .B(n_281), .C(n_307), .D(n_347), .Y(n_138) );
OAI211xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_196), .B(n_227), .C(n_267), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_175), .Y(n_141) );
AND2x2_ASAP7_75t_L g434 ( .A(n_142), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_143), .B(n_175), .Y(n_301) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g228 ( .A(n_144), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_144), .B(n_254), .Y(n_253) );
INVx5_ASAP7_75t_L g287 ( .A(n_144), .Y(n_287) );
NOR2x1_ASAP7_75t_SL g329 ( .A(n_144), .B(n_176), .Y(n_329) );
AND2x2_ASAP7_75t_L g385 ( .A(n_144), .B(n_188), .Y(n_385) );
OR2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_150), .Y(n_144) );
INVx3_ASAP7_75t_L g217 ( .A(n_146), .Y(n_217) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_147), .A2(n_507), .B(n_513), .Y(n_506) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_149), .B(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g178 ( .A(n_149), .B(n_174), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_160), .B(n_172), .Y(n_150) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_158), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
AND2x6_ASAP7_75t_L g170 ( .A(n_154), .B(n_163), .Y(n_170) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g168 ( .A(n_156), .B(n_165), .Y(n_168) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx5_ASAP7_75t_L g171 ( .A(n_158), .Y(n_171) );
AND2x2_ASAP7_75t_L g164 ( .A(n_159), .B(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_159), .Y(n_524) );
AND2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_164), .Y(n_161) );
BUFx3_ASAP7_75t_L g525 ( .A(n_162), .Y(n_525) );
INVx2_ASAP7_75t_L g531 ( .A(n_163), .Y(n_531) );
AND2x4_ASAP7_75t_L g527 ( .A(n_164), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g523 ( .A(n_165), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_171), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_170), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_171), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_171), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_171), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_171), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_171), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_171), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_171), .A2(n_465), .B(n_466), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_171), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_171), .A2(n_482), .B(n_483), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_171), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_171), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_171), .A2(n_510), .B(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_171), .A2(n_551), .B(n_552), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_172), .Y(n_236) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_172), .A2(n_241), .B(n_245), .Y(n_240) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_172), .A2(n_241), .B(n_245), .Y(n_280) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_172), .A2(n_520), .B(n_526), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_172), .A2(n_548), .B(n_549), .Y(n_547) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_187), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_176), .B(n_188), .Y(n_257) );
AND2x2_ASAP7_75t_L g318 ( .A(n_176), .B(n_287), .Y(n_318) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B(n_185), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_177), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_177), .A2(n_179), .B(n_185), .Y(n_271) );
INVx1_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_178), .A2(n_191), .B(n_192), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_178), .B(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_178), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_178), .A2(n_479), .B(n_480), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_184), .Y(n_179) );
AND2x2_ASAP7_75t_L g330 ( .A(n_187), .B(n_254), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_187), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g374 ( .A(n_187), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g407 ( .A(n_187), .B(n_228), .Y(n_407) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g251 ( .A(n_188), .Y(n_251) );
AND2x2_ASAP7_75t_L g284 ( .A(n_188), .B(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
OR2x2_ASAP7_75t_L g395 ( .A(n_188), .B(n_254), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_189), .A2(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
AOI211x1_ASAP7_75t_SL g324 ( .A1(n_198), .A2(n_316), .B(n_325), .C(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_198), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_198), .B(n_367), .Y(n_414) );
BUFx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
OAI21x1_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_207), .Y(n_200) );
INVx1_ASAP7_75t_L g208 ( .A(n_202), .Y(n_208) );
AOI322xp5_ASAP7_75t_L g227 ( .A1(n_209), .A2(n_228), .A3(n_238), .B1(n_246), .B2(n_249), .C1(n_255), .C2(n_258), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_209), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
INVx2_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
INVxp67_ASAP7_75t_L g304 ( .A(n_210), .Y(n_304) );
BUFx3_ASAP7_75t_L g368 ( .A(n_210), .Y(n_368) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_210) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_217), .A2(n_220), .B(n_226), .Y(n_219) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_217), .A2(n_220), .B(n_226), .Y(n_266) );
AO21x1_ASAP7_75t_SL g467 ( .A1(n_217), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_217), .A2(n_468), .B(n_474), .Y(n_543) );
INVx2_ASAP7_75t_L g277 ( .A(n_219), .Y(n_277) );
AND2x2_ASAP7_75t_L g326 ( .A(n_219), .B(n_240), .Y(n_326) );
AND2x2_ASAP7_75t_L g370 ( .A(n_219), .B(n_279), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_221), .B(n_225), .Y(n_220) );
AND2x2_ASAP7_75t_L g255 ( .A(n_228), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_228), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_228), .B(n_284), .Y(n_449) );
INVx4_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
AND2x2_ASAP7_75t_L g286 ( .A(n_229), .B(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_229), .Y(n_339) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_236), .B(n_237), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_235), .Y(n_230) );
AOI21x1_ASAP7_75t_L g498 ( .A1(n_236), .A2(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_238), .B(n_323), .Y(n_348) );
INVx1_ASAP7_75t_SL g387 ( .A(n_238), .Y(n_387) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x4_ASAP7_75t_L g278 ( .A(n_239), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_239), .B(n_277), .Y(n_346) );
AND2x2_ASAP7_75t_L g398 ( .A(n_239), .B(n_248), .Y(n_398) );
OR2x2_ASAP7_75t_L g422 ( .A(n_239), .B(n_240), .Y(n_422) );
AND2x2_ASAP7_75t_L g246 ( .A(n_240), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g296 ( .A(n_240), .B(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_SL g352 ( .A(n_240), .B(n_264), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_246), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
BUFx2_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
AND2x4_ASAP7_75t_SL g351 ( .A(n_248), .B(n_265), .Y(n_351) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_252), .Y(n_249) );
OR2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_253), .Y(n_299) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g268 ( .A(n_251), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g416 ( .A(n_251), .B(n_329), .Y(n_416) );
AND2x2_ASAP7_75t_L g432 ( .A(n_251), .B(n_286), .Y(n_432) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI311xp33_ASAP7_75t_L g402 ( .A1(n_253), .A2(n_341), .A3(n_403), .B(n_405), .C(n_412), .Y(n_402) );
AND2x4_ASAP7_75t_L g269 ( .A(n_254), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_254), .B(n_287), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_254), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g386 ( .A(n_254), .B(n_373), .Y(n_386) );
AND2x2_ASAP7_75t_L g272 ( .A(n_256), .B(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_257), .Y(n_290) );
OR2x2_ASAP7_75t_L g379 ( .A(n_257), .B(n_343), .Y(n_379) );
INVx1_ASAP7_75t_L g435 ( .A(n_257), .Y(n_435) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g344 ( .A(n_261), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g358 ( .A(n_261), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g433 ( .A(n_261), .B(n_306), .Y(n_433) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g276 ( .A(n_262), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g295 ( .A(n_262), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g357 ( .A(n_263), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_263), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g306 ( .A(n_264), .B(n_277), .Y(n_306) );
AND2x4_ASAP7_75t_L g359 ( .A(n_264), .B(n_266), .Y(n_359) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp33_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_272), .B(n_274), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_268), .A2(n_354), .B1(n_358), .B2(n_360), .Y(n_353) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_269), .B(n_287), .Y(n_313) );
INVx2_ASAP7_75t_L g375 ( .A(n_269), .Y(n_375) );
AND2x2_ASAP7_75t_L g389 ( .A(n_269), .B(n_385), .Y(n_389) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g285 ( .A(n_271), .Y(n_285) );
INVx1_ASAP7_75t_L g338 ( .A(n_271), .Y(n_338) );
INVx1_ASAP7_75t_L g289 ( .A(n_273), .Y(n_289) );
AND3x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_318), .C(n_319), .Y(n_317) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g381 ( .A(n_276), .Y(n_381) );
AND2x2_ASAP7_75t_L g309 ( .A(n_278), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g380 ( .A(n_278), .B(n_381), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_278), .A2(n_392), .B1(n_396), .B2(n_399), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_278), .B(n_426), .Y(n_430) );
BUFx2_ASAP7_75t_L g321 ( .A(n_279), .Y(n_321) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_280), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_291), .B1(n_293), .B2(n_294), .C(n_297), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_283), .B(n_288), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g373 ( .A(n_285), .Y(n_373) );
INVx2_ASAP7_75t_SL g362 ( .A(n_286), .Y(n_362) );
AND2x2_ASAP7_75t_L g444 ( .A(n_286), .B(n_311), .Y(n_444) );
INVx4_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
INVx1_ASAP7_75t_L g293 ( .A(n_288), .Y(n_293) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x4_ASAP7_75t_L g404 ( .A(n_292), .B(n_359), .Y(n_404) );
INVx1_ASAP7_75t_SL g443 ( .A(n_292), .Y(n_443) );
AND2x2_ASAP7_75t_L g448 ( .A(n_292), .B(n_351), .Y(n_448) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g390 ( .A(n_296), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g323 ( .A(n_304), .Y(n_323) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g320 ( .A(n_306), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g410 ( .A(n_306), .B(n_411), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_312), .B(n_314), .C(n_331), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_310), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_311), .B(n_326), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_311), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g436 ( .A(n_311), .B(n_359), .Y(n_436) );
OAI221xp5_ASAP7_75t_SL g347 ( .A1(n_312), .A2(n_336), .B1(n_348), .B2(n_349), .C(n_353), .Y(n_347) );
INVx3_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g418 ( .A(n_313), .B(n_319), .Y(n_418) );
OAI32xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_320), .A3(n_322), .B1(n_324), .B2(n_328), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_318), .Y(n_408) );
INVx2_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_319), .A2(n_371), .B(n_451), .C(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
OR2x2_ASAP7_75t_L g452 ( .A(n_321), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_325), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g413 ( .A(n_328), .Y(n_413) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g394 ( .A(n_329), .Y(n_394) );
OAI21xp33_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_340), .B(n_344), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
OR2x2_ASAP7_75t_L g371 ( .A(n_334), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_335), .B(n_338), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_337), .A2(n_369), .B1(n_438), .B2(n_441), .C(n_445), .Y(n_437) );
INVx2_ASAP7_75t_L g440 ( .A(n_337), .Y(n_440) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g361 ( .A(n_341), .B(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g428 ( .A(n_341), .B(n_386), .Y(n_428) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g426 ( .A(n_351), .Y(n_426) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_359), .B(n_389), .Y(n_446) );
INVx2_ASAP7_75t_L g453 ( .A(n_359), .Y(n_453) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_361), .A2(n_424), .B1(n_427), .B2(n_429), .C(n_431), .Y(n_423) );
AND5x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_402), .C(n_417), .D(n_437), .E(n_447), .Y(n_363) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_382), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .B1(n_374), .B2(n_376), .C(n_377), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_387), .B1(n_388), .B2(n_390), .C(n_391), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_387), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
OR2x2_ASAP7_75t_L g400 ( .A(n_395), .B(n_401), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_423), .Y(n_417) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_434), .B2(n_436), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_433), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g451 ( .A(n_444), .Y(n_451) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx4_ASAP7_75t_L g769 ( .A(n_454), .Y(n_769) );
OAI22xp5_ASAP7_75t_SL g779 ( .A1(n_454), .A2(n_769), .B1(n_780), .B2(n_781), .Y(n_779) );
AND3x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_641), .C(n_737), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_583), .C(n_610), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_493), .B(n_532), .C(n_556), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_475), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_458), .A2(n_534), .B(n_538), .C(n_544), .Y(n_533) );
OR2x2_ASAP7_75t_L g656 ( .A(n_458), .B(n_593), .Y(n_656) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g623 ( .A(n_459), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_459), .B(n_594), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_459), .B(n_739), .Y(n_754) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
AND2x2_ASAP7_75t_L g540 ( .A(n_460), .B(n_476), .Y(n_540) );
INVx1_ASAP7_75t_L g560 ( .A(n_460), .Y(n_560) );
OR2x2_ASAP7_75t_L g575 ( .A(n_460), .B(n_484), .Y(n_575) );
INVx2_ASAP7_75t_L g581 ( .A(n_460), .Y(n_581) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_460), .Y(n_636) );
INVx1_ASAP7_75t_L g713 ( .A(n_460), .Y(n_713) );
NOR2x1_ASAP7_75t_SL g562 ( .A(n_467), .B(n_484), .Y(n_562) );
AND2x2_ASAP7_75t_L g592 ( .A(n_467), .B(n_581), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
OR2x2_ASAP7_75t_L g586 ( .A(n_475), .B(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_475), .B(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g714 ( .A(n_475), .Y(n_714) );
NAND2x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_484), .Y(n_475) );
OR2x2_ASAP7_75t_SL g574 ( .A(n_476), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g578 ( .A(n_476), .Y(n_578) );
INVx4_ASAP7_75t_L g594 ( .A(n_476), .Y(n_594) );
OR2x2_ASAP7_75t_L g609 ( .A(n_476), .B(n_542), .Y(n_609) );
AND2x2_ASAP7_75t_L g648 ( .A(n_476), .B(n_562), .Y(n_648) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_476), .Y(n_660) );
OR2x6_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g541 ( .A(n_484), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g593 ( .A(n_484), .B(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g608 ( .A(n_484), .Y(n_608) );
AND2x2_ASAP7_75t_L g624 ( .A(n_484), .B(n_594), .Y(n_624) );
AND2x2_ASAP7_75t_L g637 ( .A(n_484), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g669 ( .A(n_484), .B(n_581), .Y(n_669) );
INVx2_ASAP7_75t_SL g739 ( .A(n_484), .Y(n_739) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2xp67_ASAP7_75t_L g494 ( .A(n_495), .B(n_514), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_495), .A2(n_611), .B(n_615), .C(n_631), .Y(n_610) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g706 ( .A(n_496), .B(n_545), .Y(n_706) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx2_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
AND2x4_ASAP7_75t_SL g566 ( .A(n_497), .B(n_546), .Y(n_566) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_497), .Y(n_570) );
AND2x2_ASAP7_75t_L g628 ( .A(n_497), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g702 ( .A(n_497), .Y(n_702) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_498), .Y(n_604) );
AND2x2_ASAP7_75t_L g647 ( .A(n_498), .B(n_506), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_504), .Y(n_499) );
INVx2_ASAP7_75t_L g537 ( .A(n_506), .Y(n_537) );
AND2x2_ASAP7_75t_L g597 ( .A(n_506), .B(n_546), .Y(n_597) );
INVx2_ASAP7_75t_L g629 ( .A(n_506), .Y(n_629) );
OR2x2_ASAP7_75t_L g652 ( .A(n_506), .B(n_517), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_514), .B(n_569), .Y(n_676) );
AND2x2_ASAP7_75t_L g710 ( .A(n_514), .B(n_646), .Y(n_710) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI31xp33_ASAP7_75t_SL g631 ( .A1(n_515), .A2(n_612), .A3(n_632), .B(n_639), .Y(n_631) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_516), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g582 ( .A(n_517), .B(n_545), .Y(n_582) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x4_ASAP7_75t_L g572 ( .A(n_518), .B(n_519), .Y(n_572) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_525), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
NOR2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g717 ( .A(n_535), .Y(n_717) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_537), .B(n_546), .Y(n_599) );
AND2x2_ASAP7_75t_L g640 ( .A(n_537), .B(n_555), .Y(n_640) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AND2x2_ASAP7_75t_L g620 ( .A(n_541), .B(n_578), .Y(n_620) );
AND2x2_ASAP7_75t_L g579 ( .A(n_542), .B(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_542), .Y(n_588) );
INVx2_ASAP7_75t_L g638 ( .A(n_542), .Y(n_638) );
AND2x2_ASAP7_75t_L g728 ( .A(n_542), .B(n_713), .Y(n_728) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g734 ( .A(n_544), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_545), .B(n_554), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_545), .B(n_604), .Y(n_673) );
AND2x2_ASAP7_75t_L g721 ( .A(n_545), .B(n_647), .Y(n_721) );
INVx4_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g630 ( .A(n_546), .B(n_602), .Y(n_630) );
AND2x2_ASAP7_75t_L g639 ( .A(n_546), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g651 ( .A(n_546), .Y(n_651) );
BUFx2_ASAP7_75t_L g667 ( .A(n_546), .Y(n_667) );
AND2x4_ASAP7_75t_L g701 ( .A(n_546), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g746 ( .A(n_546), .B(n_647), .Y(n_746) );
OR2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_553), .Y(n_546) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AOI222xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_563), .B1(n_567), .B2(n_573), .C1(n_576), .C2(n_582), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_558), .A2(n_622), .B1(n_625), .B2(n_630), .Y(n_621) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g605 ( .A(n_559), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_SL g619 ( .A(n_559), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_559), .B(n_624), .Y(n_757) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g718 ( .A(n_560), .B(n_624), .Y(n_718) );
OR2x2_ASAP7_75t_L g695 ( .A(n_561), .B(n_577), .Y(n_695) );
OR2x2_ASAP7_75t_L g703 ( .A(n_561), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g687 ( .A(n_562), .B(n_580), .Y(n_687) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
OR2x2_ASAP7_75t_L g595 ( .A(n_565), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g745 ( .A(n_565), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g696 ( .A(n_566), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_566), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g731 ( .A(n_566), .Y(n_731) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g716 ( .A(n_569), .Y(n_716) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g618 ( .A(n_570), .B(n_597), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_571), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g617 ( .A(n_571), .Y(n_617) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_571), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g720 ( .A(n_571), .B(n_592), .Y(n_720) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g654 ( .A(n_572), .B(n_640), .Y(n_654) );
AND2x2_ASAP7_75t_L g697 ( .A(n_572), .B(n_629), .Y(n_697) );
AND2x4_ASAP7_75t_L g612 ( .A(n_573), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g753 ( .A(n_575), .B(n_609), .Y(n_753) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_577), .B(n_592), .Y(n_736) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_578), .B(n_592), .Y(n_658) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_578), .A2(n_619), .B(n_720), .C(n_721), .Y(n_719) );
AND2x2_ASAP7_75t_L g750 ( .A(n_578), .B(n_728), .Y(n_750) );
INVx1_ASAP7_75t_L g661 ( .A(n_579), .Y(n_661) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_582), .B(n_646), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_595), .B(n_598), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_586), .A2(n_739), .B1(n_740), .B2(n_742), .Y(n_738) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g614 ( .A(n_588), .Y(n_614) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g635 ( .A(n_594), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g686 ( .A(n_594), .Y(n_686) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_605), .Y(n_598) );
INVx1_ASAP7_75t_L g677 ( .A(n_599), .Y(n_677) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B(n_621), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
OR2x2_ASAP7_75t_L g662 ( .A(n_617), .B(n_663), .Y(n_662) );
OR2x2_ASAP7_75t_L g699 ( .A(n_617), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_617), .B(n_647), .Y(n_735) );
INVx1_ASAP7_75t_L g755 ( .A(n_618), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_620), .A2(n_723), .B1(n_726), .B2(n_729), .C(n_732), .Y(n_722) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI321xp33_ASAP7_75t_L g743 ( .A1(n_625), .A2(n_660), .A3(n_744), .B1(n_747), .B2(n_749), .C(n_751), .Y(n_743) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g684 ( .A(n_629), .Y(n_684) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g678 ( .A(n_634), .Y(n_678) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g704 ( .A(n_635), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_637), .A2(n_665), .B1(n_669), .B2(n_670), .C(n_675), .Y(n_664) );
INVxp67_ASAP7_75t_L g693 ( .A(n_638), .Y(n_693) );
INVx1_ASAP7_75t_L g663 ( .A(n_640), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g641 ( .A(n_642), .B(n_688), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_664), .C(n_679), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B1(n_649), .B2(n_655), .C(n_657), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g762 ( .A(n_647), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_653), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_651), .B(n_697), .Y(n_742) );
INVx2_ASAP7_75t_SL g674 ( .A(n_652), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_653), .A2(n_658), .B1(n_659), .B2(n_662), .Y(n_657) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_661), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_662), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g668 ( .A(n_663), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g707 ( .A1(n_665), .A2(n_708), .B1(n_710), .B2(n_711), .C1(n_715), .C2(n_718), .Y(n_707) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_666), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g741 ( .A(n_666), .B(n_720), .Y(n_741) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_674), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_674), .B(n_734), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_678), .Y(n_675) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_685), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_685), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND4xp25_ASAP7_75t_SL g688 ( .A(n_689), .B(n_707), .C(n_719), .D(n_722), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_694), .B(n_696), .C(n_698), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_695), .A2(n_699), .B1(n_703), .B2(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g725 ( .A(n_697), .Y(n_725) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_714), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_731), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B(n_736), .Y(n_732) );
NOR4xp25_ASAP7_75t_L g737 ( .A(n_738), .B(n_743), .C(n_756), .D(n_758), .Y(n_737) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx4_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx3_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
OAI22x1_ASAP7_75t_L g768 ( .A1(n_765), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
endmodule