module real_aes_6723_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g279 ( .A(n_0), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_1), .A2(n_194), .B1(n_195), .B2(n_199), .Y(n_193) );
INVx1_ASAP7_75t_L g199 ( .A(n_1), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_2), .Y(n_90) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_3), .A2(n_31), .B1(n_234), .B2(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_4), .B(n_259), .Y(n_268) );
INVx1_ASAP7_75t_L g215 ( .A(n_5), .Y(n_215) );
AND2x6_ASAP7_75t_L g252 ( .A(n_5), .B(n_213), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_5), .B(n_536), .Y(n_535) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_6), .A2(n_26), .B1(n_97), .B2(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g230 ( .A(n_7), .Y(n_230) );
INVx1_ASAP7_75t_L g272 ( .A(n_8), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_9), .B(n_238), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_10), .B(n_226), .Y(n_343) );
AO32x2_ASAP7_75t_L g285 ( .A1(n_11), .A2(n_225), .A3(n_251), .B1(n_259), .B2(n_286), .Y(n_285) );
XOR2xp5_ASAP7_75t_L g544 ( .A(n_12), .B(n_86), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_13), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_13), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_13), .B(n_234), .Y(n_311) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_14), .A2(n_56), .B1(n_189), .B2(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_14), .Y(n_190) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_15), .A2(n_28), .B1(n_97), .B2(n_101), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_16), .B(n_226), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_17), .A2(n_39), .B1(n_234), .B2(n_288), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_18), .A2(n_60), .B1(n_234), .B2(n_238), .Y(n_327) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_18), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_19), .B(n_234), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_20), .Y(n_141) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_21), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_22), .B(n_254), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_23), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_24), .B(n_254), .Y(n_302) );
INVx2_ASAP7_75t_L g236 ( .A(n_25), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_27), .B(n_234), .Y(n_233) );
OAI221xp5_ASAP7_75t_L g206 ( .A1(n_28), .A2(n_44), .B1(n_55), .B2(n_207), .C(n_208), .Y(n_206) );
INVxp67_ASAP7_75t_L g209 ( .A(n_28), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_29), .B(n_254), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_30), .A2(n_41), .B1(n_151), .B2(n_157), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_32), .A2(n_58), .B1(n_171), .B2(n_177), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_33), .Y(n_83) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_34), .B(n_234), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_35), .A2(n_68), .B1(n_288), .B2(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_36), .B(n_234), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_37), .B(n_234), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_38), .B(n_246), .Y(n_266) );
AOI22xp33_ASAP7_75t_SL g341 ( .A1(n_40), .A2(n_45), .B1(n_234), .B2(n_238), .Y(n_341) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_42), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_42), .B(n_234), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_43), .B(n_234), .Y(n_306) );
AO22x2_ASAP7_75t_L g106 ( .A1(n_44), .A2(n_64), .B1(n_97), .B2(n_101), .Y(n_106) );
INVxp67_ASAP7_75t_L g210 ( .A(n_44), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_46), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_47), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_48), .B(n_234), .Y(n_280) );
INVx1_ASAP7_75t_L g229 ( .A(n_49), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_50), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_51), .A2(n_192), .B1(n_193), .B2(n_200), .Y(n_191) );
INVx1_ASAP7_75t_L g200 ( .A(n_51), .Y(n_200) );
AO32x2_ASAP7_75t_L g323 ( .A1(n_52), .A2(n_251), .A3(n_259), .B1(n_324), .B2(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g244 ( .A(n_53), .Y(n_244) );
INVx1_ASAP7_75t_L g297 ( .A(n_54), .Y(n_297) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_55), .A2(n_71), .B1(n_97), .B2(n_98), .Y(n_104) );
INVx1_ASAP7_75t_L g189 ( .A(n_56), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_57), .B(n_238), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_59), .Y(n_130) );
INVx1_ASAP7_75t_L g543 ( .A(n_60), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_61), .B(n_288), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_62), .B(n_238), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_63), .Y(n_137) );
INVx2_ASAP7_75t_L g227 ( .A(n_65), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_66), .A2(n_75), .B1(n_162), .B2(n_165), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_67), .B(n_238), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_69), .A2(n_77), .B1(n_238), .B2(n_239), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_70), .A2(n_72), .B1(n_180), .B2(n_184), .Y(n_179) );
INVx1_ASAP7_75t_L g97 ( .A(n_73), .Y(n_97) );
INVx1_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_74), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_76), .Y(n_107) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_203), .B1(n_216), .B2(n_521), .C(n_529), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_187), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_84), .B2(n_85), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AOI22xp5_ASAP7_75t_SL g530 ( .A1(n_84), .A2(n_85), .B1(n_531), .B2(n_532), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_148), .Y(n_87) );
NOR3xp33_ASAP7_75t_L g88 ( .A(n_89), .B(n_113), .C(n_136), .Y(n_88) );
OAI22xp5_ASAP7_75t_L g89 ( .A1(n_90), .A2(n_91), .B1(n_107), .B2(n_108), .Y(n_89) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_94), .B(n_102), .Y(n_93) );
INVx2_ASAP7_75t_L g176 ( .A(n_94), .Y(n_176) );
OR2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_100), .Y(n_94) );
AND2x2_ASAP7_75t_L g112 ( .A(n_95), .B(n_100), .Y(n_112) );
AND2x2_ASAP7_75t_L g156 ( .A(n_95), .B(n_128), .Y(n_156) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g117 ( .A(n_96), .B(n_100), .Y(n_117) );
AND2x2_ASAP7_75t_L g129 ( .A(n_96), .B(n_106), .Y(n_129) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_99), .Y(n_101) );
INVx2_ASAP7_75t_L g128 ( .A(n_100), .Y(n_128) );
INVx1_ASAP7_75t_L g186 ( .A(n_100), .Y(n_186) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2x1p5_ASAP7_75t_L g111 ( .A(n_103), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g178 ( .A(n_103), .B(n_156), .Y(n_178) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g119 ( .A(n_104), .Y(n_119) );
INVx1_ASAP7_75t_L g127 ( .A(n_104), .Y(n_127) );
INVx1_ASAP7_75t_L g147 ( .A(n_104), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_104), .B(n_106), .Y(n_160) );
AND2x2_ASAP7_75t_L g118 ( .A(n_105), .B(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g155 ( .A(n_106), .B(n_147), .Y(n_155) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g168 ( .A(n_112), .B(n_118), .Y(n_168) );
AND2x2_ASAP7_75t_L g183 ( .A(n_112), .B(n_155), .Y(n_183) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_120), .B1(n_121), .B2(n_130), .C(n_131), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx4_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g144 ( .A(n_117), .Y(n_144) );
AND2x2_ASAP7_75t_L g164 ( .A(n_118), .B(n_156), .Y(n_164) );
AND2x6_ASAP7_75t_L g175 ( .A(n_118), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
INVx1_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
AND2x4_ASAP7_75t_L g134 ( .A(n_129), .B(n_135), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g139 ( .A(n_129), .B(n_140), .Y(n_139) );
BUFx4f_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
BUFx12f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_141), .B2(n_142), .Y(n_136) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp67_ASAP7_75t_L g148 ( .A(n_149), .B(n_169), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_161), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x4_ASAP7_75t_L g158 ( .A(n_156), .B(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x6_ASAP7_75t_L g185 ( .A(n_160), .B(n_186), .Y(n_185) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_179), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
INVx11_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx8_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B1(n_201), .B2(n_202), .Y(n_187) );
INVx1_ASAP7_75t_L g201 ( .A(n_188), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_191), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_204), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
AND3x1_ASAP7_75t_SL g205 ( .A(n_206), .B(n_211), .C(n_214), .Y(n_205) );
INVxp67_ASAP7_75t_L g536 ( .A(n_206), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_211), .A2(n_540), .B(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g548 ( .A(n_211), .Y(n_548) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_212), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_212), .B(n_215), .Y(n_542) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OR2x2_ASAP7_75t_SL g547 ( .A(n_214), .B(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR3x1_ASAP7_75t_L g218 ( .A(n_219), .B(n_449), .C(n_498), .Y(n_218) );
NAND5xp2_ASAP7_75t_L g219 ( .A(n_220), .B(n_364), .C(n_392), .D(n_422), .E(n_436), .Y(n_219) );
AOI221xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_282), .B1(n_314), .B2(n_319), .C(n_330), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_255), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_222), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g344 ( .A(n_223), .Y(n_344) );
AND2x2_ASAP7_75t_L g352 ( .A(n_223), .B(n_258), .Y(n_352) );
AND2x2_ASAP7_75t_L g375 ( .A(n_223), .B(n_257), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_223), .B(n_269), .Y(n_390) );
OR2x2_ASAP7_75t_L g399 ( .A(n_223), .B(n_337), .Y(n_399) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_223), .Y(n_402) );
AND2x2_ASAP7_75t_L g510 ( .A(n_223), .B(n_337), .Y(n_510) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_231), .B(n_253), .Y(n_223) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_224), .A2(n_270), .B(n_281), .Y(n_269) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_226), .Y(n_259) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_227), .B(n_228), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_243), .B(n_251), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_237), .B(n_240), .Y(n_232) );
INVx3_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
BUFx3_ASAP7_75t_L g326 ( .A(n_235), .Y(n_326) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g239 ( .A(n_236), .Y(n_239) );
INVx1_ASAP7_75t_L g247 ( .A(n_236), .Y(n_247) );
INVx2_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_240), .A2(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
O2A1O1Ixp5_ASAP7_75t_SL g295 ( .A1(n_240), .A2(n_296), .B(n_297), .C(n_298), .Y(n_295) );
INVx5_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g324 ( .A1(n_241), .A2(n_250), .B1(n_325), .B2(n_327), .Y(n_324) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_242), .Y(n_250) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_242), .Y(n_277) );
INVx1_ASAP7_75t_L g309 ( .A(n_242), .Y(n_309) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_248), .C(n_249), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_245), .A2(n_267), .B(n_279), .C(n_280), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_245), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_245), .B(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_249), .A2(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_250), .A2(n_267), .B1(n_287), .B2(n_289), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_250), .A2(n_267), .B1(n_340), .B2(n_341), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_251), .B(n_338), .C(n_339), .Y(n_363) );
BUFx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_252), .A2(n_261), .B(n_264), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_252), .A2(n_271), .B(n_278), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_252), .A2(n_295), .B(n_299), .Y(n_294) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_252), .A2(n_305), .B(n_310), .Y(n_304) );
INVx4_ASAP7_75t_SL g528 ( .A(n_252), .Y(n_528) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_254), .A2(n_294), .B(n_302), .Y(n_293) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_254), .A2(n_304), .B(n_313), .Y(n_303) );
INVx2_ASAP7_75t_L g328 ( .A(n_254), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_255), .B(n_402), .Y(n_458) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OAI311xp33_ASAP7_75t_L g400 ( .A1(n_256), .A2(n_401), .A3(n_402), .B1(n_403), .C1(n_418), .Y(n_400) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_269), .Y(n_256) );
AND2x2_ASAP7_75t_L g361 ( .A(n_257), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g368 ( .A(n_257), .Y(n_368) );
AND2x2_ASAP7_75t_L g489 ( .A(n_257), .B(n_318), .Y(n_489) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_258), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g345 ( .A(n_258), .B(n_269), .Y(n_345) );
AND2x2_ASAP7_75t_L g397 ( .A(n_258), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g411 ( .A(n_258), .B(n_344), .Y(n_411) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_268), .Y(n_258) );
INVx4_ASAP7_75t_L g338 ( .A(n_259), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_266), .B(n_267), .Y(n_264) );
INVx2_ASAP7_75t_L g318 ( .A(n_269), .Y(n_318) );
AND2x2_ASAP7_75t_L g360 ( .A(n_269), .B(n_344), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B(n_274), .C(n_275), .Y(n_271) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_276), .A2(n_300), .B(n_301), .Y(n_299) );
INVx4_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g526 ( .A(n_277), .Y(n_526) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_290), .Y(n_282) );
OR2x2_ASAP7_75t_L g455 ( .A(n_283), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_283), .B(n_461), .Y(n_472) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_284), .B(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
AND2x2_ASAP7_75t_L g396 ( .A(n_285), .B(n_323), .Y(n_396) );
AND2x2_ASAP7_75t_L g407 ( .A(n_285), .B(n_303), .Y(n_407) );
AND2x2_ASAP7_75t_L g416 ( .A(n_285), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_290), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_290), .B(n_357), .Y(n_401) );
INVx2_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g388 ( .A(n_291), .B(n_347), .Y(n_388) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_303), .Y(n_291) );
INVx2_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
AND2x2_ASAP7_75t_L g415 ( .A(n_292), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g333 ( .A(n_293), .Y(n_333) );
OR2x2_ASAP7_75t_L g432 ( .A(n_293), .B(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_293), .Y(n_495) );
AND2x2_ASAP7_75t_L g334 ( .A(n_303), .B(n_329), .Y(n_334) );
INVx1_ASAP7_75t_L g355 ( .A(n_303), .Y(n_355) );
AND2x2_ASAP7_75t_L g376 ( .A(n_303), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g417 ( .A(n_303), .Y(n_417) );
INVx1_ASAP7_75t_L g433 ( .A(n_303), .Y(n_433) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_303), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_316), .B(n_421), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_316), .A2(n_406), .B1(n_455), .B2(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g498 ( .A1(n_317), .A2(n_499), .B(n_501), .C(n_519), .Y(n_498) );
INVx2_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
AND2x2_ASAP7_75t_L g409 ( .A(n_318), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g420 ( .A(n_318), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_319), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g393 ( .A(n_320), .B(n_357), .Y(n_393) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g425 ( .A(n_321), .B(n_416), .Y(n_425) );
AND2x2_ASAP7_75t_L g444 ( .A(n_321), .B(n_358), .Y(n_444) );
AND2x4_ASAP7_75t_L g380 ( .A(n_322), .B(n_354), .Y(n_380) );
AND2x2_ASAP7_75t_L g518 ( .A(n_322), .B(n_494), .Y(n_518) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_329), .Y(n_322) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
INVx1_ASAP7_75t_L g457 ( .A(n_323), .Y(n_457) );
OR2x2_ASAP7_75t_L g348 ( .A(n_329), .B(n_333), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_358), .Y(n_357) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_329), .B(n_378), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_346), .B2(n_349), .C(n_353), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_332), .A2(n_354), .B(n_356), .C(n_359), .Y(n_353) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_333), .B(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_333), .B(n_355), .Y(n_461) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_333), .Y(n_468) );
AND2x2_ASAP7_75t_L g386 ( .A(n_334), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g423 ( .A(n_334), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_345), .Y(n_335) );
INVx2_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
AOI222xp33_ASAP7_75t_L g463 ( .A1(n_336), .A2(n_347), .B1(n_464), .B2(n_466), .C1(n_467), .C2(n_469), .Y(n_463) );
AND2x2_ASAP7_75t_L g520 ( .A(n_336), .B(n_489), .Y(n_520) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .Y(n_336) );
INVx1_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
AO21x1_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B(n_342), .Y(n_337) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g362 ( .A(n_343), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g448 ( .A(n_345), .B(n_382), .Y(n_448) );
AOI21xp33_ASAP7_75t_L g459 ( .A1(n_346), .A2(n_460), .B(n_462), .Y(n_459) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_347), .B(n_354), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_347), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx3_ASAP7_75t_L g413 ( .A(n_351), .Y(n_413) );
OR2x2_ASAP7_75t_L g465 ( .A(n_351), .B(n_387), .Y(n_465) );
AND2x2_ASAP7_75t_L g381 ( .A(n_352), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g419 ( .A(n_352), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_352), .B(n_413), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_352), .B(n_409), .Y(n_435) );
AND2x2_ASAP7_75t_L g439 ( .A(n_352), .B(n_421), .Y(n_439) );
INVxp67_ASAP7_75t_L g371 ( .A(n_354), .Y(n_371) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_356), .A2(n_429), .B1(n_434), .B2(n_435), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_356), .B(n_461), .Y(n_491) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g477 ( .A(n_357), .B(n_468), .Y(n_477) );
AND2x2_ASAP7_75t_L g506 ( .A(n_357), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g511 ( .A(n_357), .B(n_461), .Y(n_511) );
INVx1_ASAP7_75t_L g424 ( .A(n_358), .Y(n_424) );
BUFx2_ASAP7_75t_L g430 ( .A(n_358), .Y(n_430) );
INVx1_ASAP7_75t_L g515 ( .A(n_359), .Y(n_515) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_360), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
NOR2x1_ASAP7_75t_L g367 ( .A(n_362), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g374 ( .A(n_362), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g383 ( .A(n_362), .Y(n_383) );
INVx3_ASAP7_75t_L g421 ( .A(n_362), .Y(n_421) );
OR2x2_ASAP7_75t_L g487 ( .A(n_362), .B(n_488), .Y(n_487) );
AOI211xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B(n_372), .C(n_384), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_365), .A2(n_502), .B1(n_509), .B2(n_511), .C(n_512), .Y(n_501) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_379), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_375), .B(n_413), .Y(n_427) );
AND2x2_ASAP7_75t_L g469 ( .A(n_375), .B(n_409), .Y(n_469) );
INVx1_ASAP7_75t_SL g482 ( .A(n_376), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_376), .B(n_430), .Y(n_485) );
INVx1_ASAP7_75t_L g503 ( .A(n_377), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_381), .A2(n_471), .B1(n_473), .B2(n_477), .C(n_478), .Y(n_470) );
AND2x2_ASAP7_75t_L g497 ( .A(n_382), .B(n_489), .Y(n_497) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g481 ( .A(n_383), .Y(n_481) );
AOI21xp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_388), .B(n_389), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g452 ( .A(n_387), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
INVx1_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B(n_397), .C(n_400), .Y(n_392) );
OAI31xp33_ASAP7_75t_L g519 ( .A1(n_393), .A2(n_431), .A3(n_518), .B(n_520), .Y(n_519) );
INVxp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g493 ( .A(n_396), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_SL g514 ( .A(n_396), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_398), .B(n_413), .Y(n_441) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g516 ( .A(n_399), .B(n_413), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_408), .B1(n_412), .B2(n_415), .Y(n_403) );
NAND2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_407), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_407), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g446 ( .A(n_407), .B(n_430), .Y(n_446) );
AND2x2_ASAP7_75t_L g500 ( .A(n_407), .B(n_495), .Y(n_500) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g475 ( .A(n_411), .Y(n_475) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g478 ( .A1(n_413), .A2(n_447), .A3(n_479), .B1(n_481), .B2(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_416), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g476 ( .A(n_420), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B(n_426), .C(n_428), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_424), .B(n_461), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_425), .A2(n_437), .B1(n_438), .B2(n_439), .C(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g437 ( .A(n_435), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_445), .B2(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_445), .B(n_503), .C(n_504), .D(n_505), .Y(n_502) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_450), .B(n_463), .C(n_470), .D(n_483), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B(n_458), .C(n_459), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g480 ( .A(n_456), .Y(n_480) );
INVx2_ASAP7_75t_L g504 ( .A(n_461), .Y(n_504) );
OR2x2_ASAP7_75t_L g513 ( .A(n_468), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_486), .B(n_490), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g509 ( .A(n_489), .B(n_510), .Y(n_509) );
AOI21xp33_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_492), .B(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_512) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx1_ASAP7_75t_L g541 ( .A(n_524), .Y(n_541) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI322xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_533), .A3(n_537), .B1(n_538), .B2(n_543), .C1(n_544), .C2(n_545), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_531), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
endmodule