module fake_jpeg_14934_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

AO21x1_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_11),
.B(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_20),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_3),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_12),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_18),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_5),
.B(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_16),
.B1(n_13),
.B2(n_9),
.Y(n_31)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

AO221x1_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.C(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_17),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.C(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_35),
.C(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_43)
);


endmodule