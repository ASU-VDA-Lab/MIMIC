module fake_jpeg_15078_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_49),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_47),
.Y(n_70)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_22),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx11_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_27),
.C(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_27),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_34),
.B1(n_23),
.B2(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_74),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_83),
.Y(n_88)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_77),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_74)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_53),
.B1(n_41),
.B2(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_58),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_38),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_38),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_38),
.C(n_40),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_78),
.B1(n_76),
.B2(n_67),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_113),
.B1(n_118),
.B2(n_124),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_78),
.B1(n_83),
.B2(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_65),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_102),
.B1(n_94),
.B2(n_100),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_106),
.B(n_86),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_22),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_130),
.Y(n_151)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_69),
.B1(n_59),
.B2(n_62),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_133),
.Y(n_139)
);

INVx2_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_103),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_78),
.B1(n_19),
.B2(n_25),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_89),
.B(n_99),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_34),
.B1(n_108),
.B2(n_30),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_132),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_125),
.B(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_85),
.C(n_92),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_150),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_107),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_100),
.Y(n_147)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_84),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_159),
.B1(n_124),
.B2(n_131),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_1),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_162),
.C(n_17),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_160),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_115),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_168),
.B1(n_175),
.B2(n_178),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_129),
.B1(n_112),
.B2(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_172),
.A2(n_177),
.B(n_187),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_174),
.B(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_113),
.B1(n_123),
.B2(n_75),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_141),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_111),
.B(n_3),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_19),
.B1(n_32),
.B2(n_29),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_143),
.C(n_145),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_185),
.C(n_30),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_141),
.C(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_144),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_37),
.B1(n_36),
.B2(n_29),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_189),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_202),
.C(n_184),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_183),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_196),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_151),
.Y(n_198)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_140),
.B1(n_158),
.B2(n_144),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_185),
.B1(n_165),
.B2(n_169),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_203),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_206),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_177),
.B1(n_179),
.B2(n_187),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_199),
.B(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_169),
.B1(n_164),
.B2(n_165),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_221),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_176),
.B1(n_164),
.B2(n_171),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_201),
.B1(n_204),
.B2(n_202),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_170),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_170),
.C(n_37),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_204),
.A2(n_146),
.B1(n_14),
.B2(n_13),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_205),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_235),
.B(n_230),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_218),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_233),
.B(n_234),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_199),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_199),
.B1(n_146),
.B2(n_28),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_208),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_227),
.B(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_217),
.C(n_211),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_214),
.B1(n_209),
.B2(n_222),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_241),
.Y(n_248)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_229),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_28),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_14),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_253),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_244),
.A2(n_13),
.B(n_12),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_10),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_237),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_2),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.C(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_2),
.Y(n_261)
);

AOI31xp33_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_256),
.C(n_255),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_265),
.A2(n_266),
.B(n_7),
.Y(n_267)
);

OAI311xp33_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.C1(n_8),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_264),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_8),
.B(n_9),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_8),
.Y(n_270)
);


endmodule