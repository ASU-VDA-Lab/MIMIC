module fake_jpeg_1007_n_127 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_50),
.Y(n_51)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_39),
.B1(n_40),
.B2(n_50),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_37),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_69),
.B1(n_58),
.B2(n_56),
.Y(n_73)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_43),
.C(n_42),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_60),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_66),
.Y(n_81)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_78),
.B1(n_62),
.B2(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_80),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_58),
.B1(n_55),
.B2(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_0),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_2),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_71),
.B1(n_65),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_95),
.B1(n_32),
.B2(n_27),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_15),
.B1(n_30),
.B2(n_28),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_72),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_2),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_105),
.B(n_18),
.C(n_16),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_26),
.B(n_21),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_20),
.C(n_19),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_109),
.C(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.C(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_14),
.C(n_5),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_107),
.B(n_106),
.C(n_6),
.D(n_7),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_4),
.B(n_5),
.Y(n_116)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_114),
.C(n_111),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_8),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_6),
.B(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_9),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_122),
.B(n_123),
.C(n_12),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_12),
.C(n_10),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_11),
.Y(n_127)
);


endmodule