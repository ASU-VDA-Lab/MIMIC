module fake_jpeg_13832_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_49),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_39),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_38),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_42),
.B1(n_37),
.B2(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_38),
.B1(n_31),
.B2(n_17),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_69),
.B1(n_8),
.B2(n_20),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_60),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

AO21x2_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_13),
.B(n_26),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_52),
.A2(n_12),
.B1(n_25),
.B2(n_21),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_27),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_74),
.B1(n_69),
.B2(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_3),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_86),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_4),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_7),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_87),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_77),
.B(n_81),
.C(n_80),
.D(n_85),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_99),
.B(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_82),
.C(n_96),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_93),
.Y(n_106)
);


endmodule