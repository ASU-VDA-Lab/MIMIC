module fake_netlist_5_186_n_1626 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1626);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1626;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_370;
wire n_976;
wire n_1449;
wire n_1566;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1598;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1617;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1591;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_1351;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_114),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_32),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_176),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_224),
.Y(n_348)
);

BUFx8_ASAP7_75t_SL g349 ( 
.A(n_251),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_174),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_178),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_21),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_197),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_15),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_171),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_222),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_309),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_94),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_140),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_235),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_228),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_218),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_125),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_15),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_18),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_34),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_268),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_260),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_191),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_3),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_138),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_261),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_180),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_188),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_170),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_335),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_271),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_200),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_199),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_85),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_280),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_93),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_86),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_186),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_291),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_301),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_319),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_341),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_90),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_50),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_71),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_213),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_10),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_80),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_290),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_75),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_211),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_79),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_243),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_130),
.Y(n_408)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_294),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_42),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_151),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_25),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_244),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_274),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_190),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_30),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_304),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_279),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_26),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_266),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_177),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_103),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_6),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_326),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_343),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_5),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_265),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_72),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_72),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_132),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_127),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_311),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_10),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_183),
.Y(n_435)
);

BUFx2_ASAP7_75t_R g436 ( 
.A(n_102),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_204),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_209),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_322),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_17),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_14),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_315),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_86),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_139),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_29),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_56),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_142),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_262),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_93),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_94),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_207),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_201),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_137),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_168),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_342),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_328),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_234),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_246),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_45),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_148),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_219),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_111),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_5),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_87),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_42),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_263),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_117),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_340),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_334),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_157),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_344),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_65),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_339),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_250),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_119),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_299),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_329),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_272),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_314),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_162),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_49),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_220),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_89),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_298),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_227),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_308),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_293),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_50),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_254),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_27),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_70),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_109),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_17),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_337),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_338),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_71),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_233),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_179),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_20),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_276),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_238),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_96),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_256),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_156),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_126),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_324),
.Y(n_506)
);

BUFx10_ASAP7_75t_L g507 ( 
.A(n_196),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_288),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_214),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_295),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_77),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_312),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_33),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_193),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_64),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_136),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_189),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_8),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_259),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_110),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_62),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_273),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_336),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_52),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_321),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_253),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_208),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_83),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_88),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_277),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_48),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_323),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_198),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_0),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_39),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_327),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_43),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_49),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g539 ( 
.A(n_317),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_13),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_154),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_185),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_303),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_24),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_47),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_249),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_166),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_57),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_247),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_28),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_63),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_248),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_267),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_141),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_16),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_48),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_67),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_163),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_242),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_13),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_223),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_210),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_2),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_101),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_221),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_215),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_24),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_63),
.Y(n_568)
);

HB1xp67_ASAP7_75t_SL g569 ( 
.A(n_226),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_4),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_97),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_167),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_87),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_332),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_164),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_67),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_100),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_134),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_287),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_85),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_255),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_283),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_479),
.B(n_0),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_360),
.B(n_1),
.Y(n_584)
);

BUFx8_ASAP7_75t_SL g585 ( 
.A(n_349),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_497),
.B(n_1),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_367),
.B(n_104),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_367),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_471),
.B(n_2),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_471),
.B(n_3),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_424),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_4),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_424),
.B(n_6),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_367),
.B(n_460),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_367),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_460),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_424),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_417),
.B(n_7),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_370),
.B(n_571),
.Y(n_599)
);

BUFx8_ASAP7_75t_SL g600 ( 
.A(n_349),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_7),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_460),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_424),
.B(n_8),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_547),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_424),
.B(n_9),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_389),
.B(n_9),
.Y(n_608)
);

BUFx8_ASAP7_75t_L g609 ( 
.A(n_424),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_547),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_11),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_424),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_487),
.B(n_11),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

BUFx8_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_395),
.B(n_12),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_573),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_407),
.B(n_12),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_426),
.B(n_14),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_573),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_576),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_576),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_547),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_512),
.B(n_16),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_550),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_576),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_549),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_550),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_435),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_502),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_18),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_426),
.B(n_19),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_409),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_454),
.B(n_492),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g640 ( 
.A(n_387),
.B(n_19),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_454),
.B(n_20),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_549),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

BUFx8_ASAP7_75t_SL g644 ( 
.A(n_387),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_500),
.B(n_21),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_500),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_353),
.B(n_22),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_370),
.B(n_22),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_429),
.B(n_23),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_350),
.Y(n_650)
);

CKINVDCx11_ASAP7_75t_R g651 ( 
.A(n_429),
.Y(n_651)
);

BUFx8_ASAP7_75t_SL g652 ( 
.A(n_430),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_571),
.B(n_23),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_351),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_435),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_352),
.B(n_105),
.Y(n_656)
);

BUFx8_ASAP7_75t_SL g657 ( 
.A(n_430),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_435),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_356),
.B(n_25),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_409),
.B(n_26),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_362),
.B(n_27),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_540),
.B(n_28),
.Y(n_662)
);

XNOR2x2_ASAP7_75t_L g663 ( 
.A(n_440),
.B(n_29),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_364),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_365),
.B(n_30),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_368),
.B(n_31),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_409),
.B(n_31),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_507),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_373),
.B(n_32),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_369),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_418),
.B(n_33),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_345),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_507),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_448),
.B(n_34),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_353),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_507),
.B(n_391),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_409),
.B(n_35),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_466),
.B(n_35),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_377),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_346),
.Y(n_680)
);

BUFx8_ASAP7_75t_L g681 ( 
.A(n_391),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_409),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_374),
.B(n_36),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_347),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_409),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_489),
.B(n_36),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_376),
.B(n_37),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_493),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_378),
.B(n_37),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_427),
.B(n_38),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_409),
.Y(n_691)
);

BUFx12f_ASAP7_75t_L g692 ( 
.A(n_390),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_493),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_384),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_385),
.B(n_106),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_397),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_392),
.Y(n_697)
);

BUFx12f_ASAP7_75t_L g698 ( 
.A(n_398),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_530),
.B(n_38),
.Y(n_699)
);

BUFx8_ASAP7_75t_SL g700 ( 
.A(n_464),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_443),
.B(n_39),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_393),
.B(n_40),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_399),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_423),
.B(n_40),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_401),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_563),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_554),
.B(n_41),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_403),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_436),
.B(n_41),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_405),
.B(n_412),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_402),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_414),
.B(n_43),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_419),
.B(n_44),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_432),
.B(n_44),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_423),
.B(n_45),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_423),
.Y(n_717)
);

INVx5_ASAP7_75t_L g718 ( 
.A(n_567),
.Y(n_718)
);

INVx5_ASAP7_75t_L g719 ( 
.A(n_567),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_423),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_423),
.B(n_46),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_371),
.B(n_46),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_437),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_406),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_404),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_447),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_451),
.B(n_47),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_410),
.B(n_51),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_423),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_363),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_455),
.B(n_51),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_456),
.B(n_52),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_413),
.B(n_53),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_420),
.B(n_53),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_450),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_458),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_459),
.B(n_54),
.Y(n_737)
);

BUFx8_ASAP7_75t_L g738 ( 
.A(n_472),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_423),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_434),
.B(n_54),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_462),
.B(n_55),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_585),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_679),
.B(n_348),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_615),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_583),
.A2(n_411),
.B1(n_562),
.B2(n_363),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_588),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_SL g747 ( 
.A1(n_640),
.A2(n_464),
.B1(n_521),
.B2(n_411),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_589),
.A2(n_490),
.B1(n_491),
.B2(n_481),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_586),
.A2(n_579),
.B1(n_582),
.B2(n_562),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_589),
.A2(n_518),
.B1(n_524),
.B2(n_515),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_623),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_598),
.A2(n_445),
.B1(n_446),
.B2(n_441),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_618),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_R g754 ( 
.A1(n_584),
.A2(n_531),
.B1(n_568),
.B2(n_538),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_629),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_618),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_598),
.A2(n_463),
.B1(n_465),
.B2(n_449),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_703),
.B(n_354),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_592),
.A2(n_582),
.B1(n_579),
.B2(n_488),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_606),
.A2(n_496),
.B1(n_499),
.B2(n_483),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_599),
.B(n_355),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_621),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_630),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_606),
.A2(n_513),
.B1(n_528),
.B2(n_511),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_672),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_633),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_634),
.A2(n_529),
.B1(n_535),
.B2(n_534),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_730),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_676),
.A2(n_544),
.B1(n_545),
.B2(n_537),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_630),
.Y(n_770)
);

XOR2xp5_ASAP7_75t_L g771 ( 
.A(n_649),
.B(n_521),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_666),
.A2(n_551),
.B1(n_555),
.B2(n_548),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_658),
.A2(n_557),
.B1(n_560),
.B2(n_556),
.Y(n_773)
);

AO22x2_ASAP7_75t_L g774 ( 
.A1(n_590),
.A2(n_580),
.B1(n_570),
.B2(n_476),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_588),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_655),
.B(n_673),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_670),
.B(n_357),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_658),
.A2(n_477),
.B1(n_486),
.B2(n_469),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_588),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_671),
.A2(n_674),
.B1(n_686),
.B2(n_678),
.Y(n_780)
);

AO22x2_ASAP7_75t_L g781 ( 
.A1(n_590),
.A2(n_498),
.B1(n_501),
.B2(n_494),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_709),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_L g783 ( 
.A1(n_709),
.A2(n_509),
.B1(n_514),
.B2(n_508),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_596),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_696),
.B(n_358),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_621),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_596),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_699),
.A2(n_361),
.B1(n_366),
.B2(n_359),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_705),
.B(n_372),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_624),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_600),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_711),
.B(n_375),
.Y(n_792)
);

INVx8_ASAP7_75t_L g793 ( 
.A(n_692),
.Y(n_793)
);

AO22x2_ASAP7_75t_L g794 ( 
.A1(n_601),
.A2(n_519),
.B1(n_520),
.B2(n_516),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_655),
.A2(n_533),
.B1(n_542),
.B2(n_523),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_725),
.B(n_655),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_684),
.B(n_553),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_707),
.A2(n_380),
.B1(n_381),
.B2(n_379),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_617),
.A2(n_575),
.B1(n_577),
.B2(n_559),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_626),
.A2(n_667),
.B1(n_677),
.B2(n_660),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_673),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_644),
.Y(n_802)
);

AO22x2_ASAP7_75t_L g803 ( 
.A1(n_601),
.A2(n_578),
.B1(n_57),
.B2(n_55),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_383),
.B1(n_386),
.B2(n_382),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_698),
.B(n_56),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_619),
.B(n_388),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_704),
.A2(n_396),
.B1(n_400),
.B2(n_394),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_596),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_668),
.B(n_408),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_624),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_722),
.A2(n_581),
.B1(n_574),
.B2(n_565),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_722),
.B(n_58),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_602),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_710),
.B(n_415),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_SL g815 ( 
.A1(n_715),
.A2(n_564),
.B1(n_561),
.B2(n_558),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_712),
.A2(n_474),
.B1(n_546),
.B2(n_543),
.Y(n_816)
);

AO22x2_ASAP7_75t_L g817 ( 
.A1(n_613),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_602),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_710),
.B(n_416),
.Y(n_819)
);

BUFx10_ASAP7_75t_L g820 ( 
.A(n_713),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_602),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_681),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_605),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_648),
.B(n_421),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_737),
.A2(n_552),
.B1(n_541),
.B2(n_536),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_721),
.A2(n_532),
.B1(n_527),
.B2(n_526),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_737),
.A2(n_525),
.B1(n_522),
.B2(n_517),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_714),
.A2(n_510),
.B1(n_506),
.B2(n_495),
.Y(n_828)
);

OAI22xp33_ASAP7_75t_L g829 ( 
.A1(n_647),
.A2(n_485),
.B1(n_484),
.B2(n_482),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_653),
.B(n_422),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_613),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_831)
);

XOR2xp5_ASAP7_75t_L g832 ( 
.A(n_663),
.B(n_425),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_659),
.A2(n_480),
.B1(n_478),
.B2(n_475),
.Y(n_833)
);

AO22x2_ASAP7_75t_L g834 ( 
.A1(n_620),
.A2(n_645),
.B1(n_641),
.B2(n_661),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_605),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_605),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_610),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_428),
.Y(n_838)
);

OAI22xp33_ASAP7_75t_R g839 ( 
.A1(n_727),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_839)
);

AO22x2_ASAP7_75t_L g840 ( 
.A1(n_620),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_840)
);

AO22x2_ASAP7_75t_L g841 ( 
.A1(n_641),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_610),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_733),
.B(n_431),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_610),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_647),
.A2(n_636),
.B1(n_593),
.B2(n_741),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_701),
.A2(n_453),
.B1(n_470),
.B2(n_468),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_813),
.A2(n_639),
.B(n_597),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_761),
.B(n_734),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_814),
.B(n_661),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_813),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_845),
.B(n_591),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_796),
.B(n_824),
.Y(n_852)
);

INVx4_ASAP7_75t_SL g853 ( 
.A(n_746),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_775),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_818),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_836),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_746),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_836),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_800),
.A2(n_593),
.B(n_603),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_779),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_784),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_787),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_808),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_780),
.B(n_806),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_821),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_823),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_830),
.B(n_740),
.Y(n_868)
);

INVxp33_ASAP7_75t_L g869 ( 
.A(n_771),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_819),
.B(n_665),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_835),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_837),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_842),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_767),
.B(n_662),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_746),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_844),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_816),
.B(n_635),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_816),
.B(n_608),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_753),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_744),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_828),
.B(n_611),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_768),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_753),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_751),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_802),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_770),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_770),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_756),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_755),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_763),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_777),
.B(n_690),
.Y(n_891)
);

XNOR2xp5_ASAP7_75t_L g892 ( 
.A(n_749),
.B(n_652),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_762),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_762),
.A2(n_597),
.B(n_607),
.Y(n_894)
);

XNOR2xp5_ASAP7_75t_L g895 ( 
.A(n_745),
.B(n_657),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_786),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_828),
.A2(n_812),
.B(n_846),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_838),
.B(n_680),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_786),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_645),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_790),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_811),
.B(n_650),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_825),
.B(n_650),
.Y(n_903)
);

XOR2xp5_ASAP7_75t_L g904 ( 
.A(n_742),
.B(n_433),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_790),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_810),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_834),
.B(n_612),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_810),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_843),
.B(n_743),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_766),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_827),
.B(n_650),
.Y(n_911)
);

AND2x2_ASAP7_75t_SL g912 ( 
.A(n_759),
.B(n_665),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_765),
.B(n_654),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_834),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_758),
.B(n_688),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_772),
.B(n_669),
.Y(n_916)
);

XOR2xp5_ASAP7_75t_L g917 ( 
.A(n_791),
.B(n_438),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_748),
.Y(n_918)
);

INVxp33_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_748),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_750),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_750),
.Y(n_922)
);

XNOR2xp5_ASAP7_75t_L g923 ( 
.A(n_832),
.B(n_700),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_809),
.B(n_669),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_797),
.B(n_637),
.Y(n_925)
);

XOR2xp5_ASAP7_75t_L g926 ( 
.A(n_760),
.B(n_439),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_774),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_789),
.B(n_792),
.Y(n_928)
);

BUFx5_ASAP7_75t_L g929 ( 
.A(n_820),
.Y(n_929)
);

XOR2xp5_ASAP7_75t_L g930 ( 
.A(n_764),
.B(n_442),
.Y(n_930)
);

AOI21x1_ASAP7_75t_L g931 ( 
.A1(n_776),
.A2(n_685),
.B(n_682),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_774),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_781),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_820),
.B(n_688),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_781),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_794),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_803),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_794),
.Y(n_938)
);

XNOR2x2_ASAP7_75t_L g939 ( 
.A(n_841),
.B(n_651),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_914),
.B(n_765),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_905),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_893),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_891),
.B(n_928),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_896),
.Y(n_944)
);

OR2x6_ASAP7_75t_L g945 ( 
.A(n_918),
.B(n_840),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_899),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_909),
.B(n_803),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_865),
.B(n_788),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_898),
.B(n_840),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_865),
.B(n_841),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_905),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_849),
.B(n_683),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_901),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_912),
.B(n_683),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_905),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_852),
.B(n_817),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_925),
.B(n_798),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_925),
.B(n_829),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_905),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_879),
.B(n_801),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_924),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_929),
.B(n_877),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_894),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_906),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_908),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_849),
.B(n_687),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_883),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_910),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_882),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_860),
.A2(n_695),
.B(n_656),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_868),
.B(n_817),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_933),
.B(n_687),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_895),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_858),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_886),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_878),
.A2(n_815),
.B1(n_826),
.B2(n_807),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_848),
.B(n_656),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_931),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_924),
.B(n_831),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_907),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_934),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_847),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_860),
.A2(n_695),
.B(n_656),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_900),
.B(n_656),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_854),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_880),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_870),
.B(n_831),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_920),
.B(n_793),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_870),
.B(n_689),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_907),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_884),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_900),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_851),
.B(n_689),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_921),
.B(n_833),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_889),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_851),
.B(n_702),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_900),
.B(n_695),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_915),
.B(n_897),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_897),
.B(n_702),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_887),
.Y(n_1000)
);

NOR2xp67_ASAP7_75t_L g1001 ( 
.A(n_885),
.B(n_822),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_850),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_877),
.B(n_731),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_855),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_900),
.B(n_695),
.Y(n_1005)
);

NAND2x1p5_ASAP7_75t_L g1006 ( 
.A(n_927),
.B(n_731),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_878),
.A2(n_799),
.B(n_732),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_912),
.B(n_732),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_900),
.B(n_643),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_902),
.B(n_643),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_881),
.B(n_724),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_881),
.B(n_752),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_902),
.A2(n_757),
.B(n_804),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_856),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_903),
.A2(n_769),
.B(n_587),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_903),
.B(n_724),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_911),
.B(n_643),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_911),
.B(n_735),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_916),
.A2(n_587),
.B(n_778),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_913),
.B(n_646),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_935),
.B(n_735),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_936),
.A2(n_754),
.B1(n_782),
.B2(n_783),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_675),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_861),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_929),
.B(n_874),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_862),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_938),
.A2(n_587),
.B(n_691),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_913),
.B(n_646),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_857),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_863),
.B(n_805),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_859),
.Y(n_1031)
);

AND2x2_ASAP7_75t_SL g1032 ( 
.A(n_937),
.B(n_839),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_888),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_890),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_864),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_929),
.B(n_675),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_929),
.B(n_646),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_964),
.Y(n_1038)
);

NOR2x1_ASAP7_75t_L g1039 ( 
.A(n_962),
.B(n_805),
.Y(n_1039)
);

AO21x2_ASAP7_75t_L g1040 ( 
.A1(n_970),
.A2(n_867),
.B(n_866),
.Y(n_1040)
);

BUFx2_ASAP7_75t_SL g1041 ( 
.A(n_969),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_993),
.B(n_929),
.Y(n_1042)
);

OR2x6_ASAP7_75t_L g1043 ( 
.A(n_969),
.B(n_793),
.Y(n_1043)
);

AND2x6_ASAP7_75t_L g1044 ( 
.A(n_992),
.B(n_871),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_961),
.B(n_937),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_961),
.B(n_872),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_993),
.B(n_929),
.Y(n_1047)
);

CKINVDCx6p67_ASAP7_75t_R g1048 ( 
.A(n_988),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_968),
.Y(n_1049)
);

OR2x2_ASAP7_75t_L g1050 ( 
.A(n_948),
.B(n_910),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_964),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_951),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1011),
.B(n_932),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1011),
.B(n_932),
.Y(n_1055)
);

CKINVDCx6p67_ASAP7_75t_R g1056 ( 
.A(n_988),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_965),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_996),
.B(n_873),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_944),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_946),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_L g1061 ( 
.A(n_980),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_943),
.B(n_919),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_957),
.B(n_919),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_946),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_1021),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_1021),
.B(n_876),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_953),
.Y(n_1067)
);

AND2x2_ASAP7_75t_SL g1068 ( 
.A(n_954),
.B(n_939),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1021),
.B(n_853),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_952),
.B(n_853),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_987),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_998),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_953),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_951),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_988),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_992),
.B(n_717),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_980),
.B(n_926),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_952),
.B(n_853),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_952),
.B(n_858),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_1016),
.Y(n_1080)
);

NAND2x1p5_ASAP7_75t_L g1081 ( 
.A(n_980),
.B(n_858),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_966),
.B(n_858),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_943),
.B(n_930),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1003),
.B(n_869),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_965),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_977),
.B(n_107),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1023),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_996),
.B(n_875),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_999),
.B(n_875),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1003),
.B(n_892),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_951),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_980),
.B(n_875),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_987),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_998),
.Y(n_1094)
);

AO21x2_ASAP7_75t_L g1095 ( 
.A1(n_983),
.A2(n_729),
.B(n_720),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1014),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1016),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1012),
.B(n_904),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1018),
.B(n_981),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_966),
.B(n_875),
.Y(n_1100)
);

BUFx4f_ASAP7_75t_L g1101 ( 
.A(n_980),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_988),
.B(n_614),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_990),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1018),
.B(n_917),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_990),
.B(n_773),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_979),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_990),
.B(n_625),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_994),
.B(n_923),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_973),
.Y(n_1109)
);

BUFx2_ASAP7_75t_SL g1110 ( 
.A(n_1001),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_951),
.Y(n_1111)
);

BUFx8_ASAP7_75t_SL g1112 ( 
.A(n_973),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_979),
.B(n_628),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_986),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_1030),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_951),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_966),
.B(n_716),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_999),
.Y(n_1118)
);

AND2x6_ASAP7_75t_L g1119 ( 
.A(n_1008),
.B(n_739),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_958),
.B(n_654),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1063),
.A2(n_954),
.B1(n_1013),
.B2(n_990),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1091),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1063),
.A2(n_954),
.B1(n_990),
.B2(n_1007),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1054),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_1091),
.Y(n_1125)
);

BUFx4_ASAP7_75t_SL g1126 ( 
.A(n_1043),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1059),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1091),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1060),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1097),
.B(n_1072),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1064),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1049),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1116),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1067),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1118),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1115),
.Y(n_1136)
);

BUFx8_ASAP7_75t_L g1137 ( 
.A(n_1071),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1077),
.A2(n_1008),
.B1(n_1025),
.B2(n_950),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1114),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1061),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1093),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1118),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1061),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1073),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_1101),
.B(n_959),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1106),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1050),
.B(n_1025),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1075),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_1116),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1101),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1116),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1096),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1072),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1097),
.B(n_950),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1094),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1045),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1038),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_1041),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1051),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1103),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1057),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1103),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1094),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_1074),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1074),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1085),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1087),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1081),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1117),
.Y(n_1169)
);

BUFx2_ASAP7_75t_SL g1170 ( 
.A(n_1070),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1053),
.B(n_949),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1070),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_1078),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1078),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1117),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1077),
.A2(n_976),
.B1(n_947),
.B2(n_971),
.Y(n_1176)
);

CKINVDCx14_ASAP7_75t_R g1177 ( 
.A(n_1109),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1043),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1081),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1092),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1084),
.Y(n_1181)
);

INVx6_ASAP7_75t_SL g1182 ( 
.A(n_1043),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1092),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1052),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1045),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1058),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1065),
.B(n_967),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1089),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1052),
.B(n_959),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1127),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1138),
.A2(n_1098),
.B1(n_1080),
.B2(n_1108),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_SL g1192 ( 
.A1(n_1147),
.A2(n_1080),
.B1(n_1042),
.B2(n_1047),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1158),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1157),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1181),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1178),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1157),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1176),
.A2(n_1062),
.B1(n_1104),
.B2(n_1099),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1121),
.A2(n_1022),
.B(n_1090),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1127),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1132),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1186),
.B(n_1055),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1177),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1165),
.Y(n_1204)
);

INVx6_ASAP7_75t_L g1205 ( 
.A(n_1137),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1132),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1178),
.Y(n_1207)
);

BUFx10_ASAP7_75t_L g1208 ( 
.A(n_1167),
.Y(n_1208)
);

INVx8_ASAP7_75t_L g1209 ( 
.A(n_1160),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1131),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1131),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1171),
.B(n_1083),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1123),
.A2(n_1068),
.B1(n_1105),
.B2(n_1015),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1130),
.A2(n_1105),
.B1(n_1089),
.B2(n_1042),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1171),
.A2(n_947),
.B1(n_971),
.B2(n_956),
.Y(n_1215)
);

BUFx8_ASAP7_75t_L g1216 ( 
.A(n_1136),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1137),
.A2(n_1032),
.B1(n_1110),
.B2(n_632),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1137),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1153),
.A2(n_1032),
.B1(n_949),
.B2(n_956),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1154),
.A2(n_940),
.B1(n_1047),
.B2(n_1039),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1153),
.A2(n_839),
.B1(n_754),
.B2(n_1088),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1155),
.A2(n_1032),
.B1(n_1066),
.B2(n_994),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1141),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1134),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1136),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1148),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1134),
.A2(n_1088),
.B1(n_940),
.B2(n_1058),
.Y(n_1227)
);

CKINVDCx14_ASAP7_75t_R g1228 ( 
.A(n_1148),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1155),
.A2(n_1066),
.B1(n_1082),
.B2(n_1079),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1163),
.B(n_1188),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1144),
.A2(n_1006),
.B1(n_1017),
.B2(n_1010),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1144),
.A2(n_1006),
.B1(n_1120),
.B2(n_941),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_1141),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1124),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1156),
.B(n_1079),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1163),
.A2(n_1082),
.B1(n_1100),
.B2(n_1046),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1169),
.A2(n_1175),
.B1(n_1185),
.B2(n_1156),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1129),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1185),
.B(n_989),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

BUFx8_ASAP7_75t_L g1241 ( 
.A(n_1146),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_SL g1242 ( 
.A(n_1146),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1188),
.A2(n_1006),
.B1(n_1120),
.B2(n_1100),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1172),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_1107),
.B1(n_1009),
.B2(n_1014),
.Y(n_1245)
);

INVx5_ASAP7_75t_L g1246 ( 
.A(n_1160),
.Y(n_1246)
);

BUFx12f_ASAP7_75t_L g1247 ( 
.A(n_1172),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1135),
.B(n_1023),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1152),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1142),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1139),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1160),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1182),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1160),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1126),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1160),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1139),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1159),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1142),
.A2(n_1187),
.B1(n_1046),
.B2(n_972),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1239),
.B(n_1173),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1213),
.A2(n_1187),
.B1(n_1019),
.B2(n_1119),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1246),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1191),
.A2(n_1187),
.B1(n_1166),
.B2(n_1033),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1199),
.A2(n_1198),
.B(n_1222),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1194),
.Y(n_1265)
);

OAI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1199),
.A2(n_1198),
.B(n_1202),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1190),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1212),
.A2(n_1030),
.B1(n_989),
.B2(n_1113),
.Y(n_1268)
);

BUFx4f_ASAP7_75t_SL g1269 ( 
.A(n_1225),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1195),
.B(n_1112),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1200),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1210),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1221),
.A2(n_1195),
.B1(n_1236),
.B2(n_1229),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1211),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1203),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1219),
.A2(n_1119),
.B1(n_1030),
.B2(n_1034),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1197),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1217),
.A2(n_1027),
.B(n_795),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1193),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1223),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1221),
.A2(n_1033),
.B1(n_681),
.B2(n_1161),
.Y(n_1281)
);

BUFx4f_ASAP7_75t_SL g1282 ( 
.A(n_1241),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1224),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1230),
.B(n_1112),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1214),
.A2(n_1119),
.B1(n_1034),
.B2(n_942),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_SL g1286 ( 
.A1(n_1215),
.A2(n_1150),
.B(n_1143),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1227),
.A2(n_1161),
.B1(n_1035),
.B2(n_1002),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1250),
.B(n_945),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1259),
.A2(n_1140),
.B1(n_1150),
.B2(n_1143),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1248),
.A2(n_1035),
.B(n_975),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1228),
.A2(n_1102),
.B1(n_1113),
.B2(n_945),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1234),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1250),
.A2(n_1140),
.B1(n_1150),
.B2(n_1143),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1220),
.A2(n_1002),
.B1(n_1029),
.B2(n_1004),
.Y(n_1294)
);

OAI222xp33_ASAP7_75t_L g1295 ( 
.A1(n_1243),
.A2(n_945),
.B1(n_1102),
.B2(n_975),
.C1(n_967),
.C2(n_1000),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1237),
.A2(n_1119),
.B1(n_942),
.B2(n_960),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1238),
.A2(n_1004),
.B1(n_1031),
.B2(n_1029),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1235),
.A2(n_1193),
.B1(n_1242),
.B2(n_1218),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1240),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1205),
.A2(n_1102),
.B1(n_1255),
.B2(n_1196),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1249),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1192),
.A2(n_1000),
.B(n_1031),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1251),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1233),
.B(n_1173),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1206),
.B(n_945),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1201),
.B(n_1172),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1257),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1242),
.A2(n_960),
.B1(n_1182),
.B2(n_1026),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1205),
.A2(n_1162),
.B1(n_738),
.B2(n_1113),
.Y(n_1309)
);

INVx5_ASAP7_75t_SL g1310 ( 
.A(n_1256),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1258),
.B(n_1173),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1231),
.A2(n_1086),
.B(n_1028),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1253),
.A2(n_1245),
.B(n_1232),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1204),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1208),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1241),
.B(n_1172),
.Y(n_1316)
);

BUFx12f_ASAP7_75t_L g1317 ( 
.A(n_1207),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1192),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1208),
.B(n_1172),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1216),
.A2(n_738),
.B1(n_1182),
.B2(n_1056),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1204),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_SL g1322 ( 
.A(n_1216),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1256),
.A2(n_997),
.B(n_984),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1246),
.A2(n_1048),
.B1(n_1162),
.B2(n_1179),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1256),
.A2(n_1036),
.B1(n_1040),
.B2(n_664),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1226),
.A2(n_1036),
.B1(n_1040),
.B2(n_664),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1246),
.A2(n_1162),
.B1(n_972),
.B2(n_1170),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1226),
.A2(n_1162),
.B1(n_972),
.B2(n_1170),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1209),
.A2(n_1026),
.B(n_1024),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1252),
.Y(n_1330)
);

OAI221xp5_ASAP7_75t_L g1331 ( 
.A1(n_1281),
.A2(n_1086),
.B1(n_1024),
.B2(n_716),
.C(n_1020),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1318),
.B(n_1179),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1281),
.A2(n_1162),
.B1(n_1254),
.B2(n_1252),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1264),
.A2(n_587),
.B1(n_609),
.B2(n_1244),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1266),
.A2(n_609),
.B1(n_1247),
.B2(n_972),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1273),
.A2(n_972),
.B1(n_991),
.B2(n_986),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1263),
.A2(n_1268),
.B1(n_1308),
.B2(n_1298),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1300),
.A2(n_1209),
.B1(n_1254),
.B2(n_972),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1280),
.B(n_1209),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1267),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1263),
.B(n_1168),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1306),
.B(n_1168),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1276),
.A2(n_1284),
.B1(n_1290),
.B2(n_1270),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1261),
.A2(n_972),
.B1(n_995),
.B2(n_991),
.Y(n_1344)
);

OAI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1278),
.A2(n_995),
.B1(n_1145),
.B2(n_1037),
.C(n_467),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1318),
.A2(n_1183),
.B1(n_1044),
.B2(n_985),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1271),
.B(n_1180),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_R g1348 ( 
.A(n_1275),
.B(n_1174),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1272),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1302),
.A2(n_1183),
.B1(n_1044),
.B2(n_985),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1291),
.A2(n_1044),
.B1(n_985),
.B2(n_1180),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1274),
.B(n_1107),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1265),
.B(n_1184),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1282),
.A2(n_1044),
.B1(n_1145),
.B2(n_1165),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1260),
.A2(n_616),
.B1(n_1076),
.B2(n_473),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1282),
.A2(n_1322),
.B1(n_1315),
.B2(n_1269),
.Y(n_1356)
);

AOI222xp33_ASAP7_75t_L g1357 ( 
.A1(n_1322),
.A2(n_444),
.B1(n_452),
.B2(n_457),
.C1(n_461),
.C2(n_719),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1260),
.A2(n_616),
.B1(n_1076),
.B2(n_1174),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1283),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1324),
.B(n_1165),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1286),
.A2(n_1320),
.B1(n_1309),
.B2(n_1328),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1279),
.A2(n_1076),
.B1(n_1174),
.B2(n_1184),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1313),
.B(n_664),
.C(n_654),
.Y(n_1363)
);

AND2x2_ASAP7_75t_SL g1364 ( 
.A(n_1326),
.B(n_1164),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1329),
.A2(n_1288),
.B1(n_1305),
.B2(n_1289),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1293),
.A2(n_1076),
.B1(n_1174),
.B2(n_1184),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1317),
.A2(n_1174),
.B1(n_1005),
.B2(n_959),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_736),
.B2(n_697),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1294),
.A2(n_1095),
.B1(n_736),
.B2(n_697),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1320),
.A2(n_1145),
.B1(n_1164),
.B2(n_1165),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1269),
.A2(n_1165),
.B1(n_1164),
.B2(n_1151),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1292),
.A2(n_1151),
.B1(n_1149),
.B2(n_1122),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1285),
.A2(n_708),
.B1(n_726),
.B2(n_723),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1287),
.A2(n_1189),
.B1(n_1069),
.B2(n_1125),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1277),
.B(n_1122),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1287),
.A2(n_1189),
.B1(n_1069),
.B2(n_1125),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1296),
.A2(n_708),
.B1(n_726),
.B2(n_723),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1297),
.A2(n_708),
.B1(n_726),
.B2(n_723),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1312),
.A2(n_1122),
.B1(n_1151),
.B2(n_1149),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1297),
.A2(n_697),
.B1(n_736),
.B2(n_694),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1304),
.A2(n_694),
.B1(n_1111),
.B2(n_1133),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1319),
.A2(n_1151),
.B1(n_1149),
.B2(n_1122),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1262),
.A2(n_1151),
.B1(n_1149),
.B2(n_1122),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1316),
.A2(n_1327),
.B1(n_1324),
.B2(n_1301),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1307),
.A2(n_694),
.B1(n_1111),
.B2(n_1133),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1330),
.A2(n_1133),
.B1(n_1128),
.B2(n_1125),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1311),
.A2(n_1128),
.B1(n_1189),
.B2(n_1149),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1262),
.A2(n_1128),
.B1(n_963),
.B2(n_688),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1326),
.A2(n_1325),
.B1(n_1323),
.B2(n_1330),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1303),
.A2(n_955),
.B1(n_963),
.B2(n_978),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1299),
.B(n_963),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1310),
.A2(n_693),
.B1(n_706),
.B2(n_719),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1314),
.A2(n_955),
.B1(n_978),
.B2(n_982),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1321),
.A2(n_955),
.B1(n_978),
.B2(n_982),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1325),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1310),
.B(n_69),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1310),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1295),
.A2(n_974),
.B1(n_955),
.B2(n_978),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1266),
.B(n_70),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1264),
.A2(n_955),
.B1(n_978),
.B2(n_594),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1332),
.B(n_73),
.Y(n_1401)
);

OAI21xp33_ASAP7_75t_L g1402 ( 
.A1(n_1399),
.A2(n_1357),
.B(n_1361),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1332),
.B(n_73),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1347),
.B(n_74),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1347),
.B(n_74),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1357),
.B(n_706),
.C(n_693),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1340),
.B(n_75),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1363),
.B(n_706),
.C(n_693),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1342),
.B(n_76),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1340),
.B(n_76),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1349),
.B(n_77),
.Y(n_1411)
);

OAI221xp5_ASAP7_75t_L g1412 ( 
.A1(n_1343),
.A2(n_719),
.B1(n_718),
.B2(n_80),
.C(n_81),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1345),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.C(n_82),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1335),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.C(n_84),
.Y(n_1414)
);

AOI211xp5_ASAP7_75t_L g1415 ( 
.A1(n_1337),
.A2(n_84),
.B(n_88),
.C(n_89),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1349),
.B(n_90),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1359),
.B(n_91),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1359),
.B(n_91),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1341),
.B(n_92),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1365),
.B(n_92),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1351),
.A2(n_718),
.B1(n_642),
.B2(n_638),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1395),
.B(n_95),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_95),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1363),
.B(n_625),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1384),
.A2(n_718),
.B1(n_642),
.B2(n_638),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1356),
.A2(n_96),
.B(n_97),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1339),
.B(n_98),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1379),
.B(n_98),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1387),
.B(n_1360),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1360),
.B(n_625),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1353),
.B(n_99),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_SL g1432 ( 
.A1(n_1338),
.A2(n_99),
.B(n_642),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1352),
.B(n_631),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1334),
.A2(n_638),
.B(n_631),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1397),
.B(n_631),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1397),
.B(n_108),
.Y(n_1436)
);

NAND4xp25_ASAP7_75t_SL g1437 ( 
.A(n_1396),
.B(n_1392),
.C(n_1367),
.D(n_1336),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1396),
.B(n_112),
.Y(n_1438)
);

OR2x2_ASAP7_75t_SL g1439 ( 
.A(n_1352),
.B(n_1348),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1375),
.B(n_113),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1364),
.B(n_1389),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1364),
.B(n_115),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1364),
.B(n_116),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1350),
.A2(n_627),
.B1(n_622),
.B2(n_604),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1391),
.B(n_118),
.Y(n_1445)
);

NAND4xp25_ASAP7_75t_L g1446 ( 
.A(n_1346),
.B(n_1333),
.C(n_1331),
.D(n_1400),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1372),
.A2(n_594),
.B(n_121),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1370),
.B(n_120),
.Y(n_1448)
);

NAND4xp25_ASAP7_75t_L g1449 ( 
.A(n_1366),
.B(n_122),
.C(n_123),
.D(n_124),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1372),
.B(n_128),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1355),
.B(n_627),
.C(n_622),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1415),
.B(n_1402),
.C(n_1413),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_L g1453 ( 
.A(n_1429),
.B(n_1398),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1414),
.A2(n_1377),
.B1(n_1344),
.B2(n_1380),
.C(n_1378),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1406),
.A2(n_1374),
.B1(n_1376),
.B2(n_1358),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1381),
.C(n_1362),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1404),
.B(n_1390),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1433),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1429),
.B(n_1441),
.Y(n_1459)
);

OA211x2_ASAP7_75t_L g1460 ( 
.A1(n_1430),
.A2(n_1424),
.B(n_1437),
.C(n_1448),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_L g1461 ( 
.A(n_1426),
.B(n_1451),
.C(n_1420),
.Y(n_1461)
);

NOR3xp33_ASAP7_75t_L g1462 ( 
.A(n_1432),
.B(n_1371),
.C(n_1354),
.Y(n_1462)
);

OAI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1425),
.A2(n_1369),
.B(n_1368),
.C(n_1382),
.Y(n_1463)
);

OR2x2_ASAP7_75t_SL g1464 ( 
.A(n_1419),
.B(n_1383),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1431),
.B(n_1385),
.C(n_1388),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1433),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1386),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1407),
.Y(n_1468)
);

NAND4xp25_ASAP7_75t_L g1469 ( 
.A(n_1423),
.B(n_1373),
.C(n_1394),
.D(n_1393),
.Y(n_1469)
);

NAND4xp75_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_129),
.C(n_131),
.D(n_133),
.Y(n_1470)
);

AO21x2_ASAP7_75t_L g1471 ( 
.A1(n_1430),
.A2(n_594),
.B(n_143),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1405),
.B(n_135),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1427),
.B(n_144),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1422),
.B(n_1407),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1417),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1422),
.B(n_145),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1401),
.B(n_147),
.Y(n_1477)
);

NOR3xp33_ASAP7_75t_L g1478 ( 
.A(n_1434),
.B(n_149),
.C(n_150),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1410),
.B(n_152),
.Y(n_1479)
);

AOI211xp5_ASAP7_75t_L g1480 ( 
.A1(n_1428),
.A2(n_153),
.B(n_155),
.C(n_158),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1401),
.B(n_159),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1439),
.B(n_1403),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1409),
.B(n_627),
.C(n_622),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1468),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1482),
.B(n_1442),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1475),
.B(n_1442),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1403),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1466),
.Y(n_1488)
);

XOR2x2_ASAP7_75t_L g1489 ( 
.A(n_1452),
.B(n_1438),
.Y(n_1489)
);

NAND4xp75_ASAP7_75t_L g1490 ( 
.A(n_1460),
.B(n_1443),
.C(n_1450),
.D(n_1417),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1474),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1474),
.B(n_1443),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1459),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1418),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1453),
.B(n_1418),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1457),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1461),
.A2(n_1449),
.B1(n_1446),
.B2(n_1450),
.Y(n_1497)
);

XNOR2xp5_ASAP7_75t_L g1498 ( 
.A(n_1464),
.B(n_1477),
.Y(n_1498)
);

NAND4xp75_ASAP7_75t_L g1499 ( 
.A(n_1479),
.B(n_1473),
.C(n_1454),
.D(n_1476),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1472),
.B(n_1436),
.Y(n_1501)
);

NAND4xp75_ASAP7_75t_L g1502 ( 
.A(n_1454),
.B(n_1424),
.C(n_1447),
.D(n_1411),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1481),
.B(n_1447),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1455),
.B(n_1447),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1483),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1471),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1408),
.B1(n_1421),
.B2(n_1445),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1471),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1480),
.B(n_1416),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1488),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1488),
.Y(n_1511)
);

XOR2x2_ASAP7_75t_L g1512 ( 
.A(n_1489),
.B(n_1470),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1484),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1496),
.Y(n_1514)
);

XNOR2x2_ASAP7_75t_L g1515 ( 
.A(n_1499),
.B(n_1465),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1491),
.Y(n_1516)
);

XOR2x2_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1456),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_R g1518 ( 
.A(n_1509),
.B(n_1435),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1486),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1495),
.Y(n_1520)
);

XOR2x2_ASAP7_75t_L g1521 ( 
.A(n_1498),
.B(n_1478),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1487),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1498),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1500),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1493),
.Y(n_1525)
);

XOR2x2_ASAP7_75t_L g1526 ( 
.A(n_1499),
.B(n_1440),
.Y(n_1526)
);

XNOR2x1_ASAP7_75t_L g1527 ( 
.A(n_1497),
.B(n_1444),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1504),
.B(n_1505),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1485),
.B(n_1463),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1492),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1486),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1494),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1492),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1485),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1503),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

AOI22x1_ASAP7_75t_L g1537 ( 
.A1(n_1515),
.A2(n_1504),
.B1(n_1506),
.B2(n_1503),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1534),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1528),
.A2(n_1509),
.B1(n_1508),
.B2(n_1501),
.Y(n_1539)
);

OAI22x1_ASAP7_75t_L g1540 ( 
.A1(n_1528),
.A2(n_1508),
.B1(n_1507),
.B2(n_1490),
.Y(n_1540)
);

XOR2x2_ASAP7_75t_L g1541 ( 
.A(n_1517),
.B(n_1502),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1523),
.Y(n_1542)
);

AOI22x1_ASAP7_75t_L g1543 ( 
.A1(n_1515),
.A2(n_1512),
.B1(n_1529),
.B2(n_1517),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1514),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1513),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1524),
.B(n_1502),
.Y(n_1546)
);

OA22x2_ASAP7_75t_L g1547 ( 
.A1(n_1512),
.A2(n_1463),
.B1(n_1469),
.B2(n_165),
.Y(n_1547)
);

XOR2x2_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_160),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1525),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1526),
.A2(n_594),
.B1(n_604),
.B2(n_595),
.Y(n_1550)
);

OAI22x1_ASAP7_75t_SL g1551 ( 
.A1(n_1523),
.A2(n_604),
.B1(n_595),
.B2(n_172),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1534),
.Y(n_1552)
);

AOI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1520),
.A2(n_1521),
.B1(n_1526),
.B2(n_1530),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1532),
.Y(n_1554)
);

AOI22x1_ASAP7_75t_L g1555 ( 
.A1(n_1533),
.A2(n_161),
.B1(n_169),
.B2(n_173),
.Y(n_1555)
);

OA22x2_ASAP7_75t_L g1556 ( 
.A1(n_1519),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_1556)
);

OAI322xp33_ASAP7_75t_L g1557 ( 
.A1(n_1543),
.A2(n_1527),
.A3(n_1535),
.B1(n_1516),
.B2(n_1522),
.C1(n_1519),
.C2(n_1531),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1549),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1536),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

AOI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1541),
.A2(n_1527),
.B1(n_1513),
.B2(n_1511),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1538),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1544),
.Y(n_1563)
);

XOR2x2_ASAP7_75t_L g1564 ( 
.A(n_1541),
.B(n_1518),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1554),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1542),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1538),
.Y(n_1567)
);

INVxp33_ASAP7_75t_SL g1568 ( 
.A(n_1542),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1554),
.Y(n_1569)
);

NOR4xp25_ASAP7_75t_L g1570 ( 
.A(n_1557),
.B(n_1546),
.C(n_1548),
.D(n_1553),
.Y(n_1570)
);

AND4x1_ASAP7_75t_L g1571 ( 
.A(n_1561),
.B(n_1550),
.C(n_1546),
.D(n_1548),
.Y(n_1571)
);

AOI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1569),
.A2(n_1539),
.B1(n_1540),
.B2(n_1551),
.C(n_1537),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1566),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1564),
.A2(n_1547),
.B1(n_1552),
.B2(n_1556),
.Y(n_1574)
);

OA22x2_ASAP7_75t_L g1575 ( 
.A1(n_1569),
.A2(n_1545),
.B1(n_1547),
.B2(n_1511),
.Y(n_1575)
);

OA22x2_ASAP7_75t_L g1576 ( 
.A1(n_1565),
.A2(n_1545),
.B1(n_1510),
.B2(n_1556),
.Y(n_1576)
);

OA22x2_ASAP7_75t_L g1577 ( 
.A1(n_1562),
.A2(n_1510),
.B1(n_1555),
.B2(n_192),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1573),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1575),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1574),
.A2(n_1568),
.B1(n_1567),
.B2(n_1563),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1572),
.A2(n_1568),
.B1(n_1558),
.B2(n_1559),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1577),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_SL g1584 ( 
.A1(n_1570),
.A2(n_1560),
.B(n_1559),
.C(n_194),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1578),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1581),
.A2(n_1560),
.B1(n_1571),
.B2(n_595),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1582),
.Y(n_1587)
);

NOR4xp25_ASAP7_75t_L g1588 ( 
.A(n_1584),
.B(n_184),
.C(n_187),
.D(n_195),
.Y(n_1588)
);

AO22x2_ASAP7_75t_L g1589 ( 
.A1(n_1580),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1579),
.A2(n_1583),
.B1(n_216),
.B2(n_217),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1582),
.B(n_212),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1587),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1585),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1589),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1586),
.A2(n_1588),
.B1(n_1590),
.B2(n_1591),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1585),
.Y(n_1596)
);

AND4x1_ASAP7_75t_L g1597 ( 
.A(n_1595),
.B(n_236),
.C(n_237),
.D(n_239),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1594),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1596),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1593),
.Y(n_1600)
);

AOI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1592),
.A2(n_240),
.B(n_241),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1601),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1600),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1599),
.B(n_245),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1597),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1598),
.B(n_252),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1605),
.Y(n_1607)
);

OAI22x1_ASAP7_75t_L g1608 ( 
.A1(n_1602),
.A2(n_257),
.B1(n_258),
.B2(n_264),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1603),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1606),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1606),
.A2(n_269),
.B1(n_270),
.B2(n_275),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1609),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1607),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1610),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1610),
.Y(n_1615)
);

OA22x2_ASAP7_75t_L g1616 ( 
.A1(n_1613),
.A2(n_1608),
.B1(n_1611),
.B2(n_1604),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1614),
.A2(n_278),
.B1(n_281),
.B2(n_282),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1615),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_1618)
);

AO22x2_ASAP7_75t_L g1619 ( 
.A1(n_1612),
.A2(n_289),
.B1(n_292),
.B2(n_296),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1616),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1619),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1620),
.A2(n_1618),
.B1(n_1617),
.B2(n_302),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1621),
.A2(n_297),
.B1(n_300),
.B2(n_305),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1622),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1624),
.A2(n_1623),
.B1(n_316),
.B2(n_318),
.C(n_325),
.Y(n_1625)
);

AOI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1625),
.A2(n_330),
.B(n_331),
.C(n_333),
.Y(n_1626)
);


endmodule