module fake_jpeg_11027_n_84 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_32),
.B1(n_34),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_38),
.B1(n_34),
.B2(n_3),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_58),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_37),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_61),
.Y(n_72)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_28),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_13),
.Y(n_61)
);

AOI22x1_ASAP7_75t_R g62 ( 
.A1(n_43),
.A2(n_38),
.B1(n_14),
.B2(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_2),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_1),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_5),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_75),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_55),
.C(n_19),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_72),
.A3(n_69),
.B1(n_65),
.B2(n_71),
.C(n_64),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_74),
.A3(n_75),
.B1(n_7),
.B2(n_8),
.C1(n_11),
.C2(n_9),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_78),
.C(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_8),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_20),
.Y(n_84)
);


endmodule