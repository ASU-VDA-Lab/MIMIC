module fake_netlist_1_8675_n_1208 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1208);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1208;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_1198;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_1202;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_1196;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_1175;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_1177;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_1185;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1197;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_1200;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1201;
wire n_1191;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_1194;
wire n_694;
wire n_301;
wire n_1179;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1174;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1078;
wire n_1016;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_1204;
wire n_652;
wire n_975;
wire n_279;
wire n_303;
wire n_968;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_1183;
wire n_567;
wire n_809;
wire n_888;
wire n_1188;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1159;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_1132;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_1180;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1160;
wire n_1184;
wire n_274;
wire n_1018;
wire n_1195;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_735;
wire n_696;
wire n_1091;
wire n_1203;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_1186;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_990;
wire n_751;
wire n_800;
wire n_626;
wire n_941;
wire n_1147;
wire n_1206;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_1178;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_1176;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_1181;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_1199;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_1193;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_1125;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1069;
wire n_1021;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_1189;
wire n_923;
wire n_1205;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1117;
wire n_859;
wire n_1027;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_1182;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_1207;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_1187;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_1190;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_1192;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_88), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_218), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_120), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_90), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_157), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_134), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_40), .B(n_196), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_236), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_234), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_60), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_71), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_183), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_226), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_238), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_245), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_86), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_251), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_69), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_102), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_71), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_47), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_55), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_165), .Y(n_281) );
BUFx2_ASAP7_75t_SL g282 ( .A(n_172), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_223), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_248), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_253), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_131), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_13), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_69), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_214), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_125), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_145), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_133), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_114), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_142), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_205), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_159), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_88), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_138), .Y(n_300) );
BUFx10_ASAP7_75t_L g301 ( .A(n_93), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_204), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_8), .B(n_32), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_113), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_126), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_154), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_100), .Y(n_307) );
CKINVDCx16_ASAP7_75t_R g308 ( .A(n_174), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_52), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_86), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_175), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_106), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_83), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_13), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_42), .Y(n_316) );
CKINVDCx16_ASAP7_75t_R g317 ( .A(n_38), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_220), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_0), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_189), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_135), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_180), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_118), .Y(n_324) );
INVxp33_ASAP7_75t_SL g325 ( .A(n_122), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_107), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_31), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_7), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_173), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_85), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_48), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_124), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_132), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_184), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_79), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_101), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_19), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_74), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_121), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_182), .Y(n_340) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_80), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_249), .Y(n_342) );
BUFx2_ASAP7_75t_SL g343 ( .A(n_244), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_139), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_168), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_31), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_169), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_190), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_68), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_240), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_44), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_105), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_232), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_77), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_111), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_49), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_176), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_195), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_14), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_109), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_237), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_64), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_194), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_123), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_30), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_73), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_243), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_115), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_61), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_197), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_21), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_36), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_23), .B(n_18), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_78), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_187), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_170), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_127), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_59), .Y(n_378) );
BUFx8_ASAP7_75t_SL g379 ( .A(n_150), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_91), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_11), .Y(n_381) );
CKINVDCx16_ASAP7_75t_R g382 ( .A(n_211), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_221), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_23), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_200), .Y(n_385) );
BUFx8_ASAP7_75t_SL g386 ( .A(n_144), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_3), .Y(n_387) );
INVxp33_ASAP7_75t_SL g388 ( .A(n_202), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_80), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_239), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_116), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_0), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_79), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_20), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_48), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_128), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_50), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_312), .B(n_1), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_316), .Y(n_399) );
OAI22x1_ASAP7_75t_SL g400 ( .A1(n_397), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_316), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_267), .A2(n_99), .B(n_98), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_316), .B(n_2), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_269), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_389), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_379), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_277), .Y(n_407) );
CKINVDCx6p67_ASAP7_75t_R g408 ( .A(n_266), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_389), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_392), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_273), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_277), .Y(n_413) );
NOR2xp33_ASAP7_75t_SL g414 ( .A(n_308), .B(n_254), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_277), .Y(n_415) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_283), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_283), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_339), .B(n_4), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_269), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_344), .B(n_4), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_283), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_257), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_259), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_279), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_317), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_283), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_385), .B(n_5), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_332), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_260), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_332), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_261), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_262), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_332), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_354), .B(n_5), .Y(n_435) );
BUFx8_ASAP7_75t_L g436 ( .A(n_332), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_345), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_267), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_415), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_415), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_415), .Y(n_441) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_403), .B(n_355), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_406), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_415), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_435), .A2(n_278), .B1(n_280), .B2(n_274), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_403), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_435), .A2(n_299), .B1(n_309), .B2(n_288), .Y(n_447) );
AOI21x1_ASAP7_75t_L g448 ( .A1(n_403), .A2(n_307), .B(n_272), .Y(n_448) );
INVx4_ASAP7_75t_L g449 ( .A(n_403), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_436), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_420), .B(n_382), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_438), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_408), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_420), .B(n_256), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_423), .B(n_256), .Y(n_458) );
NAND2xp33_ASAP7_75t_L g459 ( .A(n_423), .B(n_424), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_412), .Y(n_460) );
NAND2xp33_ASAP7_75t_R g461 ( .A(n_402), .B(n_325), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_425), .B(n_301), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_415), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_408), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_399), .Y(n_465) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_415), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_424), .B(n_285), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_399), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
AND2x6_ASAP7_75t_L g471 ( .A(n_435), .B(n_273), .Y(n_471) );
BUFx4f_ASAP7_75t_L g472 ( .A(n_402), .Y(n_472) );
NAND2xp33_ASAP7_75t_L g473 ( .A(n_430), .B(n_275), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_401), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_430), .B(n_285), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_401), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_438), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_432), .B(n_297), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
AOI21x1_ASAP7_75t_L g480 ( .A1(n_407), .A2(n_307), .B(n_272), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_432), .B(n_377), .Y(n_481) );
BUFx4f_ASAP7_75t_L g482 ( .A(n_402), .Y(n_482) );
OAI22x1_ASAP7_75t_L g483 ( .A1(n_425), .A2(n_268), .B1(n_276), .B2(n_255), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_414), .A2(n_341), .B1(n_284), .B2(n_292), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
INVx6_ASAP7_75t_L g486 ( .A(n_436), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_433), .B(n_255), .Y(n_487) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_442), .B(n_414), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_462), .B(n_398), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_443), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_453), .B(n_398), .Y(n_491) );
NAND2xp33_ASAP7_75t_L g492 ( .A(n_471), .B(n_286), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_487), .B(n_419), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_478), .B(n_419), .Y(n_494) );
BUFx2_ASAP7_75t_L g495 ( .A(n_453), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_472), .A2(n_402), .B(n_433), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_481), .B(n_421), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_465), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_484), .B(n_428), .C(n_421), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_465), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_449), .B(n_428), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_462), .B(n_452), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_449), .B(n_412), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_442), .B(n_404), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_442), .A2(n_471), .B1(n_459), .B2(n_447), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_L g507 ( .A1(n_472), .A2(n_404), .B(n_294), .C(n_291), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_456), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_449), .B(n_404), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_449), .B(n_263), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
INVx3_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_454), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_471), .B(n_322), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_484), .A2(n_271), .B1(n_292), .B2(n_284), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_469), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_458), .B(n_325), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_456), .Y(n_518) );
NOR2x2_ASAP7_75t_L g519 ( .A(n_464), .B(n_426), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_471), .B(n_396), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_446), .B(n_264), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_446), .B(n_270), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_480), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_451), .B(n_281), .Y(n_524) );
NAND2xp33_ASAP7_75t_L g525 ( .A(n_471), .B(n_396), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_474), .Y(n_526) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_483), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_451), .A2(n_331), .B1(n_394), .B2(n_258), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_472), .B(n_290), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_450), .A2(n_331), .B1(n_394), .B2(n_258), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_455), .Y(n_532) );
NAND3xp33_ASAP7_75t_SL g533 ( .A(n_445), .B(n_304), .C(n_271), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_467), .B(n_388), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_457), .A2(n_321), .B1(n_324), .B2(n_304), .Y(n_535) );
NAND3xp33_ASAP7_75t_SL g536 ( .A(n_475), .B(n_324), .C(n_321), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_455), .B(n_405), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_476), .A2(n_409), .B1(n_411), .B2(n_405), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_455), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_473), .A2(n_329), .B1(n_350), .B2(n_326), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_476), .B(n_409), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_454), .B(n_268), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_480), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_468), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_479), .B(n_411), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_479), .B(n_417), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_486), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_486), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_472), .A2(n_310), .B1(n_319), .B2(n_315), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_468), .B(n_287), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_470), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_470), .B(n_293), .Y(n_552) );
BUFx3_ASAP7_75t_L g553 ( .A(n_486), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_482), .A2(n_326), .B1(n_350), .B2(n_329), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_482), .A2(n_402), .B(n_383), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_448), .B(n_353), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_470), .B(n_318), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_460), .Y(n_558) );
AO22x1_ASAP7_75t_L g559 ( .A1(n_477), .A2(n_276), .B1(n_395), .B2(n_327), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_477), .B(n_303), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_485), .A2(n_373), .B(n_337), .C(n_338), .Y(n_561) );
INVx8_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_485), .B(n_327), .Y(n_563) );
OA22x2_ASAP7_75t_L g564 ( .A1(n_461), .A2(n_400), .B1(n_395), .B2(n_335), .Y(n_564) );
NOR2x1p5_ASAP7_75t_L g565 ( .A(n_448), .B(n_400), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_486), .B(n_340), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_439), .B(n_295), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_439), .A2(n_367), .B1(n_375), .B2(n_361), .Y(n_568) );
AND2x6_ASAP7_75t_SL g569 ( .A(n_466), .B(n_365), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_439), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_440), .B(n_296), .Y(n_571) );
AND3x1_ASAP7_75t_L g572 ( .A(n_440), .B(n_359), .C(n_371), .Y(n_572) );
AO32x1_ASAP7_75t_L g573 ( .A1(n_523), .A2(n_410), .A3(n_418), .B1(n_413), .B2(n_407), .Y(n_573) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_495), .B(n_289), .Y(n_574) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
BUFx2_ASAP7_75t_L g576 ( .A(n_508), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_490), .Y(n_577) );
AO22x1_ASAP7_75t_L g578 ( .A1(n_554), .A2(n_379), .B1(n_386), .B2(n_397), .Y(n_578) );
A2O1A1Ixp33_ASAP7_75t_L g579 ( .A1(n_499), .A2(n_359), .B(n_374), .C(n_372), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_503), .B(n_301), .Y(n_580) );
OR2x6_ASAP7_75t_SL g581 ( .A(n_519), .B(n_314), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_494), .B(n_328), .Y(n_582) );
INVx4_ASAP7_75t_L g583 ( .A(n_562), .Y(n_583) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_497), .A2(n_444), .B(n_441), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_488), .A2(n_367), .B1(n_375), .B2(n_361), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_498), .B(n_330), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_555), .A2(n_507), .B(n_556), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_489), .B(n_301), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_501), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_493), .B(n_346), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_488), .A2(n_506), .B1(n_500), .B2(n_549), .Y(n_591) );
INVxp67_ASAP7_75t_L g592 ( .A(n_518), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_491), .B(n_351), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_530), .A2(n_463), .B(n_300), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_549), .A2(n_381), .B(n_378), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_562), .Y(n_596) );
OR2x6_ASAP7_75t_L g597 ( .A(n_565), .B(n_282), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_491), .B(n_349), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_502), .A2(n_463), .B(n_306), .Y(n_599) );
NOR2xp33_ASAP7_75t_SL g600 ( .A(n_515), .B(n_386), .Y(n_600) );
INVx2_ASAP7_75t_SL g601 ( .A(n_563), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_560), .B(n_356), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_561), .A2(n_380), .B(n_393), .C(n_384), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_541), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_533), .B(n_366), .C(n_362), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_560), .B(n_369), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_510), .A2(n_313), .B(n_298), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_542), .B(n_387), .Y(n_608) );
NOR2x1_ASAP7_75t_R g609 ( .A(n_527), .B(n_343), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_517), .B(n_302), .Y(n_610) );
AOI21x1_ASAP7_75t_L g611 ( .A1(n_543), .A2(n_323), .B(n_320), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_569), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_556), .A2(n_334), .B(n_333), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_504), .A2(n_342), .B(n_336), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_509), .A2(n_348), .B(n_347), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_505), .A2(n_360), .B(n_363), .C(n_358), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_526), .A2(n_364), .B(n_376), .C(n_368), .Y(n_618) );
OR2x6_ASAP7_75t_SL g619 ( .A(n_515), .B(n_352), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_536), .B(n_265), .C(n_305), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_559), .B(n_357), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_528), .Y(n_622) );
BUFx8_ASAP7_75t_L g623 ( .A(n_531), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_534), .B(n_390), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_545), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_521), .A2(n_383), .B(n_370), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_568), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_546), .Y(n_628) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_548), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_6), .Y(n_630) );
AOI21xp5_ASAP7_75t_L g631 ( .A1(n_522), .A2(n_524), .B(n_543), .Y(n_631) );
BUFx12f_ASAP7_75t_L g632 ( .A(n_544), .Y(n_632) );
AND2x6_ASAP7_75t_L g633 ( .A(n_553), .B(n_311), .Y(n_633) );
INVx4_ASAP7_75t_L g634 ( .A(n_548), .Y(n_634) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_540), .B(n_391), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_547), .B(n_6), .Y(n_636) );
INVx5_ASAP7_75t_L g637 ( .A(n_511), .Y(n_637) );
OAI22x1_ASAP7_75t_L g638 ( .A1(n_535), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_532), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_539), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_564), .A2(n_345), .B1(n_410), .B2(n_407), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_514), .B(n_10), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_572), .B(n_410), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_520), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_512), .Y(n_645) );
INVx3_ASAP7_75t_SL g646 ( .A(n_564), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_492), .B(n_429), .C(n_422), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_513), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_513), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_551), .A2(n_434), .B(n_437), .C(n_429), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_538), .B(n_11), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g652 ( .A1(n_538), .A2(n_434), .B(n_416), .C(n_427), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_525), .B(n_12), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_550), .A2(n_466), .B(n_416), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_552), .A2(n_466), .B(n_416), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_557), .B(n_14), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_566), .B(n_15), .C(n_16), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_558), .B(n_15), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_567), .B(n_17), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_571), .B(n_17), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_571), .B(n_18), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_570), .B(n_19), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_497), .A2(n_416), .B(n_415), .Y(n_663) );
AO21x1_ASAP7_75t_L g664 ( .A1(n_555), .A2(n_427), .B(n_416), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_562), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_497), .A2(n_466), .B(n_427), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_497), .A2(n_466), .B(n_427), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_494), .B(n_21), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_497), .A2(n_427), .B(n_416), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_488), .A2(n_427), .B1(n_431), .B2(n_416), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_494), .B(n_22), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_497), .A2(n_431), .B(n_103), .Y(n_672) );
AOI21x1_ASAP7_75t_L g673 ( .A1(n_497), .A2(n_431), .B(n_104), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_537), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_491), .B(n_24), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_499), .Y(n_676) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_562), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_497), .A2(n_431), .B(n_108), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_508), .B(n_25), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_488), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_680) );
INVx3_ASAP7_75t_SL g681 ( .A(n_519), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_503), .B(n_26), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_496), .B(n_27), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_497), .A2(n_112), .B(n_110), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_577), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_682), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_627), .B(n_28), .Y(n_687) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_579), .A2(n_29), .B(n_30), .C(n_32), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_574), .B(n_29), .Y(n_689) );
OAI22x1_ASAP7_75t_L g690 ( .A1(n_681), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_601), .B(n_33), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_604), .B(n_35), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_603), .A2(n_36), .B1(n_37), .B2(n_38), .C(n_39), .Y(n_693) );
BUFx3_ASAP7_75t_L g694 ( .A(n_632), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_631), .A2(n_119), .B(n_117), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_575), .B(n_37), .Y(n_696) );
OR2x2_ASAP7_75t_L g697 ( .A(n_582), .B(n_39), .Y(n_697) );
NOR2xp33_ASAP7_75t_SL g698 ( .A(n_600), .B(n_40), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_591), .A2(n_41), .B(n_43), .C(n_44), .Y(n_699) );
AND2x6_ASAP7_75t_L g700 ( .A(n_575), .B(n_41), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_591), .A2(n_43), .B(n_45), .C(n_46), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_587), .A2(n_130), .B(n_129), .Y(n_702) );
AO31x2_ASAP7_75t_L g703 ( .A1(n_670), .A2(n_46), .A3(n_47), .B(n_49), .Y(n_703) );
AOI221xp5_ASAP7_75t_SL g704 ( .A1(n_617), .A2(n_50), .B1(n_51), .B2(n_52), .C(n_53), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_602), .B(n_51), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_618), .A2(n_53), .B(n_54), .C(n_55), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_668), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_575), .B(n_54), .Y(n_708) );
OR2x6_ASAP7_75t_L g709 ( .A(n_578), .B(n_56), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_669), .A2(n_137), .B(n_136), .Y(n_710) );
AOI221x1_ASAP7_75t_L g711 ( .A1(n_672), .A2(n_678), .B1(n_680), .B2(n_657), .C(n_684), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_671), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_588), .B(n_56), .Y(n_713) );
O2A1O1Ixp33_ASAP7_75t_L g714 ( .A1(n_630), .A2(n_57), .B(n_58), .C(n_61), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_608), .A2(n_57), .B(n_58), .C(n_62), .Y(n_715) );
AO31x2_ASAP7_75t_L g716 ( .A1(n_652), .A2(n_62), .A3(n_63), .B(n_64), .Y(n_716) );
CKINVDCx6p67_ASAP7_75t_R g717 ( .A(n_581), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_654), .A2(n_141), .B(n_140), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_655), .A2(n_179), .B(n_250), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_586), .B(n_63), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_619), .B(n_65), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_593), .B(n_65), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_585), .A2(n_66), .B1(n_67), .B2(n_70), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_605), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_593), .B(n_72), .Y(n_725) );
AND2x2_ASAP7_75t_SL g726 ( .A(n_636), .B(n_75), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_606), .B(n_75), .Y(n_727) );
CKINVDCx8_ASAP7_75t_R g728 ( .A(n_597), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_595), .A2(n_76), .B(n_77), .C(n_78), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_614), .A2(n_186), .B(n_247), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_625), .A2(n_181), .B(n_246), .Y(n_731) );
BUFx2_ASAP7_75t_SL g732 ( .A(n_636), .Y(n_732) );
AO31x2_ASAP7_75t_L g733 ( .A1(n_650), .A2(n_76), .A3(n_81), .B(n_82), .Y(n_733) );
NOR2x1_ASAP7_75t_SL g734 ( .A(n_583), .B(n_81), .Y(n_734) );
BUFx12f_ASAP7_75t_L g735 ( .A(n_623), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_576), .B(n_82), .Y(n_736) );
AO21x1_ASAP7_75t_L g737 ( .A1(n_643), .A2(n_191), .B(n_242), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g738 ( .A1(n_628), .A2(n_83), .B(n_84), .C(n_85), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_613), .A2(n_178), .B(n_241), .Y(n_739) );
AO31x2_ASAP7_75t_L g740 ( .A1(n_638), .A2(n_84), .A3(n_87), .B(n_89), .Y(n_740) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_596), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_592), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_616), .A2(n_87), .B(n_89), .C(n_90), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g744 ( .A(n_583), .B(n_91), .Y(n_744) );
AOI211x1_ASAP7_75t_L g745 ( .A1(n_651), .A2(n_92), .B(n_93), .C(n_94), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_679), .Y(n_746) );
INVx6_ASAP7_75t_SL g747 ( .A(n_597), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_622), .A2(n_192), .B(n_233), .Y(n_748) );
AO31x2_ASAP7_75t_L g749 ( .A1(n_626), .A2(n_92), .A3(n_95), .B(n_96), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_589), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_646), .Y(n_751) );
INVx4_ASAP7_75t_L g752 ( .A(n_596), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_679), .B(n_95), .Y(n_753) );
OAI21xp33_ASAP7_75t_L g754 ( .A1(n_590), .A2(n_96), .B(n_97), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_599), .A2(n_193), .B(n_143), .Y(n_755) );
INVx3_ASAP7_75t_L g756 ( .A(n_596), .Y(n_756) );
AND2x4_ASAP7_75t_L g757 ( .A(n_674), .B(n_649), .Y(n_757) );
A2O1A1Ixp33_ASAP7_75t_L g758 ( .A1(n_676), .A2(n_97), .B(n_146), .C(n_147), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_580), .B(n_148), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g760 ( .A(n_620), .B(n_149), .C(n_151), .Y(n_760) );
BUFx12f_ASAP7_75t_L g761 ( .A(n_635), .Y(n_761) );
AOI221x1_ASAP7_75t_L g762 ( .A1(n_647), .A2(n_152), .B1(n_153), .B2(n_155), .C(n_156), .Y(n_762) );
INVxp67_ASAP7_75t_SL g763 ( .A(n_665), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_641), .Y(n_764) );
BUFx10_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_594), .A2(n_158), .B(n_160), .Y(n_766) );
CKINVDCx6p67_ASAP7_75t_R g767 ( .A(n_637), .Y(n_767) );
AOI221x1_ASAP7_75t_L g768 ( .A1(n_653), .A2(n_161), .B1(n_162), .B2(n_163), .C(n_164), .Y(n_768) );
AO21x1_ASAP7_75t_L g769 ( .A1(n_683), .A2(n_166), .B(n_167), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_642), .A2(n_171), .B(n_198), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_639), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_660), .A2(n_199), .B(n_203), .C(n_206), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_637), .B(n_207), .Y(n_773) );
AOI31xp67_ASAP7_75t_L g774 ( .A1(n_573), .A2(n_208), .A3(n_209), .B(n_210), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_598), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_624), .B(n_212), .Y(n_776) );
INVx6_ASAP7_75t_SL g777 ( .A(n_624), .Y(n_777) );
AND2x6_ASAP7_75t_L g778 ( .A(n_665), .B(n_213), .Y(n_778) );
BUFx4f_ASAP7_75t_SL g779 ( .A(n_665), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_640), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_658), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_573), .A2(n_216), .B(n_217), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_610), .B(n_219), .Y(n_783) );
BUFx2_ASAP7_75t_L g784 ( .A(n_633), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g785 ( .A1(n_615), .A2(n_222), .B(n_224), .C(n_227), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_677), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_621), .B(n_228), .Y(n_787) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_677), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_656), .B(n_229), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_659), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_607), .A2(n_230), .B(n_231), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_661), .Y(n_792) );
BUFx12f_ASAP7_75t_L g793 ( .A(n_633), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_645), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_662), .Y(n_795) );
BUFx8_ASAP7_75t_L g796 ( .A(n_633), .Y(n_796) );
AO31x2_ASAP7_75t_L g797 ( .A1(n_573), .A2(n_634), .A3(n_644), .B(n_648), .Y(n_797) );
BUFx10_ASAP7_75t_L g798 ( .A(n_629), .Y(n_798) );
AO31x2_ASAP7_75t_L g799 ( .A1(n_609), .A2(n_664), .A3(n_670), .B(n_555), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_591), .A2(n_617), .B(n_604), .C(n_595), .Y(n_800) );
AO31x2_ASAP7_75t_L g801 ( .A1(n_664), .A2(n_670), .A3(n_555), .B(n_497), .Y(n_801) );
OAI22x1_ASAP7_75t_L g802 ( .A1(n_681), .A2(n_484), .B1(n_540), .B2(n_568), .Y(n_802) );
BUFx3_ASAP7_75t_L g803 ( .A(n_577), .Y(n_803) );
NOR2xp33_ASAP7_75t_SL g804 ( .A(n_681), .B(n_554), .Y(n_804) );
AND3x2_ASAP7_75t_L g805 ( .A(n_600), .B(n_453), .C(n_612), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_604), .B(n_494), .Y(n_806) );
AOI21x1_ASAP7_75t_L g807 ( .A1(n_584), .A2(n_673), .B(n_611), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_591), .A2(n_488), .B1(n_506), .B2(n_604), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_631), .A2(n_497), .B(n_507), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_574), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_682), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_682), .Y(n_812) );
AO31x2_ASAP7_75t_L g813 ( .A1(n_664), .A2(n_670), .A3(n_555), .B(n_497), .Y(n_813) );
BUFx12f_ASAP7_75t_L g814 ( .A(n_623), .Y(n_814) );
OAI21xp5_ASAP7_75t_L g815 ( .A1(n_631), .A2(n_497), .B(n_507), .Y(n_815) );
OAI21x1_ASAP7_75t_L g816 ( .A1(n_584), .A2(n_663), .B(n_666), .Y(n_816) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_575), .Y(n_817) );
NOR2x1_ASAP7_75t_SL g818 ( .A(n_583), .B(n_575), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g819 ( .A1(n_631), .A2(n_497), .B(n_507), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g820 ( .A1(n_809), .A2(n_819), .B(n_815), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_806), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_750), .Y(n_822) );
BUFx2_ASAP7_75t_L g823 ( .A(n_810), .Y(n_823) );
INVx2_ASAP7_75t_SL g824 ( .A(n_779), .Y(n_824) );
OR2x6_ASAP7_75t_L g825 ( .A(n_753), .B(n_732), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_753), .A2(n_808), .B1(n_800), .B2(n_726), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_802), .A2(n_777), .B1(n_804), .B2(n_747), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_777), .Y(n_828) );
NAND2x1p5_ASAP7_75t_L g829 ( .A(n_694), .B(n_803), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_692), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_796), .Y(n_831) );
OA21x2_ASAP7_75t_L g832 ( .A1(n_816), .A2(n_711), .B(n_807), .Y(n_832) );
INVx2_ASAP7_75t_SL g833 ( .A(n_767), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_744), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_736), .B(n_721), .Y(n_835) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_707), .A2(n_727), .B(n_705), .C(n_715), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_790), .B(n_792), .Y(n_837) );
INVx3_ASAP7_75t_SL g838 ( .A(n_717), .Y(n_838) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_736), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_691), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_775), .B(n_713), .Y(n_841) );
INVxp33_ASAP7_75t_L g842 ( .A(n_742), .Y(n_842) );
AO31x2_ASAP7_75t_L g843 ( .A1(n_768), .A2(n_762), .A3(n_737), .B(n_769), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_771), .Y(n_844) );
AO31x2_ASAP7_75t_L g845 ( .A1(n_782), .A2(n_699), .A3(n_701), .B(n_729), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_698), .A2(n_723), .B1(n_687), .B2(n_764), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_747), .A2(n_795), .B1(n_709), .B2(n_746), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_689), .B(n_757), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_722), .Y(n_849) );
INVx4_ASAP7_75t_L g850 ( .A(n_793), .Y(n_850) );
OR2x2_ASAP7_75t_L g851 ( .A(n_685), .B(n_725), .Y(n_851) );
AND2x4_ASAP7_75t_L g852 ( .A(n_757), .B(n_818), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_709), .B(n_686), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_734), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_811), .B(n_812), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_781), .B(n_697), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_720), .B(n_759), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_780), .Y(n_858) );
HB1xp67_ASAP7_75t_L g859 ( .A(n_786), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_745), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g861 ( .A(n_704), .B(n_760), .C(n_738), .Y(n_861) );
AO31x2_ASAP7_75t_L g862 ( .A1(n_702), .A2(n_758), .A3(n_772), .B(n_695), .Y(n_862) );
OAI21xp5_ASAP7_75t_L g863 ( .A1(n_730), .A2(n_743), .B(n_770), .Y(n_863) );
BUFx8_ASAP7_75t_L g864 ( .A(n_735), .Y(n_864) );
BUFx2_ASAP7_75t_R g865 ( .A(n_728), .Y(n_865) );
AO31x2_ASAP7_75t_L g866 ( .A1(n_785), .A2(n_710), .A3(n_718), .B(n_719), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_794), .B(n_776), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g868 ( .A1(n_706), .A2(n_688), .B(n_731), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_749), .Y(n_869) );
INVx6_ASAP7_75t_L g870 ( .A(n_814), .Y(n_870) );
BUFx3_ASAP7_75t_L g871 ( .A(n_751), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_755), .A2(n_714), .B(n_789), .Y(n_872) );
AOI21xp5_ASAP7_75t_SL g873 ( .A1(n_773), .A2(n_784), .B(n_791), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_783), .A2(n_754), .B(n_787), .C(n_724), .Y(n_874) );
OA21x2_ASAP7_75t_L g875 ( .A1(n_739), .A2(n_748), .B(n_766), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_703), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_752), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_703), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_741), .B(n_817), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_761), .A2(n_765), .B1(n_805), .B2(n_693), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_700), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_700), .Y(n_882) );
INVx4_ASAP7_75t_SL g883 ( .A(n_700), .Y(n_883) );
AOI21xp33_ASAP7_75t_SL g884 ( .A1(n_690), .A2(n_696), .B(n_708), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_797), .Y(n_885) );
CKINVDCx11_ASAP7_75t_R g886 ( .A(n_741), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_797), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_700), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_733), .Y(n_889) );
AO31x2_ASAP7_75t_L g890 ( .A1(n_801), .A2(n_813), .A3(n_774), .B(n_799), .Y(n_890) );
CKINVDCx6p67_ASAP7_75t_R g891 ( .A(n_778), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_799), .B(n_813), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_733), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_799), .B(n_756), .Y(n_894) );
AND2x4_ASAP7_75t_L g895 ( .A(n_788), .B(n_763), .Y(n_895) );
AOI22xp5_ASAP7_75t_SL g896 ( .A1(n_778), .A2(n_740), .B1(n_716), .B2(n_798), .Y(n_896) );
AND2x4_ASAP7_75t_L g897 ( .A(n_797), .B(n_716), .Y(n_897) );
AO31x2_ASAP7_75t_L g898 ( .A1(n_716), .A2(n_664), .A3(n_711), .B(n_808), .Y(n_898) );
BUFx3_ASAP7_75t_L g899 ( .A(n_803), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_806), .B(n_604), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_806), .B(n_604), .Y(n_901) );
INVx4_ASAP7_75t_L g902 ( .A(n_779), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_806), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_806), .B(n_726), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_806), .B(n_489), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_806), .B(n_503), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_806), .B(n_726), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_809), .A2(n_667), .B(n_666), .Y(n_908) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_804), .B(n_515), .Y(n_909) );
OAI21xp5_ASAP7_75t_L g910 ( .A1(n_800), .A2(n_587), .B(n_497), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_806), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_806), .B(n_604), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_806), .Y(n_913) );
NAND3xp33_ASAP7_75t_L g914 ( .A(n_711), .B(n_745), .C(n_704), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_806), .Y(n_915) );
A2O1A1Ixp33_ASAP7_75t_L g916 ( .A1(n_707), .A2(n_591), .B(n_712), .C(n_800), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_806), .Y(n_917) );
INVx2_ASAP7_75t_SL g918 ( .A(n_779), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_806), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_806), .Y(n_920) );
OAI21xp5_ASAP7_75t_L g921 ( .A1(n_800), .A2(n_587), .B(n_497), .Y(n_921) );
AO31x2_ASAP7_75t_L g922 ( .A1(n_711), .A2(n_664), .A3(n_808), .B(n_768), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_806), .B(n_726), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_804), .B(n_515), .Y(n_924) );
BUFx2_ASAP7_75t_L g925 ( .A(n_810), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_806), .Y(n_926) );
AO21x1_ASAP7_75t_L g927 ( .A1(n_808), .A2(n_680), .B(n_715), .Y(n_927) );
OAI21xp33_ASAP7_75t_SL g928 ( .A1(n_753), .A2(n_488), .B(n_591), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_806), .B(n_604), .Y(n_929) );
OR2x2_ASAP7_75t_L g930 ( .A(n_806), .B(n_489), .Y(n_930) );
NOR2xp33_ASAP7_75t_SL g931 ( .A(n_796), .B(n_793), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_806), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_806), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_913), .B(n_919), .Y(n_934) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_920), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_886), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_926), .B(n_826), .Y(n_937) );
OR2x6_ASAP7_75t_L g938 ( .A(n_873), .B(n_826), .Y(n_938) );
AO21x2_ASAP7_75t_L g939 ( .A1(n_910), .A2(n_921), .B(n_820), .Y(n_939) );
AND2x4_ASAP7_75t_L g940 ( .A(n_883), .B(n_881), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_869), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_876), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_928), .A2(n_904), .B1(n_907), .B2(n_923), .Y(n_943) );
INVx5_ASAP7_75t_L g944 ( .A(n_825), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_821), .B(n_903), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_911), .B(n_915), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_878), .Y(n_947) );
AND2x4_ASAP7_75t_L g948 ( .A(n_882), .B(n_888), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_879), .B(n_894), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_917), .B(n_932), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_889), .Y(n_951) );
AO21x2_ASAP7_75t_L g952 ( .A1(n_914), .A2(n_892), .B(n_908), .Y(n_952) );
BUFx2_ASAP7_75t_L g953 ( .A(n_928), .Y(n_953) );
NAND4xp25_ASAP7_75t_L g954 ( .A(n_909), .B(n_924), .C(n_827), .D(n_847), .Y(n_954) );
INVx3_ASAP7_75t_L g955 ( .A(n_891), .Y(n_955) );
OAI21xp5_ASAP7_75t_L g956 ( .A1(n_861), .A2(n_836), .B(n_874), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_893), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_860), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_933), .B(n_905), .Y(n_959) );
INVx5_ASAP7_75t_L g960 ( .A(n_825), .Y(n_960) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_823), .Y(n_961) );
OA21x2_ASAP7_75t_L g962 ( .A1(n_885), .A2(n_887), .B(n_897), .Y(n_962) );
BUFx3_ASAP7_75t_L g963 ( .A(n_852), .Y(n_963) );
HB1xp67_ASAP7_75t_L g964 ( .A(n_925), .Y(n_964) );
INVxp67_ASAP7_75t_SL g965 ( .A(n_900), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_837), .Y(n_966) );
INVx4_ASAP7_75t_L g967 ( .A(n_852), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_837), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_930), .B(n_906), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_822), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_916), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_844), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_858), .Y(n_973) );
OR2x6_ASAP7_75t_L g974 ( .A(n_825), .B(n_854), .Y(n_974) );
INVxp67_ASAP7_75t_SL g975 ( .A(n_901), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_901), .B(n_912), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_896), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_832), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_896), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_912), .B(n_929), .Y(n_980) );
INVxp67_ASAP7_75t_L g981 ( .A(n_929), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_890), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_856), .B(n_841), .Y(n_983) );
OR2x2_ASAP7_75t_L g984 ( .A(n_856), .B(n_859), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_890), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g986 ( .A1(n_868), .A2(n_846), .B(n_872), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_890), .Y(n_987) );
OR2x2_ASAP7_75t_SL g988 ( .A(n_870), .B(n_839), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_857), .B(n_840), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_855), .B(n_830), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_898), .Y(n_991) );
INVx4_ASAP7_75t_R g992 ( .A(n_824), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_849), .B(n_835), .Y(n_993) );
INVx2_ASAP7_75t_SL g994 ( .A(n_833), .Y(n_994) );
BUFx3_ASAP7_75t_L g995 ( .A(n_899), .Y(n_995) );
INVx3_ASAP7_75t_L g996 ( .A(n_877), .Y(n_996) );
BUFx2_ASAP7_75t_L g997 ( .A(n_895), .Y(n_997) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_846), .B(n_884), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_922), .Y(n_999) );
AO21x2_ASAP7_75t_L g1000 ( .A1(n_863), .A2(n_868), .B(n_872), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_848), .B(n_877), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1002 ( .A(n_842), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_884), .A2(n_857), .B1(n_853), .B2(n_880), .C(n_834), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_867), .B(n_851), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_922), .Y(n_1005) );
OA21x2_ASAP7_75t_L g1006 ( .A1(n_927), .A2(n_922), .B(n_867), .Y(n_1006) );
BUFx2_ASAP7_75t_L g1007 ( .A(n_828), .Y(n_1007) );
INVx2_ASAP7_75t_L g1008 ( .A(n_845), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_976), .B(n_831), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_976), .B(n_871), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_965), .B(n_845), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_953), .B(n_843), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_980), .A2(n_931), .B1(n_870), .B2(n_838), .Y(n_1013) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_975), .B(n_829), .Y(n_1014) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_935), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_980), .B(n_918), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_949), .B(n_986), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_978), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_969), .B(n_865), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_945), .B(n_902), .Y(n_1020) );
OAI21xp5_ASAP7_75t_SL g1021 ( .A1(n_943), .A2(n_931), .B(n_864), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_949), .B(n_862), .Y(n_1022) );
INVxp67_ASAP7_75t_L g1023 ( .A(n_961), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1024 ( .A(n_949), .B(n_866), .Y(n_1024) );
BUFx2_ASAP7_75t_L g1025 ( .A(n_938), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_942), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_945), .B(n_902), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_937), .B(n_850), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_946), .B(n_850), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_946), .B(n_864), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_942), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_947), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_948), .B(n_875), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_948), .B(n_940), .Y(n_1034) );
AND2x4_ASAP7_75t_L g1035 ( .A(n_977), .B(n_979), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g1036 ( .A(n_959), .B(n_954), .Y(n_1036) );
OR2x2_ASAP7_75t_L g1037 ( .A(n_984), .B(n_981), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1038 ( .A(n_979), .B(n_951), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_954), .A2(n_998), .B1(n_1003), .B2(n_993), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_950), .B(n_990), .Y(n_1040) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_995), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1042 ( .A(n_984), .Y(n_1042) );
INVx3_ASAP7_75t_L g1043 ( .A(n_962), .Y(n_1043) );
BUFx2_ASAP7_75t_L g1044 ( .A(n_997), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_983), .B(n_966), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_941), .B(n_1006), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1006), .B(n_939), .Y(n_1047) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_995), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1006), .B(n_939), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1006), .B(n_939), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_957), .B(n_970), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_970), .B(n_966), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_968), .B(n_972), .Y(n_1053) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_968), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1004), .B(n_989), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_982), .Y(n_1056) );
OR2x2_ASAP7_75t_L g1057 ( .A(n_1004), .B(n_989), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_972), .B(n_973), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1059 ( .A1(n_944), .A2(n_960), .B1(n_988), .B2(n_967), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_973), .B(n_1000), .Y(n_1060) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_963), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1018), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_1054), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1017), .B(n_952), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1017), .B(n_952), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1060), .B(n_952), .Y(n_1066) );
NAND2xp5_ASAP7_75t_SL g1067 ( .A(n_1059), .B(n_944), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1042), .B(n_958), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_1018), .Y(n_1069) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_1015), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1052), .B(n_958), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1060), .B(n_962), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1052), .B(n_934), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1056), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1022), .B(n_962), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1040), .B(n_964), .Y(n_1076) );
OR2x2_ASAP7_75t_L g1077 ( .A(n_1055), .B(n_1008), .Y(n_1077) );
INVx3_ASAP7_75t_L g1078 ( .A(n_1043), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1045), .B(n_1002), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1046), .B(n_1000), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1037), .B(n_971), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1046), .B(n_1000), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1055), .B(n_985), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1051), .B(n_1005), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1057), .B(n_997), .Y(n_1085) );
AND2x2_ASAP7_75t_SL g1086 ( .A(n_1025), .B(n_967), .Y(n_1086) );
INVx4_ASAP7_75t_L g1087 ( .A(n_1061), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1026), .Y(n_1088) );
INVx1_ASAP7_75t_SL g1089 ( .A(n_1041), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_1057), .B(n_987), .Y(n_1090) );
INVx1_ASAP7_75t_SL g1091 ( .A(n_1041), .Y(n_1091) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_1044), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_1036), .B(n_1001), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1051), .B(n_1005), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1026), .Y(n_1095) );
AND2x4_ASAP7_75t_SL g1096 ( .A(n_1034), .B(n_967), .Y(n_1096) );
BUFx2_ASAP7_75t_L g1097 ( .A(n_1044), .Y(n_1097) );
OR2x2_ASAP7_75t_L g1098 ( .A(n_1035), .B(n_999), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1012), .B(n_991), .Y(n_1099) );
INVxp67_ASAP7_75t_SL g1100 ( .A(n_1043), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1031), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1053), .B(n_1001), .Y(n_1102) );
NAND4xp25_ASAP7_75t_L g1103 ( .A(n_1039), .B(n_956), .C(n_1007), .D(n_955), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1032), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1032), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1062), .Y(n_1106) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1075), .B(n_1033), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1070), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1080), .B(n_1024), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1080), .B(n_1024), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1082), .B(n_1024), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1082), .B(n_1047), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1071), .B(n_1058), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1088), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_1083), .B(n_1011), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1088), .Y(n_1116) );
NAND2x1p5_ASAP7_75t_L g1117 ( .A(n_1086), .B(n_944), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1095), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1064), .B(n_1047), .Y(n_1119) );
INVx4_ASAP7_75t_L g1120 ( .A(n_1096), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1101), .Y(n_1121) );
AND2x4_ASAP7_75t_SL g1122 ( .A(n_1087), .B(n_1034), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1084), .B(n_1058), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1090), .B(n_1038), .Y(n_1124) );
INVx3_ASAP7_75t_L g1125 ( .A(n_1078), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1065), .B(n_1049), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_1065), .B(n_1050), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1101), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1075), .B(n_1050), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1062), .Y(n_1130) );
INVxp67_ASAP7_75t_L g1131 ( .A(n_1089), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1084), .B(n_1038), .Y(n_1132) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1069), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1104), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1105), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1074), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1077), .B(n_1038), .Y(n_1137) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1077), .B(n_1038), .Y(n_1138) );
NOR2xp33_ASAP7_75t_L g1139 ( .A(n_1093), .B(n_1030), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1131), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1141 ( .A(n_1112), .B(n_1066), .Y(n_1141) );
INVx3_ASAP7_75t_L g1142 ( .A(n_1120), .Y(n_1142) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1106), .Y(n_1143) );
NOR2xp33_ASAP7_75t_L g1144 ( .A(n_1108), .B(n_936), .Y(n_1144) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1106), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1114), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1114), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1112), .B(n_1094), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_1120), .A2(n_1021), .B1(n_1103), .B2(n_1013), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_1107), .B(n_1078), .Y(n_1150) );
OR2x2_ASAP7_75t_L g1151 ( .A(n_1119), .B(n_1072), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1129), .B(n_1072), .Y(n_1152) );
CKINVDCx5p33_ASAP7_75t_R g1153 ( .A(n_1139), .Y(n_1153) );
OAI32xp33_ASAP7_75t_L g1154 ( .A1(n_1117), .A2(n_1091), .A3(n_1103), .B1(n_1014), .B2(n_1048), .Y(n_1154) );
INVx1_ASAP7_75t_SL g1155 ( .A(n_1122), .Y(n_1155) );
OR2x2_ASAP7_75t_L g1156 ( .A(n_1126), .B(n_1098), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1126), .B(n_1094), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1127), .B(n_1099), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_1123), .B(n_1048), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1116), .Y(n_1160) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1130), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1133), .Y(n_1162) );
NAND2x1_ASAP7_75t_SL g1163 ( .A(n_1142), .B(n_1087), .Y(n_1163) );
AOI31xp33_ASAP7_75t_L g1164 ( .A1(n_1149), .A2(n_1117), .A3(n_1067), .B(n_1028), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1140), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1149), .B(n_1023), .C(n_1079), .Y(n_1166) );
NOR2xp33_ASAP7_75t_L g1167 ( .A(n_1153), .B(n_994), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1168 ( .A1(n_1154), .A2(n_1122), .B(n_1086), .Y(n_1168) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1144), .B(n_1076), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1143), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1143), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1151), .B(n_1127), .Y(n_1172) );
NAND2xp5_ASAP7_75t_SL g1173 ( .A(n_1155), .B(n_1087), .Y(n_1173) );
OAI21xp5_ASAP7_75t_L g1174 ( .A1(n_1154), .A2(n_1063), .B(n_1029), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1145), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1156), .Y(n_1176) );
OAI22xp33_ASAP7_75t_SL g1177 ( .A1(n_1173), .A2(n_1151), .B1(n_1150), .B2(n_1159), .Y(n_1177) );
NAND3xp33_ASAP7_75t_L g1178 ( .A(n_1166), .B(n_1019), .C(n_1010), .Y(n_1178) );
OAI21xp33_ASAP7_75t_L g1179 ( .A1(n_1164), .A2(n_1141), .B(n_1148), .Y(n_1179) );
OAI321xp33_ASAP7_75t_L g1180 ( .A1(n_1174), .A2(n_1115), .A3(n_1124), .B1(n_1132), .B2(n_1138), .C(n_1137), .Y(n_1180) );
INVxp67_ASAP7_75t_L g1181 ( .A(n_1165), .Y(n_1181) );
AOI21xp5_ASAP7_75t_L g1182 ( .A1(n_1168), .A2(n_1096), .B(n_1157), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_1167), .A2(n_1009), .B1(n_1020), .B2(n_1027), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1176), .B(n_1152), .Y(n_1184) );
OR3x1_ASAP7_75t_L g1185 ( .A(n_1163), .B(n_1147), .C(n_1146), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1186 ( .A1(n_1169), .A2(n_1158), .B1(n_1068), .B2(n_1110), .C(n_1111), .Y(n_1186) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_1172), .A2(n_1158), .B1(n_1110), .B2(n_1111), .C(n_1109), .Y(n_1187) );
AOI322xp5_ASAP7_75t_L g1188 ( .A1(n_1170), .A2(n_1113), .A3(n_1102), .B1(n_1016), .B2(n_1085), .C1(n_1160), .C2(n_1081), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_1171), .A2(n_1092), .B1(n_1097), .B2(n_1135), .C(n_1136), .Y(n_1189) );
AOI21xp5_ASAP7_75t_L g1190 ( .A1(n_1171), .A2(n_1096), .B(n_1100), .Y(n_1190) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1181), .B(n_1179), .Y(n_1191) );
AOI221xp5_ASAP7_75t_L g1192 ( .A1(n_1180), .A2(n_1177), .B1(n_1178), .B2(n_1182), .C(n_1186), .Y(n_1192) );
AND4x1_ASAP7_75t_L g1193 ( .A(n_1183), .B(n_1187), .C(n_1190), .D(n_1189), .Y(n_1193) );
NAND3xp33_ASAP7_75t_SL g1194 ( .A(n_1188), .B(n_1185), .C(n_1183), .Y(n_1194) );
INVxp67_ASAP7_75t_L g1195 ( .A(n_1191), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1193), .Y(n_1196) );
NOR2x1_ASAP7_75t_L g1197 ( .A(n_1194), .B(n_992), .Y(n_1197) );
NAND3xp33_ASAP7_75t_SL g1198 ( .A(n_1196), .B(n_1192), .C(n_992), .Y(n_1198) );
AND3x1_ASAP7_75t_L g1199 ( .A(n_1197), .B(n_1184), .C(n_1175), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1195), .B(n_1175), .Y(n_1200) );
INVx2_ASAP7_75t_SL g1201 ( .A(n_1200), .Y(n_1201) );
XNOR2x1_ASAP7_75t_L g1202 ( .A(n_1199), .B(n_974), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1201), .B(n_1198), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_1203), .A2(n_1202), .B1(n_960), .B2(n_974), .Y(n_1204) );
AOI222xp33_ASAP7_75t_L g1205 ( .A1(n_1204), .A2(n_1092), .B1(n_1125), .B2(n_996), .C1(n_1116), .C2(n_1118), .Y(n_1205) );
OA21x2_ASAP7_75t_L g1206 ( .A1(n_1205), .A2(n_1128), .B(n_1134), .Y(n_1206) );
AOI21xp5_ASAP7_75t_L g1207 ( .A1(n_1206), .A2(n_1073), .B(n_1121), .Y(n_1207) );
AOI21xp5_ASAP7_75t_L g1208 ( .A1(n_1207), .A2(n_1162), .B(n_1161), .Y(n_1208) );
endmodule