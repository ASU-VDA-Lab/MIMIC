module fake_jpeg_21361_n_319 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_13),
.B1(n_19),
.B2(n_21),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_13),
.B1(n_19),
.B2(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_13),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_19),
.B(n_15),
.C(n_11),
.Y(n_60)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_13),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_51),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_19),
.B1(n_37),
.B2(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_19),
.B1(n_29),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_37),
.B1(n_29),
.B2(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_61),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_67),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_72),
.B(n_48),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_45),
.B1(n_41),
.B2(n_44),
.Y(n_85)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_54),
.B1(n_36),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_44),
.B1(n_40),
.B2(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_56),
.B1(n_55),
.B2(n_58),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_88),
.B(n_99),
.C(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_48),
.C(n_58),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_27),
.C(n_26),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_95),
.B(n_17),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_44),
.B1(n_40),
.B2(n_45),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_64),
.B1(n_76),
.B2(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_71),
.A2(n_40),
.B1(n_43),
.B2(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_61),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_65),
.B1(n_78),
.B2(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_102),
.B1(n_95),
.B2(n_96),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_63),
.B1(n_64),
.B2(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_107),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_116),
.C(n_27),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_105),
.A2(n_124),
.B1(n_22),
.B2(n_15),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_70),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_94),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_81),
.C(n_80),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_16),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_108),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_74),
.B1(n_30),
.B2(n_46),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_35),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_74),
.B1(n_18),
.B2(n_21),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_74),
.B1(n_18),
.B2(n_21),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_123),
.B(n_15),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_27),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_126),
.A2(n_147),
.B1(n_11),
.B2(n_32),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_14),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_154),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_150),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_141),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_82),
.B1(n_98),
.B2(n_22),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_138),
.B1(n_118),
.B2(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_117),
.B(n_101),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_155),
.B(n_11),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_36),
.B1(n_22),
.B2(n_50),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_21),
.B1(n_18),
.B2(n_36),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_153),
.B1(n_35),
.B2(n_17),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_21),
.B1(n_22),
.B2(n_36),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_152),
.C(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_32),
.C(n_26),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_15),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_12),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_14),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_124),
.B(n_120),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_156),
.B(n_129),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_112),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_167),
.B(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_168),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_126),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_130),
.B(n_124),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_173),
.C(n_152),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_182),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_124),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_124),
.C(n_118),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_119),
.B1(n_22),
.B2(n_11),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_129),
.B1(n_147),
.B2(n_128),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_176),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_140),
.Y(n_207)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_146),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_155),
.B1(n_144),
.B2(n_145),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_177),
.B1(n_175),
.B2(n_12),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_192),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_200),
.C(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_197),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_14),
.B1(n_12),
.B2(n_16),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_133),
.C(n_139),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_140),
.B(n_150),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_208),
.B(n_180),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_209),
.B1(n_163),
.B2(n_167),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_154),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_185),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_206),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_23),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_23),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_168),
.B1(n_161),
.B2(n_180),
.Y(n_215)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_159),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_176),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_188),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_236),
.B1(n_17),
.B2(n_23),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_178),
.C(n_186),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_222),
.C(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_163),
.B1(n_164),
.B2(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_187),
.C(n_159),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_177),
.C(n_24),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_35),
.C(n_28),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_209),
.C(n_194),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_16),
.B1(n_17),
.B2(n_35),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_232),
.A2(n_199),
.B1(n_208),
.B2(n_207),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_219),
.B1(n_222),
.B2(n_220),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_17),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_201),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_250),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_210),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_246),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_211),
.C(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_230),
.C(n_231),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_202),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_198),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_234),
.A2(n_14),
.B(n_16),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_10),
.B(n_9),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_235),
.B1(n_226),
.B2(n_229),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_268),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_260),
.C(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_223),
.C(n_227),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_233),
.C(n_236),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_226),
.B1(n_17),
.B2(n_7),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_255),
.B1(n_254),
.B2(n_247),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_17),
.C(n_23),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_241),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_9),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_239),
.C(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_281),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_256),
.A2(n_243),
.B(n_246),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_2),
.B(n_3),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_265),
.C(n_266),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_249),
.C(n_17),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_249),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_264),
.B1(n_8),
.B2(n_7),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_278),
.Y(n_289)
);

AOI321xp33_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_8),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_0),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_6),
.C(n_4),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_0),
.C(n_1),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_0),
.C(n_2),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_294),
.A2(n_4),
.B(n_5),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_3),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_4),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_4),
.C(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_5),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_303),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_274),
.B(n_5),
.C(n_6),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_5),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_300),
.B(n_289),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_306),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_313),
.B(n_309),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_307),
.B(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_286),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_288),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_6),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_6),
.Y(n_319)
);


endmodule