module fake_netlist_5_892_n_150 (n_29, n_16, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_150);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_150;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_124;
wire n_86;
wire n_136;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_126;
wire n_84;
wire n_130;
wire n_79;
wire n_131;
wire n_47;
wire n_53;
wire n_44;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVxp33_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_15),
.B(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_1),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_4),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_5),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_65),
.Y(n_81)
);

OR2x6_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_7),
.B1(n_20),
.B2(n_21),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_66),
.B(n_61),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_57),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_59),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_52),
.B(n_50),
.C(n_49),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_60),
.B(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

AND2x6_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_56),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_47),
.B(n_28),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_47),
.B(n_32),
.C(n_34),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_79),
.B1(n_82),
.B2(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_82),
.B1(n_75),
.B2(n_81),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_84),
.B(n_76),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_81),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_71),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_80),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_76),
.B1(n_80),
.B2(n_36),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_106),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_100),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_98),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_93),
.B(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_97),
.Y(n_126)
);

NAND4xp25_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_92),
.C(n_102),
.D(n_37),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_121),
.B1(n_120),
.B2(n_114),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_76),
.B1(n_35),
.B2(n_40),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_27),
.B1(n_112),
.B2(n_111),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_111),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_119),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_119),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_119),
.Y(n_135)
);

OR2x6_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_127),
.B1(n_119),
.B2(n_116),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_130),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_137),
.B(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_136),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_138),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

NOR2xp67_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_144),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_138),
.B1(n_136),
.B2(n_140),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_125),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_116),
.B(n_125),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_112),
.B1(n_78),
.B2(n_148),
.Y(n_150)
);


endmodule