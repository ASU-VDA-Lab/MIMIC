module real_jpeg_4297_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_255;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_295;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_18)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_71),
.B1(n_82),
.B2(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_1),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_1),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_83),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_5),
.B(n_9),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_5),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_90),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_6),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_9),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_62),
.B(n_66),
.C(n_70),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_9),
.A2(n_56),
.B1(n_90),
.B2(n_94),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_56),
.B1(n_98),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_56),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_9),
.B(n_101),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_143),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_9),
.B(n_247),
.C(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_9),
.B(n_204),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_9),
.B(n_48),
.C(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_11),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_206),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_192),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_121),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_60),
.C(n_95),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_16),
.A2(n_95),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_16),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_16),
.A2(n_196),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_18),
.A2(n_54),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_26),
.B(n_27),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_26),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_27),
.Y(n_204)
);

AOI22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_30),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_30),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_30),
.Y(n_167)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_31),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_31),
.Y(n_245)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_46),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_54),
.B(n_190),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_60),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_61),
.A2(n_72),
.B1(n_73),
.B2(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_61),
.Y(n_216)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_101)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_72),
.A2(n_73),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_73),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_73),
.B(n_239),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_73),
.B(n_176),
.C(n_257),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_74),
.B(n_89),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_74),
.A2(n_81),
.B1(n_89),
.B2(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_80),
.Y(n_220)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_86),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx8_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_87),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_89),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_118),
.B2(n_120),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_96),
.A2(n_100),
.B1(n_118),
.B2(n_120),
.Y(n_188)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_177),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_139),
.B2(n_176),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_129),
.B1(n_130),
.B2(n_135),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_182),
.B(n_185),
.Y(n_181)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_129),
.B(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_139),
.A2(n_176),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_140),
.A2(n_141),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_164),
.B1(n_169),
.B2(n_175),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_164),
.B1(n_169),
.B2(n_175),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_142),
.A2(n_169),
.B(n_175),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.Y(n_143)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_176),
.B(n_280),
.C(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_179),
.A2(n_180),
.B1(n_243),
.B2(n_251),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_251),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_179),
.A2(n_180),
.B1(n_202),
.B2(n_213),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_179),
.B(n_202),
.C(n_264),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_202),
.C(n_205),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_187),
.A2(n_188),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.C(n_200),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_218),
.C(n_221),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_226),
.B(n_295),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_223),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_208),
.B(n_223),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_217),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_209),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_217),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_242),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_285)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_289),
.B(n_294),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_277),
.B(n_288),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_261),
.B(n_276),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_253),
.B(n_260),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_241),
.B(n_252),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_238),
.B(n_240),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_259),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_274),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_274),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_282),
.B1(n_283),
.B2(n_286),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);


endmodule