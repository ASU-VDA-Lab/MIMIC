module fake_ibex_1082_n_17 (n_1, n_4, n_3, n_6, n_5, n_2, n_0, n_17);

input n_1;
input n_4;
input n_3;
input n_6;
input n_5;
input n_2;
input n_0;

output n_17;


BUFx16f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);


endmodule