module real_jpeg_9128_n_16 (n_5, n_4, n_8, n_0, n_12, n_309, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_309;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx24_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_54),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_40),
.B1(n_50),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_2),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_104),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_104),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_104),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_4),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_155),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_4),
.A2(n_40),
.B1(n_50),
.B2(n_155),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_5),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_146),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_146),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_40),
.B1(n_50),
.B2(n_146),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_36),
.B1(n_40),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_6),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_12),
.A2(n_58),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_12),
.B(n_58),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_12),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_12),
.A2(n_27),
.B1(n_33),
.B2(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_12),
.B(n_52),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_12),
.A2(n_42),
.B(n_46),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_12),
.A2(n_40),
.B1(n_50),
.B2(n_164),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_15),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_77),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_15),
.A2(n_40),
.B1(n_50),
.B2(n_77),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_112),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_92),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_21),
.A2(n_22),
.B1(n_72),
.B2(n_73),
.Y(n_300)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_55),
.B2(n_71),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_25),
.A2(n_38),
.B(n_71),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_25),
.A2(n_26),
.B1(n_56),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_27),
.A2(n_33),
.B1(n_145),
.B2(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_27),
.A2(n_98),
.B(n_148),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_27),
.A2(n_34),
.B(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_27),
.A2(n_33),
.B1(n_211),
.B2(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_27),
.A2(n_197),
.B(n_233),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_28),
.B(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_28),
.A2(n_32),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_29),
.A2(n_30),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_29),
.B(n_65),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_29),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_30),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_32),
.B(n_97),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_33),
.B(n_164),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_33),
.A2(n_96),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_48),
.B(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_39),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_39),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_39),
.A2(n_44),
.B1(n_247),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_39),
.A2(n_44),
.B1(n_103),
.B2(n_256),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B(n_43),
.C(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_40),
.A2(n_41),
.B(n_164),
.C(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_44),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_79),
.B(n_81),
.C(n_82),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_79),
.Y(n_81)
);

HAxp5_ASAP7_75t_SL g189 ( 
.A(n_46),
.B(n_164),
.CON(n_189),
.SN(n_189)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_49),
.B(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_52),
.A2(n_120),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_56),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_66),
.B(n_68),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_64),
.B1(n_66),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_57),
.A2(n_64),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_57),
.A2(n_64),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_57),
.A2(n_64),
.B1(n_154),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_57),
.A2(n_64),
.B1(n_179),
.B2(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_57),
.A2(n_85),
.B(n_187),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_59),
.B1(n_79),
.B2(n_80),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_58),
.B(n_79),
.Y(n_195)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_59),
.A2(n_81),
.B1(n_189),
.B2(n_195),
.Y(n_194)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_64),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_64),
.A2(n_88),
.B(n_100),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_69),
.A2(n_87),
.B(n_90),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_84),
.B(n_91),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_78),
.A2(n_82),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_78),
.A2(n_127),
.B(n_259),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_82),
.B(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_114),
.B1(n_115),
.B2(n_132),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_91),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_92),
.A2(n_93),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.C(n_106),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_94),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_95),
.B(n_99),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_108),
.B(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_108),
.A2(n_124),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_108),
.A2(n_124),
.B1(n_207),
.B2(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_133),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_124),
.A2(n_243),
.B(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_284),
.A3(n_296),
.B1(n_301),
.B2(n_307),
.C(n_309),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_249),
.C(n_280),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_223),
.B(n_248),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_200),
.B(n_222),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_182),
.B(n_199),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_173),
.B(n_181),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_161),
.B(n_172),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_149),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_160),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_160),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_167),
.B(n_171),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_175),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_183),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.CI(n_180),
.CON(n_176),
.SN(n_176)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_193),
.B2(n_198),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_186),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_188),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_192),
.C(n_198),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_193),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_196),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_216),
.B2(n_217),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_219),
.C(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_215),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_212),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_218),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_237),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_236),
.C(n_237),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_232),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_244),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_241),
.C(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_267),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_267),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_261),
.C(n_265),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_254),
.C(n_260),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_260),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_267)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_276),
.C(n_277),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_285),
.A2(n_302),
.B(n_306),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_287),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_293),
.C(n_295),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B(n_305),
.Y(n_302)
);


endmodule