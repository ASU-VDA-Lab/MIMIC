module real_aes_2497_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_570;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_231;
wire n_547;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_481;
wire n_498;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_623;
wire n_249;
wire n_446;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_294;
wire n_393;
wire n_258;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_0), .A2(n_196), .B1(n_274), .B2(n_277), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_1), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_2), .A2(n_115), .B1(n_277), .B2(n_310), .Y(n_309) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_3), .A2(n_154), .B1(n_244), .B2(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g590 ( .A(n_3), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_4), .A2(n_103), .B1(n_267), .B2(n_270), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_5), .A2(n_194), .B1(n_549), .B2(n_551), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_6), .A2(n_48), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_7), .A2(n_142), .B1(n_295), .B2(n_298), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_8), .A2(n_51), .B1(n_301), .B2(n_315), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_9), .A2(n_84), .B1(n_402), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_10), .A2(n_158), .B1(n_284), .B2(n_321), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_11), .A2(n_71), .B1(n_373), .B2(n_376), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_12), .A2(n_81), .B1(n_300), .B2(n_301), .Y(n_319) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_13), .A2(n_53), .B1(n_244), .B2(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_13), .B(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_14), .A2(n_33), .B1(n_300), .B2(n_318), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_15), .A2(n_145), .B1(n_411), .B2(n_483), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_16), .A2(n_116), .B1(n_287), .B2(n_291), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_17), .A2(n_32), .B1(n_604), .B2(n_605), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_18), .A2(n_223), .B(n_230), .C(n_592), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_19), .A2(n_47), .B1(n_410), .B2(n_411), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_20), .A2(n_70), .B1(n_295), .B2(n_297), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_21), .A2(n_175), .B1(n_284), .B2(n_321), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_22), .A2(n_220), .B1(n_300), .B2(n_301), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_23), .A2(n_203), .B1(n_549), .B2(n_551), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_24), .A2(n_140), .B1(n_398), .B2(n_400), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_25), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_26), .A2(n_159), .B1(n_287), .B2(n_301), .Y(n_366) );
AOI222xp33_ASAP7_75t_L g627 ( .A1(n_27), .A2(n_110), .B1(n_221), .B2(n_395), .C1(n_400), .C2(n_568), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_28), .A2(n_210), .B1(n_300), .B2(n_301), .Y(n_352) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_29), .A2(n_38), .B1(n_520), .B2(n_521), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_30), .A2(n_169), .B1(n_404), .B2(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_31), .A2(n_212), .B1(n_614), .B2(n_616), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_34), .A2(n_86), .B1(n_413), .B2(n_416), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_35), .B(n_240), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_36), .A2(n_168), .B1(n_444), .B2(n_446), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_37), .A2(n_217), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_39), .A2(n_179), .B1(n_438), .B2(n_568), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_40), .A2(n_72), .B1(n_601), .B2(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_41), .A2(n_177), .B1(n_314), .B2(n_315), .Y(n_313) );
AO222x2_ASAP7_75t_L g343 ( .A1(n_42), .A2(n_52), .B1(n_156), .B2(n_240), .C1(n_258), .C2(n_262), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_43), .A2(n_63), .B1(n_365), .B2(n_574), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g340 ( .A(n_44), .B(n_341), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_45), .A2(n_173), .B1(n_292), .B2(n_300), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_46), .A2(n_162), .B1(n_314), .B2(n_317), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_49), .A2(n_96), .B1(n_277), .B2(n_310), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_50), .A2(n_137), .B1(n_267), .B2(n_270), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_54), .A2(n_58), .B1(n_310), .B2(n_346), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_55), .A2(n_208), .B1(n_258), .B2(n_262), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_56), .A2(n_128), .B1(n_434), .B2(n_435), .Y(n_433) );
XNOR2x2_ASAP7_75t_L g458 ( .A(n_57), .B(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_59), .A2(n_166), .B1(n_438), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_60), .A2(n_141), .B1(n_314), .B2(n_317), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_61), .B(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_62), .A2(n_138), .B1(n_481), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_64), .A2(n_191), .B1(n_291), .B2(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_65), .A2(n_111), .B1(n_513), .B2(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_66), .A2(n_87), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx3_ASAP7_75t_L g244 ( .A(n_67), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_68), .A2(n_134), .B1(n_405), .B2(n_566), .Y(n_565) );
AO22x2_ASAP7_75t_L g562 ( .A1(n_69), .A2(n_563), .B1(n_577), .B2(n_578), .Y(n_562) );
INVx1_ASAP7_75t_L g577 ( .A(n_69), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_73), .B(n_435), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_74), .A2(n_152), .B1(n_315), .B2(n_318), .Y(n_355) );
XOR2x2_ASAP7_75t_L g304 ( .A(n_75), .B(n_305), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_76), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_77), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_78), .A2(n_176), .B1(n_258), .B2(n_262), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_79), .A2(n_207), .B1(n_629), .B2(n_630), .Y(n_628) );
AO22x1_ASAP7_75t_L g461 ( .A1(n_80), .A2(n_129), .B1(n_462), .B2(n_463), .Y(n_461) );
INVx1_ASAP7_75t_SL g245 ( .A(n_82), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_82), .B(n_104), .Y(n_591) );
INVx2_ASAP7_75t_L g229 ( .A(n_83), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_85), .A2(n_190), .B1(n_379), .B2(n_381), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_88), .A2(n_122), .B1(n_479), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_89), .A2(n_178), .B1(n_483), .B2(n_485), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_90), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_91), .A2(n_102), .B1(n_317), .B2(n_318), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_92), .A2(n_107), .B1(n_501), .B2(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_93), .A2(n_101), .B1(n_301), .B2(n_546), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_94), .A2(n_183), .B1(n_410), .B2(n_411), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_95), .A2(n_112), .B1(n_553), .B2(n_556), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_97), .A2(n_113), .B1(n_404), .B2(n_632), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_98), .A2(n_205), .B1(n_267), .B2(n_270), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_99), .B(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_100), .A2(n_193), .B1(n_314), .B2(n_337), .Y(n_336) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_104), .A2(n_164), .B1(n_244), .B2(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_105), .B(n_240), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_106), .A2(n_161), .B1(n_379), .B2(n_435), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_108), .B(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_109), .A2(n_136), .B1(n_398), .B2(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_114), .A2(n_187), .B1(n_258), .B2(n_262), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_117), .B(n_369), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_118), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_119), .A2(n_131), .B1(n_481), .B2(n_574), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_120), .A2(n_127), .B1(n_284), .B2(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_121), .A2(n_199), .B1(n_420), .B2(n_555), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_123), .Y(n_256) );
INVx1_ASAP7_75t_L g246 ( .A(n_124), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g281 ( .A1(n_125), .A2(n_172), .B1(n_282), .B2(n_284), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_126), .A2(n_150), .B1(n_520), .B2(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_130), .A2(n_144), .B1(n_291), .B2(n_454), .Y(n_572) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_132), .B(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_133), .A2(n_151), .B1(n_284), .B2(n_321), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_135), .A2(n_216), .B1(n_282), .B2(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g266 ( .A1(n_139), .A2(n_214), .B1(n_267), .B2(n_270), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_143), .A2(n_188), .B1(n_544), .B2(n_547), .Y(n_543) );
XNOR2x1_ASAP7_75t_L g327 ( .A(n_146), .B(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_147), .A2(n_167), .B1(n_419), .B2(n_420), .Y(n_418) );
AO22x1_ASAP7_75t_L g465 ( .A1(n_148), .A2(n_211), .B1(n_435), .B2(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_149), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_153), .A2(n_180), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_155), .A2(n_209), .B1(n_444), .B2(n_481), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_157), .A2(n_195), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_160), .A2(n_197), .B1(n_470), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_163), .A2(n_198), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_165), .A2(n_174), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_170), .A2(n_202), .B1(n_513), .B2(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_171), .B(n_395), .Y(n_394) );
XOR2x2_ASAP7_75t_L g530 ( .A(n_181), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_182), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g586 ( .A(n_182), .Y(n_586) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_184), .A2(n_594), .B1(n_595), .B2(n_617), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_184), .Y(n_617) );
OA22x2_ASAP7_75t_L g622 ( .A1(n_185), .A2(n_623), .B1(n_624), .B2(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_185), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_186), .A2(n_213), .B1(n_379), .B2(n_381), .Y(n_396) );
INVx1_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
AND2x2_ASAP7_75t_R g619 ( .A(n_189), .B(n_586), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_192), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_200), .B(n_228), .Y(n_227) );
XNOR2x1_ASAP7_75t_L g391 ( .A(n_201), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g302 ( .A(n_204), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_206), .A2(n_219), .B1(n_274), .B2(n_346), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_215), .Y(n_499) );
OA22x2_ASAP7_75t_L g356 ( .A1(n_218), .A2(n_357), .B1(n_358), .B2(n_385), .Y(n_356) );
INVx1_ASAP7_75t_L g385 ( .A(n_218), .Y(n_385) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_224), .B(n_227), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g646 ( .A(n_225), .B(n_227), .Y(n_646) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_226), .B(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_488), .B1(n_581), .B2(n_582), .C(n_583), .Y(n_230) );
INVx1_ASAP7_75t_L g581 ( .A(n_231), .Y(n_581) );
XNOR2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_388), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B1(n_323), .B2(n_324), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OA22x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_303), .B1(n_304), .B2(n_322), .Y(n_234) );
INVx1_ASAP7_75t_L g322 ( .A(n_235), .Y(n_322) );
XOR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_302), .Y(n_235) );
NAND2x1_ASAP7_75t_L g236 ( .A(n_237), .B(n_279), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_265), .Y(n_237) );
OAI21xp5_ASAP7_75t_SL g238 ( .A1(n_239), .A2(n_256), .B(n_257), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_249), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_241), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g346 ( .A(n_241), .B(n_278), .Y(n_346) );
AND2x2_ASAP7_75t_L g371 ( .A(n_241), .B(n_249), .Y(n_371) );
AND2x4_ASAP7_75t_L g377 ( .A(n_241), .B(n_271), .Y(n_377) );
AND2x4_ASAP7_75t_L g402 ( .A(n_241), .B(n_278), .Y(n_402) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
AND2x2_ASAP7_75t_L g260 ( .A(n_242), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_242), .Y(n_263) );
INVx2_ASAP7_75t_L g276 ( .A(n_242), .Y(n_276) );
OAI22x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B1(n_245), .B2(n_246), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g248 ( .A(n_244), .Y(n_248) );
INVx2_ASAP7_75t_L g252 ( .A(n_244), .Y(n_252) );
INVx1_ASAP7_75t_L g255 ( .A(n_244), .Y(n_255) );
INVx2_ASAP7_75t_L g261 ( .A(n_247), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_247), .B(n_276), .Y(n_275) );
BUFx2_ASAP7_75t_L g285 ( .A(n_247), .Y(n_285) );
AND2x4_ASAP7_75t_L g289 ( .A(n_249), .B(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g296 ( .A(n_249), .B(n_260), .Y(n_296) );
AND2x6_ASAP7_75t_L g300 ( .A(n_249), .B(n_275), .Y(n_300) );
AND2x2_ASAP7_75t_L g315 ( .A(n_249), .B(n_290), .Y(n_315) );
AND2x2_ASAP7_75t_L g317 ( .A(n_249), .B(n_260), .Y(n_317) );
AND2x2_ASAP7_75t_L g337 ( .A(n_249), .B(n_260), .Y(n_337) );
AND2x2_ASAP7_75t_L g415 ( .A(n_249), .B(n_275), .Y(n_415) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g259 ( .A(n_251), .B(n_253), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_254), .Y(n_264) );
INVx1_ASAP7_75t_L g269 ( .A(n_251), .Y(n_269) );
INVxp67_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g268 ( .A(n_254), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g274 ( .A(n_259), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g292 ( .A(n_259), .B(n_290), .Y(n_292) );
AND2x2_ASAP7_75t_L g310 ( .A(n_259), .B(n_275), .Y(n_310) );
AND2x2_ASAP7_75t_L g318 ( .A(n_259), .B(n_290), .Y(n_318) );
AND2x2_ASAP7_75t_L g380 ( .A(n_259), .B(n_260), .Y(n_380) );
AND2x4_ASAP7_75t_L g399 ( .A(n_259), .B(n_275), .Y(n_399) );
AND2x4_ASAP7_75t_L g267 ( .A(n_260), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g375 ( .A(n_260), .B(n_268), .Y(n_375) );
AND2x4_ASAP7_75t_L g290 ( .A(n_261), .B(n_276), .Y(n_290) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g383 ( .A(n_263), .B(n_264), .Y(n_383) );
AND2x4_ASAP7_75t_L g284 ( .A(n_264), .B(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g298 ( .A(n_264), .B(n_290), .Y(n_298) );
AND2x4_ASAP7_75t_L g314 ( .A(n_264), .B(n_290), .Y(n_314) );
AND2x4_ASAP7_75t_L g365 ( .A(n_264), .B(n_285), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_273), .Y(n_265) );
AND2x2_ASAP7_75t_L g283 ( .A(n_268), .B(n_275), .Y(n_283) );
AND2x6_ASAP7_75t_L g301 ( .A(n_268), .B(n_290), .Y(n_301) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_275), .Y(n_321) );
AND2x2_ASAP7_75t_SL g351 ( .A(n_268), .B(n_275), .Y(n_351) );
AND2x4_ASAP7_75t_L g422 ( .A(n_268), .B(n_290), .Y(n_422) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_269), .Y(n_272) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_293), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_286), .Y(n_280) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g445 ( .A(n_283), .Y(n_445) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_283), .Y(n_574) );
INVx3_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g419 ( .A(n_288), .Y(n_419) );
INVx2_ASAP7_75t_L g454 ( .A(n_288), .Y(n_454) );
INVx2_ASAP7_75t_SL g478 ( .A(n_288), .Y(n_478) );
INVx2_ASAP7_75t_SL g520 ( .A(n_288), .Y(n_520) );
INVx4_ASAP7_75t_L g555 ( .A(n_288), .Y(n_555) );
INVx8_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g557 ( .A(n_291), .Y(n_557) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g417 ( .A(n_292), .Y(n_417) );
BUFx3_ASAP7_75t_L g479 ( .A(n_292), .Y(n_479) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_292), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_299), .Y(n_293) );
BUFx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx3_ASAP7_75t_L g410 ( .A(n_296), .Y(n_410) );
INVx6_ASAP7_75t_L g484 ( .A(n_296), .Y(n_484) );
BUFx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
INVx2_ASAP7_75t_L g486 ( .A(n_298), .Y(n_486) );
BUFx2_ASAP7_75t_SL g514 ( .A(n_298), .Y(n_514) );
BUFx2_ASAP7_75t_SL g560 ( .A(n_298), .Y(n_560) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_306), .B(n_312), .Y(n_305) );
NAND4xp25_ASAP7_75t_SL g306 ( .A(n_307), .B(n_308), .C(n_309), .D(n_311), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .C(n_319), .D(n_320), .Y(n_312) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OA22x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_356), .B1(n_386), .B2(n_387), .Y(n_325) );
INVx1_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
XOR2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_340), .Y(n_326) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_334), .Y(n_328) );
NAND4xp25_ASAP7_75t_SL g329 ( .A(n_330), .B(n_331), .C(n_332), .D(n_333), .Y(n_329) );
NAND4xp25_ASAP7_75t_SL g334 ( .A(n_335), .B(n_336), .C(n_338), .D(n_339), .Y(n_334) );
NAND2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_348), .Y(n_341) );
NOR2x1_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_353), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NOR2xp67_ASAP7_75t_L g358 ( .A(n_359), .B(n_367), .Y(n_358) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .C(n_366), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx5_ASAP7_75t_SL g447 ( .A(n_365), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g367 ( .A(n_368), .B(n_372), .C(n_378), .D(n_384), .Y(n_367) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx4_ASAP7_75t_SL g395 ( .A(n_370), .Y(n_395) );
INVx3_ASAP7_75t_SL g431 ( .A(n_370), .Y(n_431) );
INVx4_ASAP7_75t_SL g472 ( .A(n_370), .Y(n_472) );
INVx3_ASAP7_75t_L g599 ( .A(n_370), .Y(n_599) );
INVx6_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g462 ( .A(n_374), .Y(n_462) );
INVx1_ASAP7_75t_L g502 ( .A(n_374), .Y(n_502) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_375), .Y(n_404) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_375), .Y(n_566) );
BUFx2_ASAP7_75t_SL g602 ( .A(n_376), .Y(n_602) );
BUFx6f_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g406 ( .A(n_377), .Y(n_406) );
BUFx3_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
INVx2_ASAP7_75t_L g464 ( .A(n_377), .Y(n_464) );
BUFx4f_ASAP7_75t_L g632 ( .A(n_377), .Y(n_632) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_379), .Y(n_604) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx3_ASAP7_75t_L g434 ( .A(n_380), .Y(n_434) );
INVx2_ASAP7_75t_L g467 ( .A(n_380), .Y(n_467) );
BUFx5_ASAP7_75t_L g630 ( .A(n_380), .Y(n_630) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_381), .Y(n_539) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g606 ( .A(n_382), .Y(n_606) );
INVx2_ASAP7_75t_L g629 ( .A(n_382), .Y(n_629) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx12f_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_423), .B1(n_424), .B2(n_487), .Y(n_388) );
INVx2_ASAP7_75t_L g487 ( .A(n_389), .Y(n_487) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_407), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .C(n_397), .D(n_403), .Y(n_393) );
BUFx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_399), .Y(n_470) );
BUFx3_ASAP7_75t_L g568 ( .A(n_399), .Y(n_568) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_401), .A2(n_506), .B1(n_507), .B2(n_509), .Y(n_505) );
INVx2_ASAP7_75t_SL g608 ( .A(n_401), .Y(n_608) );
INVx6_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .C(n_412), .D(n_418), .Y(n_407) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
INVx2_ASAP7_75t_SL g523 ( .A(n_414), .Y(n_523) );
INVx2_ASAP7_75t_L g615 ( .A(n_414), .Y(n_615) );
INVx2_ASAP7_75t_SL g637 ( .A(n_414), .Y(n_637) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g449 ( .A(n_415), .Y(n_449) );
BUFx2_ASAP7_75t_L g546 ( .A(n_415), .Y(n_546) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g450 ( .A(n_421), .Y(n_450) );
INVx2_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
INVx1_ASAP7_75t_SL g521 ( .A(n_421), .Y(n_521) );
INVx2_ASAP7_75t_L g547 ( .A(n_421), .Y(n_547) );
INVx2_ASAP7_75t_SL g635 ( .A(n_421), .Y(n_635) );
INVx8_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_426), .B1(n_456), .B2(n_457), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
XNOR2x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_455), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_441), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_436), .Y(n_428) );
OAI21xp33_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B(n_433), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_430), .A2(n_494), .B1(n_495), .B2(n_496), .C(n_497), .Y(n_493) );
INVx2_ASAP7_75t_L g541 ( .A(n_430), .Y(n_541) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g496 ( .A(n_434), .Y(n_496) );
BUFx6f_ASAP7_75t_SL g538 ( .A(n_434), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
BUFx6f_ASAP7_75t_SL g534 ( .A(n_440), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_451), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g517 ( .A(n_445), .Y(n_517) );
INVx1_ASAP7_75t_L g550 ( .A(n_445), .Y(n_550) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
INVx2_ASAP7_75t_L g551 ( .A(n_447), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_473), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .C(n_468), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_471), .Y(n_468) );
BUFx4f_ASAP7_75t_SL g508 ( .A(n_470), .Y(n_508) );
BUFx2_ASAP7_75t_L g536 ( .A(n_470), .Y(n_536) );
AND4x1_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .C(n_480), .D(n_482), .Y(n_473) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g513 ( .A(n_484), .Y(n_513) );
INVx1_ASAP7_75t_SL g559 ( .A(n_484), .Y(n_559) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g640 ( .A(n_486), .Y(n_640) );
INVx1_ASAP7_75t_L g582 ( .A(n_488), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_527), .B1(n_528), .B2(n_580), .Y(n_488) );
INVx1_ASAP7_75t_L g580 ( .A(n_489), .Y(n_580) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_510), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_505), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_503), .B2(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_515), .Y(n_511) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_526), .Y(n_616) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_530), .B1(n_561), .B2(n_579), .Y(n_528) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_532), .B(n_542), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .C(n_537), .D(n_540), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .C(n_552), .D(n_558), .Y(n_542) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g579 ( .A(n_561), .Y(n_579) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g578 ( .A(n_563), .Y(n_578) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_571), .Y(n_563) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .C(n_569), .D(n_570), .Y(n_564) );
BUFx6f_ASAP7_75t_SL g601 ( .A(n_566), .Y(n_601) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .C(n_575), .D(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_585), .B(n_588), .Y(n_643) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_618), .B1(n_620), .B2(n_623), .C1(n_641), .C2(n_644), .Y(n_592) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_609), .Y(n_595) );
NAND4xp25_ASAP7_75t_SL g596 ( .A(n_597), .B(n_600), .C(n_603), .D(n_607), .Y(n_596) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .C(n_612), .D(n_613), .Y(n_609) );
BUFx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_633), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .C(n_631), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .C(n_638), .D(n_639), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_642), .Y(n_641) );
CKINVDCx6p67_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_645), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_646), .Y(n_645) );
endmodule