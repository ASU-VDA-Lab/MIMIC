module fake_jpeg_9518_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_47),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_55),
.B1(n_58),
.B2(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_25),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_22),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_72),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_25),
.B1(n_22),
.B2(n_28),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_19),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_26),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_89)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_30),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_14),
.B(n_10),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_75),
.A2(n_59),
.B(n_74),
.C(n_73),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_35),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_80),
.Y(n_133)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_82),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_81),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_97),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_95),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_46),
.B1(n_27),
.B2(n_23),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_98),
.B1(n_29),
.B2(n_17),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_35),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_24),
.B(n_29),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_54),
.B(n_28),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_46),
.B1(n_26),
.B2(n_34),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_24),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_108),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_35),
.B1(n_15),
.B2(n_8),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_56),
.A2(n_35),
.B1(n_14),
.B2(n_13),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_56),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_48),
.Y(n_116)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_138),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_0),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_122),
.B(n_24),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_57),
.B(n_61),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_62),
.B1(n_57),
.B2(n_65),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_125),
.B1(n_127),
.B2(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_62),
.B1(n_65),
.B2(n_26),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_136),
.B(n_142),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_90),
.B1(n_101),
.B2(n_98),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_26),
.B1(n_29),
.B2(n_17),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_75),
.B(n_111),
.C(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_69),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_29),
.B(n_34),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_102),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_168),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_145),
.B(n_154),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_107),
.B1(n_80),
.B2(n_94),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_178)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_139),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_87),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_159),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_107),
.B1(n_75),
.B2(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_92),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_93),
.B1(n_87),
.B2(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_166),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_0),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_167),
.B(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_36),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_164),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_36),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_165),
.B(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_134),
.B(n_7),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_34),
.B(n_29),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_76),
.B(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_38),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_78),
.B1(n_92),
.B2(n_39),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_175),
.B1(n_129),
.B2(n_139),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_39),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_121),
.A2(n_78),
.B1(n_39),
.B2(n_40),
.Y(n_175)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_12),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_185),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_141),
.B1(n_126),
.B2(n_125),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_182),
.A2(n_147),
.B1(n_150),
.B2(n_172),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_117),
.B(n_124),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_210),
.B(n_177),
.Y(n_222)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_117),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_198),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_135),
.B(n_117),
.C(n_84),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_153),
.B1(n_162),
.B2(n_167),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_38),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_206),
.C(n_59),
.Y(n_234)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_176),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_208),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_18),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

AO32x1_ASAP7_75t_L g210 ( 
.A1(n_150),
.A2(n_59),
.A3(n_29),
.B1(n_73),
.B2(n_74),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_157),
.B(n_168),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_216),
.B1(n_226),
.B2(n_233),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_218),
.B(n_225),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_171),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_238),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_156),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_228),
.C(n_234),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_157),
.CI(n_160),
.CON(n_225),
.SN(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_147),
.B1(n_167),
.B2(n_152),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_230),
.B1(n_235),
.B2(n_204),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_160),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_178),
.A2(n_161),
.B1(n_172),
.B2(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_114),
.B1(n_86),
.B2(n_83),
.Y(n_233)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_59),
.B1(n_105),
.B2(n_114),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_38),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_178),
.C(n_182),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_199),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_189),
.B(n_29),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_180),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_241),
.B(n_249),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_246),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_205),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_247),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_221),
.B(n_180),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_252),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_237),
.B(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_220),
.B(n_203),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_258),
.C(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_213),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_226),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_219),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_191),
.C(n_201),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_266),
.C(n_272),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_260),
.B1(n_246),
.B2(n_259),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_243),
.B(n_236),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_216),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_201),
.C(n_227),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_222),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_230),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_225),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_202),
.C(n_181),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_257),
.B1(n_240),
.B2(n_254),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_294),
.B1(n_270),
.B2(n_277),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_200),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_276),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_295),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_247),
.B(n_257),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_211),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_279),
.Y(n_297)
);

AOI21x1_ASAP7_75t_SL g291 ( 
.A1(n_263),
.A2(n_240),
.B(n_225),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_292),
.B(n_268),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_245),
.B(n_239),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_294),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_262),
.A2(n_192),
.B1(n_209),
.B2(n_203),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_265),
.C(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_299),
.Y(n_310)
);

AO221x1_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_288),
.B1(n_289),
.B2(n_284),
.C(n_192),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_300),
.A2(n_293),
.B1(n_286),
.B2(n_283),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_307),
.B1(n_1),
.B2(n_2),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_200),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_309),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_287),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_286),
.B1(n_283),
.B2(n_281),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_266),
.B1(n_185),
.B2(n_3),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_312),
.A2(n_314),
.B(n_308),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_313),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_281),
.B(n_7),
.C(n_11),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_24),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_302),
.B(n_1),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_309),
.Y(n_320)
);

AOI31xp67_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_321),
.A3(n_2),
.B(n_4),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_298),
.Y(n_321)
);

OAI221xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_315),
.B1(n_311),
.B2(n_312),
.C(n_313),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_301),
.C(n_307),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_18),
.C(n_3),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_329),
.B(n_325),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

OAI311xp33_ASAP7_75t_L g333 ( 
.A1(n_331),
.A2(n_326),
.A3(n_322),
.B1(n_5),
.C1(n_4),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_4),
.C(n_5),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_4),
.Y(n_336)
);


endmodule