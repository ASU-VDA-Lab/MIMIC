module real_jpeg_29510_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_1),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_1),
.A2(n_59),
.B1(n_60),
.B2(n_100),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_100),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_1),
.A2(n_25),
.B1(n_30),
.B2(n_100),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_2),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_79),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_25),
.B1(n_30),
.B2(n_79),
.Y(n_193)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_69),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_69),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_7),
.A2(n_25),
.B1(n_30),
.B2(n_69),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_25),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_8),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_25),
.B1(n_30),
.B2(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_10),
.A2(n_58),
.B(n_59),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_10),
.B(n_39),
.Y(n_204)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_10),
.A2(n_39),
.B(n_43),
.C(n_204),
.D(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_73),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_24),
.B(n_217),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g245 ( 
.A1(n_10),
.A2(n_60),
.B(n_72),
.C(n_156),
.D(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_10),
.B(n_60),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_39),
.B(n_44),
.C(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_12),
.A2(n_41),
.B1(n_59),
.B2(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_41),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_15),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_15),
.A2(n_25),
.B1(n_30),
.B2(n_66),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_249)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_20),
.B(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_91),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_21),
.B(n_83),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_51),
.B1(n_52),
.B2(n_82),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_23),
.B(n_37),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_24),
.A2(n_35),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_24),
.A2(n_29),
.B1(n_34),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_24),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_24),
.A2(n_34),
.B1(n_150),
.B2(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_24),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_24),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_25),
.A2(n_30),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_25),
.B(n_45),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_30),
.A2(n_40),
.A3(n_46),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_30),
.B(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_33),
.A2(n_95),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_33),
.B(n_218),
.Y(n_217)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_34),
.B(n_144),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_45),
.Y(n_44)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_39),
.A2(n_59),
.A3(n_246),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_40),
.B(n_77),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_42),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_47),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_43),
.A2(n_47),
.B1(n_87),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_43),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_43),
.A2(n_47),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_50),
.A2(n_97),
.B(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_50),
.B(n_172),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_50),
.A2(n_170),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_50),
.B(n_144),
.Y(n_230)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_70),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_70),
.C(n_82),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_64),
.B(n_67),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_55),
.B(n_68),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_55),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_62),
.B(n_144),
.C(n_145),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_67),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_71),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_73),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_72),
.A2(n_73),
.B1(n_154),
.B2(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_77),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_80),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_105),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_80),
.A2(n_103),
.B(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_89),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_89),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_90),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_90),
.A2(n_224),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.C(n_101),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_134),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_126),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_116),
.B1(n_117),
.B2(n_125),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_115),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_112),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_123),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_121),
.B(n_144),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_159),
.B(n_275),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_157),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_131),
.B(n_157),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.C(n_136),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_132),
.B(n_135),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_137),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_151),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_139),
.B1(n_151),
.B2(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_148),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_196),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_182),
.B(n_195),
.Y(n_161)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_162),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_179),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_179),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_185),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_190),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_189),
.B(n_190),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_191),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_192),
.B(n_194),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_273),
.C(n_274),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_268),
.B(n_272),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_257),
.B(n_267),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_241),
.B(n_256),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_220),
.B(n_240),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_208),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_202),
.B(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_206),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_214),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_216),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_228),
.B(n_239),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_227),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_226),
.A2(n_233),
.B(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_234),
.B(n_238),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_247),
.C(n_250),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_253),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.C(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);


endmodule