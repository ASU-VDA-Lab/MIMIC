module real_jpeg_23493_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_25),
.B1(n_32),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_3),
.Y(n_97)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_37),
.C(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_30),
.B1(n_72),
.B2(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_89),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_121),
.B1(n_160),
.B2(n_164),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_8),
.A2(n_25),
.B1(n_32),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_8),
.A2(n_65),
.B1(n_82),
.B2(n_83),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_8),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_65),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_32),
.C(n_33),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_25),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_12),
.A2(n_72),
.B1(n_73),
.B2(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_91),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_13),
.A2(n_72),
.B1(n_73),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_100),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_15),
.Y(n_164)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_15),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_103),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_103),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_51),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B(n_27),
.C(n_31),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_23),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_23),
.A2(n_33),
.B1(n_82),
.B2(n_84),
.Y(n_81)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_25),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_25),
.B(n_30),
.CON(n_118),
.SN(n_118)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_27),
.A2(n_60),
.B1(n_80),
.B2(n_85),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_30),
.CON(n_27),
.SN(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_30),
.B(n_98),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_30),
.B(n_167),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g119 ( 
.A(n_32),
.B(n_69),
.C(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_43),
.B2(n_47),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_35),
.A2(n_54),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_36),
.A2(n_37),
.B1(n_96),
.B2(n_97),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_36),
.B(n_166),
.Y(n_165)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_38),
.B(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_38),
.Y(n_161)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_53),
.B(n_55),
.Y(n_52)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_46),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.C(n_62),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_71),
.B2(n_75),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_64),
.A2(n_67),
.B1(n_89),
.B2(n_118),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_76),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_72),
.B(n_117),
.C(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_73),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_87),
.Y(n_78)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_99),
.B(n_101),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_112),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_93),
.A2(n_110),
.B1(n_112),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_98),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_113),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_104),
.A2(n_105),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_108),
.A2(n_113),
.B1(n_114),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_153),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_181),
.B(n_187),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_171),
.B(n_180),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_149),
.B(n_170),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_133),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_144),
.C(n_147),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_156),
.B(n_169),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_155),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_162),
.B(n_168),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_179),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);


endmodule