module fake_jpeg_16081_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_25),
.Y(n_66)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_26),
.B1(n_39),
.B2(n_47),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_59),
.B(n_32),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_37),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_26),
.B1(n_17),
.B2(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_17),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_33),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_69),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_72),
.B1(n_31),
.B2(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_33),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_33),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_32),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_19),
.B1(n_23),
.B2(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_92),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_47),
.B1(n_45),
.B2(n_19),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_99),
.B1(n_93),
.B2(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_99),
.B(n_88),
.C(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_87),
.A2(n_89),
.B(n_32),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_28),
.B1(n_24),
.B2(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_96),
.Y(n_124)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_49),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_23),
.C(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_59),
.A2(n_21),
.B1(n_70),
.B2(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_36),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_70),
.B1(n_49),
.B2(n_50),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_61),
.B1(n_70),
.B2(n_50),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_56),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_84),
.CI(n_90),
.CON(n_105),
.SN(n_105)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_76),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_111),
.B1(n_131),
.B2(n_74),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_119),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_103),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_101),
.B(n_76),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_61),
.B1(n_54),
.B2(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_127),
.B1(n_128),
.B2(n_32),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_54),
.B1(n_67),
.B2(n_56),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_67),
.B1(n_56),
.B2(n_21),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_116),
.B(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_21),
.B1(n_36),
.B2(n_18),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_38),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_96),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_96),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_141),
.B(n_147),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_73),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_158),
.B1(n_162),
.B2(n_130),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_91),
.C(n_85),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_140),
.C(n_143),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_85),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_85),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_152),
.B(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_132),
.A3(n_104),
.B1(n_124),
.B2(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_149),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_80),
.C(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_151),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_80),
.B(n_94),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_125),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_161),
.B1(n_118),
.B2(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_95),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_75),
.B1(n_52),
.B2(n_12),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_27),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_117),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_106),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_27),
.C(n_75),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_165),
.B(n_166),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_113),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_167),
.A2(n_178),
.B(n_30),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_168),
.A2(n_179),
.B1(n_193),
.B2(n_154),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_160),
.B1(n_134),
.B2(n_162),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_170),
.B(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_112),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_194),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_157),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_120),
.B1(n_106),
.B2(n_104),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_191),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_106),
.B1(n_120),
.B2(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_183),
.A2(n_38),
.B1(n_48),
.B2(n_42),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_115),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_129),
.C(n_127),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_42),
.C(n_75),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_139),
.B(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_111),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_125),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_159),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_137),
.A2(n_118),
.B1(n_107),
.B2(n_108),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_108),
.B(n_107),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_32),
.B(n_38),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_138),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_219),
.C(n_220),
.Y(n_242)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_202),
.B(n_203),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_142),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_206),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_171),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_141),
.B(n_161),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_225),
.B(n_167),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_178),
.A2(n_152),
.B1(n_142),
.B2(n_154),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_216),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_221),
.B(n_185),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_52),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_222),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_30),
.C(n_18),
.Y(n_220)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_182),
.B1(n_172),
.B2(n_191),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_166),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_195),
.A2(n_0),
.B(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_222),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_230),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_197),
.B(n_174),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_227),
.B(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_252),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_235),
.B1(n_239),
.B2(n_218),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_234),
.B(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_183),
.B1(n_172),
.B2(n_190),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_197),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_240),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_188),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_238),
.A2(n_245),
.B(n_211),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_180),
.B(n_167),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_187),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_186),
.C(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_248),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_209),
.B(n_208),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_180),
.C(n_170),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_190),
.C(n_179),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_251),
.A2(n_201),
.B(n_173),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_257),
.A2(n_231),
.B(n_241),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_204),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_265),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_210),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_263),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_214),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_218),
.B1(n_225),
.B2(n_215),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_267),
.B1(n_8),
.B2(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_223),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_165),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_273),
.C(n_236),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_227),
.B(n_202),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_198),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_274),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_18),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_9),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_280),
.C(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_233),
.B1(n_250),
.B2(n_229),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_279),
.A2(n_285),
.B1(n_263),
.B2(n_271),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_248),
.C(n_229),
.Y(n_280)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_239),
.C(n_234),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_226),
.C(n_231),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_287),
.C(n_254),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_259),
.B(n_262),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_9),
.Y(n_287)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_296),
.C(n_8),
.Y(n_317)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_298),
.B(n_302),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_304),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.Y(n_312)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_258),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_10),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_299),
.A2(n_276),
.B(n_283),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_0),
.B(n_3),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_296),
.A2(n_284),
.B1(n_280),
.B2(n_278),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_318),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_292),
.B1(n_287),
.B2(n_261),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_295),
.B1(n_297),
.B2(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_11),
.C(n_13),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_10),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_330),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_294),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_328),
.C(n_311),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_294),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_325),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_308),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_326),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_3),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_3),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_327),
.B(n_314),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_337),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_312),
.Y(n_337)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_313),
.Y(n_339)
);

OAI221xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_340),
.B1(n_335),
.B2(n_312),
.C(n_333),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_342),
.A2(n_343),
.B(n_330),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_321),
.C(n_310),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_341),
.B(n_4),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_4),
.C(n_5),
.Y(n_346)
);

A2O1A1O1Ixp25_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_4),
.B(n_5),
.C(n_339),
.D(n_267),
.Y(n_347)
);


endmodule