module fake_netlist_6_2553_n_2108 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2108);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2108;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_83),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_202),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_98),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_87),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_93),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_33),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_89),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_112),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_44),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_54),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_107),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_39),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_24),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_161),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_126),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_146),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_22),
.Y(n_254)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_81),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_14),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_188),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_180),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_154),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_153),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_88),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_68),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_101),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_64),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_54),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_116),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_44),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_158),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_170),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_67),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_97),
.Y(n_275)
);

BUFx2_ASAP7_75t_SL g276 ( 
.A(n_41),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_71),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_91),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_63),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_69),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_120),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_34),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_90),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_122),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_102),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_139),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_123),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_7),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_189),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_84),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_219),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_64),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_53),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_216),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_32),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_152),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_160),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_94),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_168),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_218),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_130),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_132),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_156),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_27),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_131),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_179),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_111),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_195),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_76),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_194),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_12),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_99),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_215),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_57),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_49),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_18),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_187),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_63),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_7),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_148),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_196),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_61),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_59),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_78),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_171),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_39),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_53),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_14),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_16),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_29),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_8),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_41),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_117),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_35),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_197),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_136),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_151),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_47),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_19),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_157),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_37),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_164),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_19),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_100),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_214),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_45),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_169),
.Y(n_357)
);

BUFx8_ASAP7_75t_SL g358 ( 
.A(n_105),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_142),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_185),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_147),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_166),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_67),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_176),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_81),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_21),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_143),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_52),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_26),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_46),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_60),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_42),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_192),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_106),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_11),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_50),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_118),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_109),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_208),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_49),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_210),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_13),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_95),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_52),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_65),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_162),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_184),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_31),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_135),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_198),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_68),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_121),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_199),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_206),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_174),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_61),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_203),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_129),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_0),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_115),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_11),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_200),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_0),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_40),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_85),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_59),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_76),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_138),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_25),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_172),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_74),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_134),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_36),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_1),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_15),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_159),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_43),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_74),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_177),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_137),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_62),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_28),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_48),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_173),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_50),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_4),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_149),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_178),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_71),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_321),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_261),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_265),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_358),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_338),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_346),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_345),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_349),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_372),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_224),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_228),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_229),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_355),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_233),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_230),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_233),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_335),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_258),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_238),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_335),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_241),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_351),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_247),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_250),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_252),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_351),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_223),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_223),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_338),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_253),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_231),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_260),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_258),
.B(n_2),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_277),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_277),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_262),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_276),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_273),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_303),
.B(n_431),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_282),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_277),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_225),
.B(n_3),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_287),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_385),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_385),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_288),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_225),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_292),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_276),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_293),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_297),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_226),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_301),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_226),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_305),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_306),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_308),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_309),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_310),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_311),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_239),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_239),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_395),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_240),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_323),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_324),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_330),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_291),
.B(n_3),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_303),
.B(n_4),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_240),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_245),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_331),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_343),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_245),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_344),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_350),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_320),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_431),
.B(n_5),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_352),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_246),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_354),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_246),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_266),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_284),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_317),
.B(n_5),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_266),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_362),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_361),
.B(n_9),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_395),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_365),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_376),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_380),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_381),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_274),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_274),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_382),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_280),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_243),
.Y(n_544)
);

INVxp67_ASAP7_75t_SL g545 ( 
.A(n_284),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_280),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_384),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_440),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_470),
.B(n_361),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_479),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_515),
.B(n_304),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_479),
.B(n_361),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_441),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_442),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_283),
.B1(n_312),
.B2(n_254),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_434),
.A2(n_422),
.B1(n_427),
.B2(n_319),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_442),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_480),
.B(n_231),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_453),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_544),
.B(n_286),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_478),
.B(n_279),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_480),
.B(n_232),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_493),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_498),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_498),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_455),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_438),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_545),
.B(n_432),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_500),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_455),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_457),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_451),
.B(n_221),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_507),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_469),
.A2(n_267),
.B1(n_332),
.B2(n_347),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_386),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_435),
.B(n_436),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_508),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_457),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_486),
.B(n_232),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_458),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_461),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_454),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_464),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_489),
.B(n_391),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g605 ( 
.A(n_437),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_510),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_462),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_489),
.B(n_396),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_509),
.B(n_285),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_468),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_475),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_490),
.B(n_491),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_475),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_490),
.B(n_397),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_477),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_516),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_459),
.B(n_257),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_491),
.B(n_236),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_477),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_516),
.B(n_398),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_520),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_534),
.A2(n_237),
.B(n_236),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_528),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_448),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_443),
.A2(n_255),
.B1(n_342),
.B2(n_341),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_528),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_529),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_529),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_532),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_532),
.B(n_220),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_540),
.A2(n_244),
.B(n_237),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_482),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_535),
.B(n_285),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_582),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_557),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_557),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_570),
.B(n_279),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_620),
.A2(n_587),
.B1(n_465),
.B2(n_483),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_629),
.A2(n_524),
.B1(n_445),
.B2(n_487),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_553),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_570),
.A2(n_531),
.B1(n_307),
.B2(n_329),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g647 ( 
.A(n_628),
.B(n_481),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_577),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_576),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_577),
.B(n_449),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_583),
.B(n_450),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_629),
.A2(n_517),
.B1(n_514),
.B2(n_222),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_580),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_L g655 ( 
.A(n_591),
.B(n_495),
.C(n_526),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_557),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_577),
.B(n_456),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_580),
.Y(n_660)
);

AND3x2_ASAP7_75t_L g661 ( 
.A(n_582),
.B(n_234),
.C(n_220),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_614),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_576),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_561),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_561),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_565),
.B(n_279),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_561),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_626),
.B(n_234),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_553),
.Y(n_670)
);

BUFx6f_ASAP7_75t_SL g671 ( 
.A(n_628),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_570),
.B(n_279),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_570),
.A2(n_307),
.B1(n_329),
.B2(n_296),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_580),
.A2(n_496),
.B1(n_499),
.B2(n_494),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_614),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_554),
.A2(n_264),
.B1(n_269),
.B2(n_244),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_593),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_580),
.A2(n_502),
.B1(n_504),
.B2(n_501),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_577),
.B(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_577),
.B(n_463),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_551),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_580),
.A2(n_554),
.B1(n_636),
.B2(n_609),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_565),
.B(n_540),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_576),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_577),
.B(n_466),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_576),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_583),
.B(n_259),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_551),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_576),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_570),
.A2(n_333),
.B1(n_334),
.B2(n_296),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_576),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_SL g693 ( 
.A(n_628),
.B(n_505),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_565),
.B(n_279),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_628),
.B(n_467),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_551),
.B(n_264),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_548),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_570),
.B(n_279),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_563),
.Y(n_699)
);

NOR2x1p5_ASAP7_75t_L g700 ( 
.A(n_609),
.B(n_227),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_637),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_636),
.B(n_473),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_579),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_476),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_563),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_637),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_554),
.B(n_304),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_549),
.Y(n_709)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_593),
.Y(n_710)
);

HB1xp67_ASAP7_75t_SL g711 ( 
.A(n_575),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_579),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_566),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_579),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_548),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_570),
.A2(n_334),
.B1(n_337),
.B2(n_333),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_575),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_607),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_548),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_553),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_592),
.B(n_485),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_579),
.Y(n_723)
);

INVxp33_ASAP7_75t_L g724 ( 
.A(n_607),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_604),
.B(n_488),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_631),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_554),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_572),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_572),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_570),
.B(n_604),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_573),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_549),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_608),
.B(n_259),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_566),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_566),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_548),
.Y(n_737)
);

AND2x4_ASAP7_75t_L g738 ( 
.A(n_549),
.B(n_269),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_570),
.A2(n_371),
.B1(n_400),
.B2(n_337),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_608),
.B(n_492),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_562),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_623),
.B(n_503),
.C(n_497),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_631),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_616),
.B(n_268),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_574),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_616),
.B(n_506),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_602),
.B(n_512),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_623),
.B(n_302),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_562),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_574),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_631),
.B(n_268),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_578),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_552),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_571),
.B(n_513),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_554),
.A2(n_373),
.B1(n_400),
.B2(n_403),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_554),
.A2(n_519),
.B1(n_511),
.B2(n_527),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_602),
.B(n_518),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_578),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_555),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_571),
.B(n_521),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_552),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_584),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_584),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_568),
.B(n_522),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_571),
.B(n_525),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_631),
.B(n_272),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_555),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_605),
.B(n_537),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_635),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_596),
.B(n_533),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_634),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_626),
.A2(n_373),
.B1(n_353),
.B2(n_408),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_564),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_555),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_559),
.A2(n_539),
.B1(n_538),
.B2(n_536),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_559),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_552),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_552),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_588),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_596),
.B(n_542),
.Y(n_781)
);

NOR2x1p5_ASAP7_75t_L g782 ( 
.A(n_588),
.B(n_235),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_548),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_631),
.B(n_272),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_564),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_548),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_550),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_635),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_560),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_589),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_591),
.A2(n_547),
.B1(n_452),
.B2(n_444),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_596),
.B(n_439),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_711),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_669),
.A2(n_626),
.B1(n_635),
.B2(n_621),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_662),
.B(n_302),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_775),
.B(n_316),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_709),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_662),
.B(n_302),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_652),
.B(n_626),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_709),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_755),
.B(n_357),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_742),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_727),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_761),
.B(n_360),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_662),
.B(n_302),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_L g806 ( 
.A(n_702),
.B(n_560),
.C(n_621),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_742),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_727),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_750),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_782),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_768),
.B(n_302),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_766),
.B(n_242),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_718),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_771),
.B(n_248),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_774),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_768),
.B(n_302),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_705),
.B(n_621),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_731),
.B(n_320),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_722),
.B(n_631),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_643),
.B(n_251),
.C(n_249),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_718),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_687),
.A2(n_594),
.B(n_606),
.C(n_633),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_682),
.A2(n_409),
.B1(n_423),
.B2(n_399),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_728),
.A2(n_300),
.B1(n_275),
.B2(n_377),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_725),
.B(n_635),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_781),
.B(n_404),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_645),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_L g828 ( 
.A1(n_708),
.A2(n_327),
.B1(n_313),
.B2(n_299),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_774),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_741),
.B(n_635),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_656),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_669),
.B(n_320),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_785),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_776),
.B(n_263),
.C(n_256),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_747),
.B(n_270),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_770),
.A2(n_300),
.B(n_289),
.C(n_294),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_644),
.B(n_567),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_646),
.A2(n_634),
.B1(n_299),
.B2(n_340),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_728),
.A2(n_406),
.B1(n_414),
.B2(n_416),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_785),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_655),
.B(n_792),
.C(n_765),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_760),
.A2(n_420),
.B1(n_428),
.B2(n_634),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_654),
.B(n_320),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_756),
.B(n_278),
.C(n_271),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_770),
.A2(n_634),
.B1(n_313),
.B2(n_289),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_644),
.B(n_567),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_760),
.B(n_286),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_695),
.B(n_286),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_654),
.A2(n_275),
.B1(n_294),
.B2(n_315),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_653),
.B(n_290),
.C(n_281),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_733),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_748),
.B(n_295),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_663),
.A2(n_315),
.B1(n_327),
.B2(n_340),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_SL g854 ( 
.A1(n_647),
.A2(n_286),
.B1(n_243),
.B2(n_410),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_644),
.B(n_569),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_657),
.B(n_569),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_675),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_657),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_639),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_724),
.B(n_589),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_674),
.B(n_678),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_660),
.A2(n_359),
.B1(n_368),
.B2(n_377),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_681),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_733),
.B(n_590),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_657),
.B(n_598),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_772),
.B(n_320),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_688),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_660),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_670),
.B(n_598),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_708),
.A2(n_389),
.B1(n_424),
.B2(n_412),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_670),
.B(n_598),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_772),
.B(n_320),
.Y(n_873)
);

BUFx8_ASAP7_75t_L g874 ( 
.A(n_671),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_772),
.B(n_320),
.Y(n_875)
);

OAI221xp5_ASAP7_75t_L g876 ( 
.A1(n_773),
.A2(n_353),
.B1(n_366),
.B2(n_371),
.C(n_375),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_670),
.B(n_598),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_729),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_721),
.B(n_600),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_642),
.B(n_590),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_640),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_719),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_721),
.B(n_683),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_730),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_640),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_732),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_719),
.B(n_366),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_739),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_701),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_721),
.B(n_600),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_748),
.B(n_298),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_683),
.B(n_600),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_788),
.B(n_320),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_746),
.B(n_600),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_658),
.Y(n_895)
);

NOR2xp67_ASAP7_75t_L g896 ( 
.A(n_743),
.B(n_594),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_751),
.B(n_611),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_753),
.B(n_611),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_724),
.B(n_707),
.Y(n_899)
);

NAND2x1_ASAP7_75t_L g900 ( 
.A(n_648),
.B(n_754),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_658),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_665),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_759),
.B(n_611),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_788),
.B(n_320),
.Y(n_904)
);

NOR2x1p5_ASAP7_75t_L g905 ( 
.A(n_758),
.B(n_314),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_763),
.B(n_611),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_665),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_666),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_666),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_708),
.A2(n_359),
.B1(n_368),
.B2(n_389),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_780),
.B(n_612),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_790),
.B(n_612),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_687),
.A2(n_412),
.B1(n_402),
.B2(n_424),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_758),
.B(n_318),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_738),
.B(n_612),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_668),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_754),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_651),
.B(n_393),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_738),
.B(n_612),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_668),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_691),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_754),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_738),
.B(n_622),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_762),
.B(n_622),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_693),
.B(n_597),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_671),
.A2(n_393),
.B1(n_394),
.B2(n_401),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_691),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_707),
.B(n_322),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_676),
.B(n_597),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_R g931 ( 
.A(n_638),
.B(n_325),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_762),
.B(n_394),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_671),
.A2(n_696),
.B1(n_700),
.B2(n_734),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_762),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_699),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_778),
.B(n_622),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_778),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_696),
.B(n_606),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_696),
.B(n_617),
.Y(n_939)
);

AO221x1_ASAP7_75t_L g940 ( 
.A1(n_778),
.A2(n_403),
.B1(n_429),
.B2(n_375),
.C(n_415),
.Y(n_940)
);

INVx8_ASAP7_75t_L g941 ( 
.A(n_638),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_699),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_779),
.B(n_734),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_706),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_L g945 ( 
.A(n_757),
.B(n_617),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_779),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_777),
.B(n_326),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_779),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_706),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_713),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_659),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_745),
.B(n_622),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_791),
.B(n_619),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_713),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_679),
.B(n_619),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_735),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_745),
.B(n_581),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_735),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_680),
.B(n_581),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_789),
.B(n_328),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_769),
.B(n_624),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_882),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_859),
.A2(n_883),
.B(n_819),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_859),
.A2(n_685),
.B(n_783),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_817),
.B(n_673),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_802),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_801),
.B(n_804),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_959),
.A2(n_672),
.B(n_641),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_865),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_690),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_797),
.B(n_667),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_865),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_865),
.Y(n_974)
);

AND3x1_ASAP7_75t_SL g975 ( 
.A(n_905),
.B(n_415),
.C(n_408),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_821),
.B(n_710),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_807),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_899),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_841),
.B(n_661),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_837),
.A2(n_672),
.B(n_641),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_846),
.A2(n_698),
.B(n_649),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_797),
.B(n_667),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_855),
.A2(n_698),
.B(n_649),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_799),
.A2(n_740),
.B(n_717),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_796),
.B(n_703),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_804),
.B(n_786),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_835),
.B(n_786),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_832),
.A2(n_749),
.B(n_712),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_857),
.A2(n_649),
.B(n_716),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_861),
.B(n_624),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_866),
.A2(n_720),
.B(n_716),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_832),
.A2(n_749),
.B(n_784),
.C(n_767),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_795),
.A2(n_715),
.B(n_704),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_835),
.B(n_726),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_796),
.B(n_812),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_852),
.B(n_632),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_806),
.B(n_723),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_812),
.B(n_786),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_814),
.B(n_787),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_814),
.B(n_787),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_797),
.B(n_726),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_852),
.A2(n_401),
.B(n_402),
.C(n_767),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_827),
.B(n_787),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_870),
.A2(n_720),
.B(n_716),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_831),
.B(n_858),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_L g1006 ( 
.A(n_941),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_938),
.B(n_667),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_L g1008 ( 
.A1(n_795),
.A2(n_784),
.B(n_752),
.C(n_736),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_893),
.A2(n_752),
.B(n_632),
.C(n_633),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_807),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_891),
.A2(n_736),
.B(n_429),
.C(n_425),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_825),
.A2(n_694),
.B(n_667),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_938),
.B(n_667),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_L g1014 ( 
.A1(n_798),
.A2(n_737),
.B(n_720),
.C(n_630),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_938),
.B(n_667),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_L g1016 ( 
.A(n_941),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_809),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_797),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_939),
.B(n_694),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_803),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_941),
.Y(n_1021)
);

AOI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_891),
.A2(n_369),
.B(n_364),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_939),
.B(n_694),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_915),
.A2(n_425),
.B(n_417),
.C(n_630),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_836),
.A2(n_417),
.B(n_541),
.C(n_543),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_872),
.A2(n_737),
.B(n_726),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_939),
.B(n_694),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_877),
.A2(n_890),
.B(n_879),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_803),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_793),
.B(n_889),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_869),
.B(n_694),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_876),
.A2(n_694),
.B1(n_410),
.B2(n_243),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_869),
.B(n_726),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_803),
.B(n_744),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_830),
.A2(n_737),
.B(n_744),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_798),
.A2(n_744),
.B(n_714),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_805),
.A2(n_920),
.B(n_916),
.Y(n_1037)
);

BUFx4f_ASAP7_75t_L g1038 ( 
.A(n_887),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_805),
.A2(n_744),
.B(n_714),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_924),
.A2(n_714),
.B(n_650),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_892),
.A2(n_714),
.B(n_650),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_893),
.A2(n_625),
.B(n_627),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_808),
.B(n_851),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_845),
.A2(n_648),
.B1(n_692),
.B2(n_689),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_794),
.A2(n_818),
.B(n_943),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_803),
.B(n_650),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_818),
.A2(n_692),
.B(n_689),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_838),
.A2(n_940),
.B1(n_904),
.B2(n_820),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_800),
.Y(n_1049)
);

AO21x1_ASAP7_75t_L g1050 ( 
.A1(n_828),
.A2(n_541),
.B(n_543),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_808),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_SL g1052 ( 
.A1(n_904),
.A2(n_546),
.B(n_630),
.C(n_625),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_915),
.A2(n_625),
.B(n_627),
.C(n_613),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_947),
.A2(n_627),
.B(n_585),
.C(n_613),
.Y(n_1054)
);

NOR3xp33_ASAP7_75t_L g1055 ( 
.A(n_960),
.B(n_407),
.C(n_336),
.Y(n_1055)
);

AOI22x1_ASAP7_75t_L g1056 ( 
.A1(n_918),
.A2(n_686),
.B1(n_684),
.B2(n_664),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_955),
.A2(n_692),
.B(n_689),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_851),
.B(n_650),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_929),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_900),
.A2(n_692),
.B(n_689),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_800),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_960),
.B(n_947),
.C(n_862),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_880),
.B(n_664),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_948),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_874),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_878),
.B(n_664),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_884),
.B(n_664),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_896),
.B(n_664),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_810),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_933),
.B(n_684),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_864),
.B(n_868),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_886),
.B(n_684),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_953),
.A2(n_585),
.B(n_610),
.C(n_613),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_957),
.A2(n_686),
.B(n_684),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_952),
.A2(n_686),
.B(n_684),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_811),
.A2(n_816),
.B(n_925),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_815),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_874),
.B(n_677),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_888),
.B(n_686),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_854),
.B(n_421),
.C(n_348),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_910),
.B(n_686),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_829),
.B(n_833),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_867),
.A2(n_697),
.B(n_558),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_829),
.B(n_599),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_867),
.A2(n_697),
.B(n_558),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_873),
.A2(n_697),
.B(n_558),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_873),
.A2(n_618),
.B(n_615),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_874),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_961),
.B(n_847),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_833),
.B(n_648),
.Y(n_1090)
);

AND2x2_ASAP7_75t_SL g1091 ( 
.A(n_834),
.B(n_546),
.Y(n_1091)
);

AO21x2_ASAP7_75t_L g1092 ( 
.A1(n_875),
.A2(n_618),
.B(n_615),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_822),
.A2(n_585),
.B(n_610),
.C(n_618),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_875),
.A2(n_697),
.B(n_550),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_948),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_931),
.A2(n_339),
.B(n_356),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_840),
.B(n_599),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_951),
.A2(n_697),
.B(n_550),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_840),
.B(n_599),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_930),
.A2(n_615),
.B(n_610),
.C(n_410),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_871),
.A2(n_418),
.B(n_370),
.C(n_374),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_923),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_951),
.B(n_648),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_811),
.A2(n_410),
.B(n_378),
.C(n_379),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_816),
.A2(n_603),
.B(n_601),
.C(n_599),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_887),
.B(n_363),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_936),
.A2(n_550),
.B(n_556),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_887),
.B(n_383),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_826),
.B(n_581),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_934),
.B(n_581),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_843),
.A2(n_550),
.B(n_556),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_894),
.A2(n_388),
.B(n_390),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_897),
.A2(n_556),
.B(n_550),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_937),
.B(n_581),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_946),
.B(n_581),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_856),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_898),
.A2(n_556),
.B(n_558),
.Y(n_1117)
);

NOR2x1_ASAP7_75t_L g1118 ( 
.A(n_848),
.B(n_945),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_SL g1119 ( 
.A(n_844),
.B(n_405),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_903),
.A2(n_556),
.B(n_558),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_906),
.A2(n_556),
.B(n_558),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_823),
.A2(n_430),
.B1(n_413),
.B2(n_419),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_856),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_860),
.B(n_586),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_912),
.A2(n_603),
.B(n_601),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_842),
.A2(n_426),
.B1(n_411),
.B2(n_599),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_919),
.A2(n_595),
.B1(n_586),
.B2(n_599),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_839),
.B(n_586),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_L g1129 ( 
.A1(n_913),
.A2(n_932),
.B(n_958),
.Y(n_1129)
);

BUFx4f_ASAP7_75t_L g1130 ( 
.A(n_949),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_860),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_914),
.A2(n_603),
.B1(n_601),
.B2(n_599),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_926),
.B(n_10),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_824),
.A2(n_10),
.B(n_12),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_881),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_L g1136 ( 
.A(n_850),
.B(n_13),
.C(n_16),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_911),
.A2(n_927),
.B(n_853),
.C(n_950),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_954),
.A2(n_595),
.B(n_586),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_881),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_885),
.A2(n_595),
.B(n_586),
.Y(n_1140)
);

NOR3xp33_ASAP7_75t_L g1141 ( 
.A(n_849),
.B(n_17),
.C(n_20),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_932),
.B(n_17),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_885),
.A2(n_595),
.B(n_586),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_895),
.B(n_595),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_931),
.B(n_595),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_956),
.B(n_944),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_863),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1087),
.A2(n_956),
.B(n_944),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_967),
.A2(n_942),
.B1(n_935),
.B2(n_928),
.Y(n_1149)
);

BUFx2_ASAP7_75t_SL g1150 ( 
.A(n_1021),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_995),
.B(n_895),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1049),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_996),
.B(n_901),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_971),
.A2(n_942),
.B(n_935),
.C(n_928),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_963),
.A2(n_922),
.B(n_921),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1011),
.A2(n_922),
.B(n_921),
.C(n_917),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1017),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_SL g1158 ( 
.A(n_1080),
.B(n_20),
.C(n_23),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1062),
.B(n_901),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1135),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1059),
.B(n_917),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_990),
.B(n_902),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_970),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1069),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1064),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_962),
.B(n_902),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_985),
.B(n_909),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_994),
.A2(n_908),
.B(n_907),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_962),
.Y(n_1169)
);

AND2x6_ASAP7_75t_SL g1170 ( 
.A(n_1030),
.B(n_1106),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_985),
.B(n_909),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1088),
.B(n_1030),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_976),
.B(n_907),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1062),
.B(n_908),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1089),
.A2(n_603),
.B(n_601),
.C(n_27),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1064),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_978),
.B(n_1089),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_969),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_L g1179 ( 
.A(n_1095),
.B(n_603),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1139),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1045),
.A2(n_603),
.B(n_601),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1131),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_966),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1055),
.A2(n_603),
.B1(n_601),
.B2(n_82),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_965),
.A2(n_601),
.B1(n_213),
.B2(n_211),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1071),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1064),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1022),
.B(n_23),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1064),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1037),
.A2(n_144),
.B(n_207),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_977),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1065),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_L g1193 ( 
.A(n_1055),
.B(n_209),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1010),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1147),
.A2(n_205),
.B1(n_191),
.B2(n_190),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1024),
.A2(n_30),
.B(n_33),
.C(n_35),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_SL g1197 ( 
.A(n_1006),
.B(n_186),
.Y(n_1197)
);

NOR3xp33_ASAP7_75t_L g1198 ( 
.A(n_979),
.B(n_36),
.C(n_37),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1091),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1071),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1002),
.A2(n_46),
.B(n_47),
.C(n_51),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_993),
.A2(n_92),
.B(n_182),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1139),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1049),
.B(n_86),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_997),
.A2(n_51),
.B(n_55),
.C(n_56),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1018),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1091),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_997),
.A2(n_110),
.B(n_175),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_973),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1018),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1116),
.Y(n_1211)
);

AND2x6_ASAP7_75t_SL g1212 ( 
.A(n_1030),
.B(n_60),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1005),
.B(n_65),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_R g1214 ( 
.A(n_1006),
.B(n_114),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_998),
.A2(n_119),
.B(n_167),
.Y(n_1215)
);

OAI21xp33_ASAP7_75t_SL g1216 ( 
.A1(n_984),
.A2(n_66),
.B(n_70),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1070),
.A2(n_66),
.B(n_70),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_999),
.A2(n_124),
.B(n_165),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1133),
.A2(n_72),
.B(n_73),
.C(n_75),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1000),
.A2(n_104),
.B(n_150),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_974),
.A2(n_103),
.B1(n_145),
.B2(n_141),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1077),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1133),
.A2(n_72),
.B(n_73),
.C(n_75),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1020),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1049),
.Y(n_1225)
);

CKINVDCx11_ASAP7_75t_R g1226 ( 
.A(n_1049),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_987),
.A2(n_125),
.B(n_133),
.Y(n_1227)
);

AO32x1_ASAP7_75t_L g1228 ( 
.A1(n_1126),
.A2(n_77),
.A3(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1061),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1035),
.A2(n_127),
.B(n_183),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1061),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_979),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1123),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1063),
.A2(n_1125),
.B(n_1068),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1142),
.A2(n_992),
.B(n_1137),
.C(n_1048),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_986),
.B(n_1145),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1051),
.B(n_1029),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1123),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1102),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1051),
.B(n_1029),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1142),
.A2(n_1054),
.B(n_1053),
.C(n_1136),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_1118),
.B1(n_1048),
.B2(n_1108),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1061),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1038),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1096),
.B(n_1106),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1082),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1146),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1129),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1136),
.A2(n_1141),
.B1(n_1050),
.B2(n_1122),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1066),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1130),
.A2(n_1043),
.B1(n_1061),
.B2(n_1070),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1130),
.B(n_1038),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1016),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1020),
.B(n_1095),
.Y(n_1254)
);

NOR3xp33_ASAP7_75t_SL g1255 ( 
.A(n_1108),
.B(n_1101),
.C(n_1112),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1033),
.B(n_1028),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_968),
.A2(n_980),
.B(n_964),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1007),
.A2(n_1015),
.B1(n_1019),
.B2(n_1013),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1100),
.A2(n_1009),
.B(n_1104),
.C(n_1076),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1078),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_988),
.A2(n_1012),
.B(n_981),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1141),
.A2(n_1073),
.B(n_1052),
.C(n_1025),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1067),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1072),
.B(n_1079),
.Y(n_1264)
);

BUFx8_ASAP7_75t_SL g1265 ( 
.A(n_1016),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1081),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1003),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1008),
.A2(n_1014),
.B(n_983),
.C(n_1027),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1134),
.A2(n_1023),
.B1(n_1032),
.B2(n_1128),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_975),
.A2(n_1063),
.B1(n_1068),
.B2(n_1031),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1058),
.A2(n_1046),
.B1(n_1001),
.B2(n_1034),
.Y(n_1271)
);

CKINVDCx16_ASAP7_75t_R g1272 ( 
.A(n_975),
.Y(n_1272)
);

AO32x1_ASAP7_75t_L g1273 ( 
.A1(n_1132),
.A2(n_1044),
.A3(n_1056),
.B1(n_1105),
.B2(n_1093),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1041),
.A2(n_989),
.B(n_1109),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1032),
.Y(n_1275)
);

OAI21xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1046),
.A2(n_1034),
.B(n_1001),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1103),
.B(n_1042),
.Y(n_1277)
);

INVx3_ASAP7_75t_SL g1278 ( 
.A(n_1084),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1075),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1092),
.B(n_1084),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1047),
.A2(n_1040),
.B(n_1039),
.C(n_1036),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1092),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_SL g1283 ( 
.A1(n_1097),
.A2(n_1099),
.B(n_1115),
.C(n_1114),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1097),
.B(n_1099),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1110),
.B(n_1090),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1124),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1057),
.B(n_1098),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1144),
.B(n_1026),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1074),
.A2(n_1094),
.B(n_1086),
.C(n_1083),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_SL g1290 ( 
.A(n_1107),
.B(n_1117),
.C(n_1121),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1060),
.B(n_1120),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1113),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1127),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_972),
.B(n_982),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1140),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_SL g1296 ( 
.A(n_1085),
.B(n_1138),
.C(n_1143),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1111),
.B(n_976),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_970),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_963),
.A2(n_859),
.B(n_1045),
.Y(n_1299)
);

NOR2x1_ASAP7_75t_L g1300 ( 
.A(n_1021),
.B(n_841),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_978),
.B(n_1049),
.Y(n_1301)
);

AOI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_967),
.A2(n_995),
.B(n_804),
.Y(n_1302)
);

XNOR2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1065),
.B(n_593),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1062),
.B(n_995),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1302),
.A2(n_1245),
.B(n_1235),
.C(n_1242),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1299),
.A2(n_1256),
.B(n_1261),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1239),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1299),
.A2(n_1261),
.B(n_1236),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1304),
.A2(n_1174),
.B(n_1241),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1169),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1186),
.B(n_1200),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1257),
.A2(n_1288),
.B(n_1279),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1186),
.B(n_1200),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1279),
.A2(n_1274),
.B(n_1287),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1177),
.B(n_1169),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1274),
.A2(n_1264),
.B(n_1171),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1151),
.B(n_1246),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1155),
.A2(n_1168),
.B(n_1234),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1291),
.A2(n_1248),
.B(n_1181),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_L g1321 ( 
.A(n_1255),
.B(n_1249),
.C(n_1207),
.Y(n_1321)
);

INVx5_ASAP7_75t_L g1322 ( 
.A(n_1265),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1259),
.A2(n_1268),
.A3(n_1282),
.B(n_1281),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1167),
.A2(n_1277),
.B(n_1153),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1182),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1226),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1225),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1289),
.A2(n_1285),
.B(n_1273),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1255),
.B(n_1199),
.C(n_1158),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1247),
.B(n_1162),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1154),
.A2(n_1156),
.B(n_1283),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1243),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_SL g1333 ( 
.A1(n_1208),
.A2(n_1219),
.B(n_1223),
.C(n_1175),
.Y(n_1333)
);

AOI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1159),
.A2(n_1271),
.B(n_1251),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1241),
.A2(n_1216),
.B(n_1270),
.C(n_1193),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1250),
.B(n_1263),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1154),
.A2(n_1156),
.B(n_1258),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1183),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1202),
.A2(n_1295),
.B(n_1230),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1266),
.B(n_1267),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1217),
.A2(n_1185),
.A3(n_1190),
.B(n_1230),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1190),
.A2(n_1290),
.B(n_1262),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1273),
.A2(n_1290),
.B(n_1292),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1269),
.A2(n_1213),
.B1(n_1161),
.B2(n_1211),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1163),
.B(n_1298),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1294),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1286),
.A2(n_1293),
.B(n_1215),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1262),
.A2(n_1280),
.B(n_1179),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1297),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1243),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1301),
.B(n_1252),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1237),
.A2(n_1240),
.B(n_1218),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1243),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1215),
.A2(n_1218),
.B(n_1227),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1220),
.A2(n_1227),
.B(n_1149),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1220),
.A2(n_1195),
.A3(n_1221),
.B(n_1222),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1233),
.A2(n_1238),
.B(n_1197),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1198),
.A2(n_1300),
.B1(n_1301),
.B2(n_1209),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1170),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1191),
.Y(n_1360)
);

OAI22x1_ASAP7_75t_L g1361 ( 
.A1(n_1232),
.A2(n_1244),
.B1(n_1203),
.B2(n_1180),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1184),
.A2(n_1205),
.B(n_1173),
.C(n_1201),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1194),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1198),
.A2(n_1205),
.B(n_1201),
.C(n_1196),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1206),
.A2(n_1210),
.B(n_1224),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1160),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1243),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1178),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1166),
.A2(n_1228),
.A3(n_1296),
.B(n_1196),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1178),
.A2(n_1209),
.B1(n_1192),
.B2(n_1272),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1260),
.B(n_1164),
.Y(n_1371)
);

OAI22x1_ASAP7_75t_L g1372 ( 
.A1(n_1278),
.A2(n_1253),
.B1(n_1204),
.B2(n_1284),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1284),
.B(n_1187),
.Y(n_1373)
);

AO31x2_ASAP7_75t_L g1374 ( 
.A1(n_1228),
.A2(n_1296),
.A3(n_1278),
.B(n_1158),
.Y(n_1374)
);

AOI221x1_ASAP7_75t_L g1375 ( 
.A1(n_1228),
.A2(n_1176),
.B1(n_1187),
.B2(n_1165),
.C(n_1189),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1224),
.A2(n_1150),
.B(n_1152),
.C(n_1229),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1254),
.A2(n_1165),
.B(n_1189),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1214),
.A2(n_1212),
.B1(n_1152),
.B2(n_1229),
.C(n_1231),
.Y(n_1378)
);

INVx5_ASAP7_75t_L g1379 ( 
.A(n_1165),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1172),
.B(n_1229),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1254),
.A2(n_1165),
.B(n_1189),
.Y(n_1381)
);

O2A1O1Ixp5_ASAP7_75t_L g1382 ( 
.A1(n_1254),
.A2(n_1172),
.B(n_1189),
.C(n_1231),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1303),
.A2(n_967),
.B(n_995),
.C(n_1302),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1231),
.B(n_899),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1242),
.B(n_1062),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1186),
.B(n_899),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1226),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1212),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1302),
.A2(n_967),
.B(n_995),
.C(n_1062),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1226),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1395)
);

OAI21xp33_ASAP7_75t_L g1396 ( 
.A1(n_1188),
.A2(n_967),
.B(n_995),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1302),
.A2(n_967),
.B(n_995),
.C(n_1062),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1301),
.B(n_1252),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1186),
.B(n_899),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1235),
.A2(n_967),
.B(n_1261),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1302),
.B(n_967),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1302),
.A2(n_967),
.B(n_995),
.C(n_1245),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1186),
.B(n_899),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_SL g1404 ( 
.A1(n_1235),
.A2(n_967),
.B(n_995),
.C(n_1302),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1163),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1265),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1265),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1302),
.B(n_995),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1235),
.A2(n_1259),
.A3(n_1268),
.B(n_1299),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1302),
.B(n_995),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_SL g1415 ( 
.A(n_1242),
.B(n_1062),
.C(n_995),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1235),
.A2(n_967),
.B1(n_995),
.B2(n_1186),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1164),
.Y(n_1417)
);

OAI22x1_ASAP7_75t_L g1418 ( 
.A1(n_1242),
.A2(n_1232),
.B1(n_1245),
.B2(n_1188),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1302),
.B(n_967),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1235),
.A2(n_967),
.B1(n_995),
.B2(n_1186),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1302),
.B(n_967),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1235),
.A2(n_967),
.B1(n_995),
.B2(n_1186),
.Y(n_1423)
);

AOI21xp33_ASAP7_75t_L g1424 ( 
.A1(n_1302),
.A2(n_967),
.B(n_995),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1302),
.B(n_967),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1302),
.A2(n_967),
.B(n_995),
.C(n_1245),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1427)
);

OAI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1235),
.A2(n_967),
.B1(n_995),
.B2(n_1186),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1163),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1302),
.B(n_967),
.Y(n_1431)
);

AOI221x1_ASAP7_75t_L g1432 ( 
.A1(n_1302),
.A2(n_967),
.B1(n_1062),
.B2(n_1198),
.C(n_1235),
.Y(n_1432)
);

CKINVDCx11_ASAP7_75t_R g1433 ( 
.A(n_1212),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1235),
.A2(n_1259),
.A3(n_1268),
.B(n_1299),
.Y(n_1434)
);

AO22x2_ASAP7_75t_L g1435 ( 
.A1(n_1198),
.A2(n_1062),
.B1(n_995),
.B2(n_967),
.Y(n_1435)
);

AO31x2_ASAP7_75t_L g1436 ( 
.A1(n_1235),
.A2(n_1259),
.A3(n_1268),
.B(n_1299),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1302),
.B(n_995),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1302),
.B(n_967),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1439)
);

AO31x2_ASAP7_75t_L g1440 ( 
.A1(n_1235),
.A2(n_1259),
.A3(n_1268),
.B(n_1299),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1261),
.A2(n_1235),
.B(n_1299),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1242),
.B(n_1062),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1261),
.A2(n_1235),
.B(n_1299),
.Y(n_1444)
);

AOI221x1_ASAP7_75t_L g1445 ( 
.A1(n_1302),
.A2(n_967),
.B1(n_1062),
.B2(n_1198),
.C(n_1235),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1212),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_SL g1450 ( 
.A1(n_1235),
.A2(n_967),
.B(n_995),
.C(n_1302),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1235),
.A2(n_967),
.B1(n_995),
.B2(n_1186),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1226),
.Y(n_1452)
);

NOR2x1p5_ASAP7_75t_L g1453 ( 
.A(n_1164),
.B(n_1021),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1257),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1302),
.B(n_967),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1157),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1245),
.A2(n_1062),
.B1(n_967),
.B2(n_995),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1226),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1302),
.B(n_967),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1299),
.A2(n_859),
.B(n_1256),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1406),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1321),
.A2(n_1437),
.B1(n_1412),
.B2(n_1414),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1321),
.A2(n_1458),
.B1(n_1358),
.B2(n_1305),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1430),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1409),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1459),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1417),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1329),
.A2(n_1445),
.B1(n_1432),
.B2(n_1418),
.Y(n_1469)
);

INVx6_ASAP7_75t_L g1470 ( 
.A(n_1379),
.Y(n_1470)
);

BUFx8_ASAP7_75t_L g1471 ( 
.A(n_1459),
.Y(n_1471)
);

INVx8_ASAP7_75t_L g1472 ( 
.A(n_1379),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1345),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1329),
.A2(n_1435),
.B1(n_1416),
.B2(n_1429),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1396),
.A2(n_1415),
.B1(n_1385),
.B2(n_1442),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1453),
.Y(n_1476)
);

BUFx10_ASAP7_75t_L g1477 ( 
.A(n_1459),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1435),
.A2(n_1451),
.B1(n_1423),
.B2(n_1420),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1327),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1327),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1416),
.A2(n_1423),
.B1(n_1451),
.B2(n_1420),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1379),
.B(n_1349),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1424),
.A2(n_1429),
.B1(n_1460),
.B2(n_1421),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1327),
.Y(n_1484)
);

INVx6_ASAP7_75t_L g1485 ( 
.A(n_1322),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1325),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1400),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1338),
.Y(n_1488)
);

BUFx10_ASAP7_75t_L g1489 ( 
.A(n_1326),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1401),
.A2(n_1431),
.B1(n_1460),
.B2(n_1425),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1424),
.A2(n_1431),
.B1(n_1438),
.B2(n_1421),
.Y(n_1491)
);

INVx6_ASAP7_75t_L g1492 ( 
.A(n_1322),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1318),
.A2(n_1426),
.B1(n_1402),
.B2(n_1370),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1401),
.A2(n_1425),
.B1(n_1438),
.B2(n_1455),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1318),
.A2(n_1335),
.B1(n_1383),
.B2(n_1340),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1400),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1340),
.A2(n_1419),
.B1(n_1455),
.B2(n_1336),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1351),
.A2(n_1398),
.B1(n_1378),
.B2(n_1371),
.Y(n_1498)
);

INVx6_ASAP7_75t_L g1499 ( 
.A(n_1322),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1419),
.A2(n_1359),
.B1(n_1349),
.B2(n_1310),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1452),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1457),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1363),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1310),
.A2(n_1316),
.B1(n_1410),
.B2(n_1351),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1380),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1410),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1312),
.A2(n_1344),
.B1(n_1378),
.B2(n_1403),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1344),
.A2(n_1388),
.B1(n_1399),
.B2(n_1336),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1314),
.A2(n_1441),
.B1(n_1444),
.B2(n_1330),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1314),
.A2(n_1441),
.B1(n_1444),
.B2(n_1330),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1368),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1390),
.A2(n_1449),
.B1(n_1433),
.B2(n_1372),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1332),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1323),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1343),
.A2(n_1355),
.B1(n_1360),
.B2(n_1324),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1366),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1311),
.A2(n_1328),
.B1(n_1347),
.B2(n_1342),
.Y(n_1518)
);

INVx3_ASAP7_75t_SL g1519 ( 
.A(n_1389),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1380),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1410),
.Y(n_1521)
);

INVx11_ASAP7_75t_L g1522 ( 
.A(n_1393),
.Y(n_1522)
);

BUFx4_ASAP7_75t_SL g1523 ( 
.A(n_1382),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1373),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1364),
.A2(n_1317),
.B1(n_1346),
.B2(n_1354),
.Y(n_1525)
);

BUFx4_ASAP7_75t_SL g1526 ( 
.A(n_1376),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1350),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1350),
.Y(n_1528)
);

INVx6_ASAP7_75t_L g1529 ( 
.A(n_1353),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1353),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1333),
.A2(n_1306),
.B1(n_1450),
.B2(n_1404),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1367),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1362),
.A2(n_1392),
.B1(n_1397),
.B2(n_1357),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1309),
.A2(n_1337),
.B1(n_1313),
.B2(n_1348),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1427),
.A2(n_1461),
.B1(n_1391),
.B2(n_1394),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1427),
.A2(n_1461),
.B1(n_1395),
.B2(n_1422),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1405),
.A2(n_1456),
.B1(n_1407),
.B2(n_1411),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1367),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1375),
.A2(n_1334),
.B1(n_1377),
.B2(n_1443),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1381),
.A2(n_1352),
.B1(n_1367),
.B2(n_1315),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1408),
.A2(n_1447),
.B1(n_1331),
.B2(n_1320),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1339),
.A2(n_1319),
.B1(n_1365),
.B2(n_1387),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1308),
.B(n_1428),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1323),
.Y(n_1544)
);

BUFx4_ASAP7_75t_R g1545 ( 
.A(n_1374),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1413),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1413),
.A2(n_1436),
.B1(n_1440),
.B2(n_1434),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1374),
.B(n_1356),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1374),
.A2(n_1436),
.B1(n_1440),
.B2(n_1434),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1413),
.Y(n_1550)
);

CKINVDCx11_ASAP7_75t_R g1551 ( 
.A(n_1356),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1436),
.A2(n_1440),
.B1(n_1369),
.B2(n_1341),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1369),
.A2(n_1341),
.B1(n_1356),
.B2(n_1386),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1439),
.A2(n_1446),
.B1(n_1448),
.B2(n_1454),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1369),
.B(n_1341),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_995),
.B2(n_1242),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1452),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1326),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_995),
.B2(n_1275),
.Y(n_1561)
);

CKINVDCx11_ASAP7_75t_R g1562 ( 
.A(n_1452),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1349),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1379),
.Y(n_1565)
);

BUFx8_ASAP7_75t_L g1566 ( 
.A(n_1459),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_995),
.B2(n_1242),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1418),
.A2(n_1062),
.B1(n_1245),
.B2(n_995),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1452),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1409),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1307),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1577)
);

BUFx4f_ASAP7_75t_L g1578 ( 
.A(n_1459),
.Y(n_1578)
);

BUFx8_ASAP7_75t_L g1579 ( 
.A(n_1459),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1313),
.A2(n_1461),
.B(n_1427),
.Y(n_1580)
);

OAI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_995),
.B2(n_1275),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1409),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_SL g1583 ( 
.A1(n_1321),
.A2(n_642),
.B(n_559),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1584)
);

CKINVDCx11_ASAP7_75t_R g1585 ( 
.A(n_1452),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1406),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_SL g1587 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1406),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_995),
.B2(n_1275),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1418),
.A2(n_1245),
.B1(n_1188),
.B2(n_1361),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1453),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1345),
.Y(n_1592)
);

BUFx4_ASAP7_75t_R g1593 ( 
.A(n_1406),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1418),
.A2(n_1062),
.B1(n_1245),
.B2(n_995),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1326),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1321),
.A2(n_693),
.B1(n_647),
.B2(n_1245),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1406),
.Y(n_1597)
);

INVx5_ASAP7_75t_L g1598 ( 
.A(n_1379),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1321),
.A2(n_967),
.B1(n_1414),
.B2(n_1412),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1550),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1494),
.B(n_1491),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1482),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1515),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1573),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1524),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1515),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1557),
.A2(n_1567),
.B(n_1569),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1546),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1546),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1580),
.A2(n_1543),
.B(n_1536),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1487),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1582),
.Y(n_1612)
);

INVx6_ASAP7_75t_L g1613 ( 
.A(n_1598),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1487),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1547),
.B(n_1533),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1496),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1563),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1491),
.B(n_1478),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1544),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1473),
.B(n_1592),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1555),
.B(n_1490),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1483),
.B(n_1474),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1463),
.B(n_1556),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1548),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1466),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1485),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1483),
.B(n_1481),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1552),
.Y(n_1628)
);

BUFx2_ASAP7_75t_SL g1629 ( 
.A(n_1598),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1485),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1552),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1502),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1509),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1560),
.B(n_1564),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1509),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1510),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1535),
.A2(n_1536),
.B(n_1537),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1539),
.A2(n_1554),
.B(n_1553),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1510),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1490),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1549),
.Y(n_1641)
);

INVx4_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1545),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1497),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1598),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1553),
.Y(n_1646)
);

AOI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1561),
.A2(n_1581),
.B(n_1589),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1503),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1511),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1508),
.B(n_1475),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1485),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1511),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1574),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1535),
.A2(n_1537),
.B(n_1542),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1568),
.B(n_1577),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1594),
.A2(n_1599),
.B(n_1556),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1551),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1501),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1505),
.B(n_1518),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1571),
.B(n_1572),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1472),
.Y(n_1661)
);

BUFx3_ASAP7_75t_L g1662 ( 
.A(n_1492),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1495),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1505),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1578),
.B(n_1559),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1518),
.B(n_1512),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1469),
.B(n_1493),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1492),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1492),
.B(n_1499),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1472),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1525),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1539),
.Y(n_1673)
);

AOI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1527),
.A2(n_1538),
.B(n_1517),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1587),
.B(n_1596),
.C(n_1599),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1593),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1516),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1516),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1540),
.Y(n_1679)
);

AOI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1486),
.A2(n_1488),
.B(n_1523),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1534),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1498),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1542),
.A2(n_1534),
.B(n_1541),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1541),
.Y(n_1684)
);

CKINVDCx11_ASAP7_75t_R g1685 ( 
.A(n_1558),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1571),
.B(n_1576),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1531),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1523),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1472),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1462),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1572),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1499),
.B(n_1506),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1575),
.A2(n_1576),
.B1(n_1584),
.B2(n_1583),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1507),
.B(n_1575),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1507),
.A2(n_1584),
.B(n_1513),
.Y(n_1695)
);

BUFx4f_ASAP7_75t_SL g1696 ( 
.A(n_1595),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1521),
.B(n_1590),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1561),
.A2(n_1589),
.B(n_1581),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1500),
.B(n_1504),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1588),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1526),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1513),
.A2(n_1526),
.B(n_1565),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1465),
.B(n_1597),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1499),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1528),
.A2(n_1532),
.B(n_1591),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1632),
.Y(n_1706)
);

AO32x2_ASAP7_75t_L g1707 ( 
.A1(n_1693),
.A2(n_1476),
.A3(n_1520),
.B1(n_1530),
.B2(n_1529),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1705),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1607),
.A2(n_1578),
.B(n_1597),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1647),
.A2(n_1586),
.B(n_1465),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1656),
.A2(n_1468),
.B(n_1479),
.C(n_1484),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1621),
.B(n_1467),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1579),
.C(n_1471),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1644),
.B(n_1514),
.Y(n_1714)
);

AO21x1_ASAP7_75t_L g1715 ( 
.A1(n_1634),
.A2(n_1470),
.B(n_1565),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1621),
.B(n_1519),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1667),
.B(n_1468),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1620),
.B(n_1625),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1685),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1675),
.A2(n_1480),
.B1(n_1479),
.B2(n_1519),
.C(n_1514),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1644),
.B(n_1470),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1655),
.A2(n_1585),
.B1(n_1570),
.B2(n_1562),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1643),
.B(n_1477),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_SL g1724 ( 
.A1(n_1701),
.A2(n_1471),
.B1(n_1566),
.B2(n_1579),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1602),
.B(n_1477),
.Y(n_1725)
);

A2O1A1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1695),
.A2(n_1566),
.B(n_1489),
.C(n_1529),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1617),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1602),
.B(n_1489),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1668),
.A2(n_1522),
.B(n_1666),
.C(n_1623),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1643),
.B(n_1601),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1604),
.B(n_1612),
.Y(n_1731)
);

AO21x2_ASAP7_75t_L g1732 ( 
.A1(n_1610),
.A2(n_1683),
.B(n_1654),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1664),
.B(n_1697),
.Y(n_1733)
);

AND2x6_ASAP7_75t_L g1734 ( 
.A(n_1663),
.B(n_1627),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1705),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1611),
.B(n_1614),
.Y(n_1736)
);

OA21x2_ASAP7_75t_L g1737 ( 
.A1(n_1683),
.A2(n_1654),
.B(n_1637),
.Y(n_1737)
);

OAI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1686),
.A2(n_1668),
.B(n_1695),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1663),
.B(n_1657),
.Y(n_1739)
);

OA21x2_ASAP7_75t_L g1740 ( 
.A1(n_1637),
.A2(n_1610),
.B(n_1673),
.Y(n_1740)
);

A2O1A1Ixp33_ASAP7_75t_L g1741 ( 
.A1(n_1627),
.A2(n_1622),
.B(n_1666),
.C(n_1694),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1660),
.A2(n_1691),
.B1(n_1650),
.B2(n_1618),
.C(n_1698),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_SL g1743 ( 
.A1(n_1679),
.A2(n_1691),
.B(n_1673),
.C(n_1640),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1614),
.B(n_1616),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1640),
.B(n_1649),
.Y(n_1745)
);

A2O1A1Ixp33_ASAP7_75t_L g1746 ( 
.A1(n_1694),
.A2(n_1618),
.B(n_1650),
.C(n_1660),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1615),
.A2(n_1677),
.B(n_1678),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1652),
.B(n_1616),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1698),
.A2(n_1615),
.B(n_1701),
.C(n_1682),
.Y(n_1749)
);

NAND2x1_ASAP7_75t_L g1750 ( 
.A(n_1705),
.B(n_1613),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1615),
.A2(n_1682),
.B1(n_1699),
.B2(n_1641),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1690),
.B(n_1700),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1652),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1674),
.Y(n_1754)
);

INVx3_ASAP7_75t_SL g1755 ( 
.A(n_1676),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1615),
.A2(n_1678),
.B(n_1677),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1648),
.Y(n_1757)
);

AO32x2_ASAP7_75t_L g1758 ( 
.A1(n_1651),
.A2(n_1669),
.A3(n_1642),
.B1(n_1631),
.B2(n_1628),
.Y(n_1758)
);

AO32x2_ASAP7_75t_L g1759 ( 
.A1(n_1651),
.A2(n_1669),
.A3(n_1642),
.B1(n_1631),
.B2(n_1628),
.Y(n_1759)
);

CKINVDCx6p67_ASAP7_75t_R g1760 ( 
.A(n_1658),
.Y(n_1760)
);

OR2x6_ASAP7_75t_L g1761 ( 
.A(n_1659),
.B(n_1629),
.Y(n_1761)
);

NAND2x1_ASAP7_75t_L g1762 ( 
.A(n_1613),
.B(n_1670),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1699),
.A2(n_1702),
.B(n_1688),
.C(n_1672),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1670),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1698),
.A2(n_1687),
.B(n_1688),
.C(n_1684),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1681),
.A2(n_1679),
.B(n_1646),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1703),
.B(n_1665),
.Y(n_1767)
);

INVx5_ASAP7_75t_L g1768 ( 
.A(n_1645),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1638),
.A2(n_1681),
.B(n_1659),
.Y(n_1769)
);

OAI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1680),
.A2(n_1702),
.B(n_1633),
.Y(n_1770)
);

XNOR2xp5_ASAP7_75t_L g1771 ( 
.A(n_1626),
.B(n_1630),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1605),
.B(n_1641),
.Y(n_1772)
);

AO32x2_ASAP7_75t_L g1773 ( 
.A1(n_1642),
.A2(n_1671),
.A3(n_1661),
.B1(n_1689),
.B2(n_1646),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1761),
.B(n_1609),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1633),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1706),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1735),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1766),
.B(n_1635),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1757),
.Y(n_1779)
);

NOR2x1p5_ASAP7_75t_L g1780 ( 
.A(n_1713),
.B(n_1630),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_L g1781 ( 
.A(n_1734),
.B(n_1613),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1708),
.B(n_1638),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1742),
.B(n_1635),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1737),
.B(n_1636),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1754),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1708),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1742),
.A2(n_1741),
.B1(n_1746),
.B2(n_1722),
.C(n_1720),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1730),
.B(n_1639),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1769),
.B(n_1603),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1740),
.B(n_1600),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1727),
.B(n_1603),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1769),
.B(n_1606),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1727),
.B(n_1606),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1758),
.B(n_1608),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1753),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1748),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1748),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1736),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1744),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1758),
.B(n_1759),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1768),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1772),
.B(n_1624),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1772),
.B(n_1624),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1773),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1747),
.B(n_1659),
.Y(n_1805)
);

BUFx3_ASAP7_75t_L g1806 ( 
.A(n_1750),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1747),
.B(n_1659),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1745),
.B(n_1738),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1758),
.B(n_1619),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1759),
.B(n_1619),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1759),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1745),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1732),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1713),
.A2(n_1734),
.B1(n_1715),
.B2(n_1720),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1738),
.B(n_1653),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1714),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1808),
.B(n_1752),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1785),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_L g1819 ( 
.A1(n_1787),
.A2(n_1709),
.B(n_1710),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1801),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1787),
.B(n_1716),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1808),
.B(n_1756),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1798),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1786),
.B(n_1756),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1790),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1809),
.B(n_1733),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1809),
.B(n_1773),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1814),
.A2(n_1711),
.B1(n_1726),
.B2(n_1709),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1786),
.B(n_1732),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1809),
.B(n_1773),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1806),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1810),
.B(n_1717),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_1783),
.B(n_1765),
.C(n_1729),
.Y(n_1833)
);

OR2x2_ASAP7_75t_SL g1834 ( 
.A(n_1783),
.B(n_1712),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1804),
.B(n_1788),
.Y(n_1835)
);

INVxp67_ASAP7_75t_SL g1836 ( 
.A(n_1812),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1816),
.B(n_1765),
.Y(n_1837)
);

OAI33xp33_ASAP7_75t_L g1838 ( 
.A1(n_1802),
.A2(n_1751),
.A3(n_1714),
.B1(n_1721),
.B2(n_1749),
.B3(n_1739),
.Y(n_1838)
);

OAI211xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1815),
.A2(n_1729),
.B(n_1749),
.C(n_1763),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1775),
.B(n_1770),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1776),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1815),
.B(n_1710),
.C(n_1751),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1812),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1776),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1796),
.B(n_1721),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1782),
.B(n_1743),
.C(n_1770),
.Y(n_1846)
);

BUFx2_ASAP7_75t_L g1847 ( 
.A(n_1806),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1799),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1790),
.Y(n_1849)
);

AOI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1800),
.A2(n_1719),
.B(n_1724),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1799),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1806),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1780),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1782),
.A2(n_1762),
.B(n_1767),
.C(n_1723),
.Y(n_1854)
);

AND4x1_ASAP7_75t_L g1855 ( 
.A(n_1800),
.B(n_1731),
.C(n_1718),
.D(n_1760),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1775),
.B(n_1764),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1779),
.Y(n_1857)
);

AOI211xp5_ASAP7_75t_L g1858 ( 
.A1(n_1805),
.A2(n_1807),
.B(n_1789),
.C(n_1792),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1789),
.A2(n_1692),
.B1(n_1707),
.B2(n_1771),
.C(n_1662),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1779),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1801),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1848),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1827),
.B(n_1830),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1811),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1825),
.B(n_1801),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1830),
.B(n_1811),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1811),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1840),
.B(n_1778),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1837),
.B(n_1836),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1849),
.B(n_1801),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1840),
.B(n_1778),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1835),
.B(n_1784),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1851),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1858),
.B(n_1784),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1843),
.B(n_1818),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1820),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1821),
.B(n_1728),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1857),
.Y(n_1878)
);

HB1xp67_ASAP7_75t_L g1879 ( 
.A(n_1823),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1858),
.B(n_1832),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1832),
.B(n_1784),
.Y(n_1882)
);

AND2x4_ASAP7_75t_SL g1883 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1820),
.B(n_1774),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1841),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1829),
.Y(n_1886)
);

OAI33xp33_ASAP7_75t_L g1887 ( 
.A1(n_1833),
.A2(n_1791),
.A3(n_1793),
.B1(n_1803),
.B2(n_1802),
.B3(n_1795),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1841),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1826),
.B(n_1794),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1829),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1844),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1844),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1856),
.B(n_1777),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1860),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1818),
.B(n_1797),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1880),
.B(n_1831),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1883),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1887),
.A2(n_1819),
.B1(n_1833),
.B2(n_1839),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1880),
.B(n_1831),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1869),
.B(n_1845),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1878),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1895),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1880),
.B(n_1847),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1877),
.B(n_1658),
.Y(n_1905)
);

CKINVDCx16_ASAP7_75t_R g1906 ( 
.A(n_1881),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1895),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1868),
.B(n_1834),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1885),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1885),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1885),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1888),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1888),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1878),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1869),
.B(n_1822),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1888),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1891),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1879),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1878),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1874),
.B(n_1822),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1878),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1868),
.B(n_1834),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1874),
.B(n_1817),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1875),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1863),
.B(n_1847),
.Y(n_1925)
);

NAND2x1p5_ASAP7_75t_L g1926 ( 
.A(n_1876),
.B(n_1781),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1884),
.B(n_1696),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1892),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1891),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1868),
.B(n_1856),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1891),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1894),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1894),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1894),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1883),
.Y(n_1935)
);

NOR2x1p5_ASAP7_75t_SL g1936 ( 
.A(n_1886),
.B(n_1813),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1879),
.Y(n_1937)
);

NAND2x1p5_ASAP7_75t_L g1938 ( 
.A(n_1876),
.B(n_1861),
.Y(n_1938)
);

NOR3x1_ASAP7_75t_L g1939 ( 
.A(n_1876),
.B(n_1854),
.C(n_1828),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1862),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1863),
.B(n_1852),
.Y(n_1941)
);

AOI22xp33_ASAP7_75t_L g1942 ( 
.A1(n_1887),
.A2(n_1819),
.B1(n_1842),
.B2(n_1838),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1863),
.B(n_1852),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1862),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1892),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1892),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1909),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1898),
.B(n_1863),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1925),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1874),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1925),
.B(n_1884),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1909),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1941),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1938),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1908),
.B(n_1871),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1941),
.B(n_1884),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1943),
.B(n_1881),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1908),
.B(n_1871),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1943),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1910),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1906),
.B(n_1884),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1922),
.B(n_1871),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_L g1963 ( 
.A1(n_1904),
.A2(n_1842),
.B1(n_1846),
.B2(n_1850),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1896),
.B(n_1889),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1910),
.Y(n_1965)
);

NAND2x1_ASAP7_75t_L g1966 ( 
.A(n_1897),
.B(n_1884),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1922),
.B(n_1893),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1940),
.B(n_1864),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1911),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1896),
.B(n_1884),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1899),
.B(n_1883),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1911),
.Y(n_1972)
);

XNOR2x1_ASAP7_75t_L g1973 ( 
.A(n_1899),
.B(n_1846),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1928),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1928),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1912),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1912),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1903),
.B(n_1883),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1903),
.B(n_1889),
.Y(n_1979)
);

INVx2_ASAP7_75t_SL g1980 ( 
.A(n_1938),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1926),
.B(n_1889),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1913),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1926),
.B(n_1889),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1937),
.B(n_1893),
.Y(n_1984)
);

INVxp33_ASAP7_75t_L g1985 ( 
.A(n_1905),
.Y(n_1985)
);

NAND2x1p5_ASAP7_75t_L g1986 ( 
.A(n_1939),
.B(n_1855),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1947),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1986),
.A2(n_1859),
.B1(n_1850),
.B2(n_1935),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1985),
.B(n_1927),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1948),
.B(n_1918),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1986),
.A2(n_1938),
.B(n_1926),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1986),
.A2(n_1973),
.B1(n_1963),
.B2(n_1950),
.Y(n_1992)
);

OAI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1986),
.A2(n_1855),
.B1(n_1920),
.B2(n_1937),
.C(n_1915),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1973),
.A2(n_1853),
.B1(n_1897),
.B2(n_1780),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1963),
.A2(n_1944),
.B(n_1900),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1947),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1948),
.B(n_1950),
.Y(n_1997)
);

OAI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1973),
.A2(n_1923),
.B1(n_1881),
.B2(n_1944),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1952),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1949),
.B(n_1924),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1964),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1966),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1952),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1961),
.A2(n_1881),
.B1(n_1734),
.B2(n_1902),
.Y(n_2004)
);

OAI33xp33_ASAP7_75t_L g2005 ( 
.A1(n_1984),
.A2(n_1907),
.A3(n_1931),
.B1(n_1934),
.B2(n_1933),
.B3(n_1932),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1960),
.Y(n_2006)
);

O2A1O1Ixp5_ASAP7_75t_L g2007 ( 
.A1(n_1954),
.A2(n_1966),
.B(n_1949),
.C(n_1959),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1967),
.B(n_1930),
.Y(n_2008)
);

AOI222xp33_ASAP7_75t_L g2009 ( 
.A1(n_1968),
.A2(n_1936),
.B1(n_1873),
.B2(n_1907),
.C1(n_1864),
.C2(n_1866),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1971),
.Y(n_2010)
);

CKINVDCx14_ASAP7_75t_R g2011 ( 
.A(n_1971),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1960),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1965),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1949),
.B(n_1873),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1964),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1992),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1987),
.Y(n_2017)
);

OAI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1995),
.A2(n_1968),
.B1(n_1967),
.B2(n_1955),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_1995),
.B(n_1954),
.Y(n_2019)
);

CKINVDCx16_ASAP7_75t_R g2020 ( 
.A(n_2011),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1997),
.A2(n_1980),
.B(n_1961),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1990),
.B(n_1955),
.Y(n_2022)
);

OAI211xp5_ASAP7_75t_L g2023 ( 
.A1(n_1993),
.A2(n_1954),
.B(n_1980),
.C(n_1962),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2002),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2010),
.B(n_1953),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_2001),
.Y(n_2026)
);

AOI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1993),
.A2(n_1959),
.B1(n_1953),
.B2(n_1964),
.C(n_1957),
.Y(n_2027)
);

AOI21xp33_ASAP7_75t_L g2028 ( 
.A1(n_1989),
.A2(n_1980),
.B(n_1954),
.Y(n_2028)
);

AOI21xp33_ASAP7_75t_L g2029 ( 
.A1(n_1998),
.A2(n_1962),
.B(n_1958),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1996),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1999),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_2015),
.B(n_1978),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1991),
.B(n_1957),
.Y(n_2033)
);

O2A1O1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1988),
.A2(n_1958),
.B(n_1984),
.C(n_1959),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_2008),
.B(n_2014),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2000),
.B(n_1953),
.Y(n_2036)
);

OAI211xp5_ASAP7_75t_SL g2037 ( 
.A1(n_2009),
.A2(n_1965),
.B(n_1972),
.C(n_1969),
.Y(n_2037)
);

OAI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1994),
.A2(n_1824),
.B1(n_1881),
.B2(n_1930),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2026),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_2016),
.A2(n_1978),
.B1(n_2004),
.B2(n_2005),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_2020),
.B(n_2007),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2017),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_2019),
.Y(n_2043)
);

OAI21xp5_ASAP7_75t_SL g2044 ( 
.A1(n_2016),
.A2(n_1957),
.B(n_1970),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_2024),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2018),
.A2(n_2005),
.B1(n_2007),
.B2(n_2012),
.C(n_2006),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2032),
.B(n_1970),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2030),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2031),
.Y(n_2049)
);

NAND2x1p5_ASAP7_75t_L g2050 ( 
.A(n_2033),
.B(n_2022),
.Y(n_2050)
);

AOI211xp5_ASAP7_75t_L g2051 ( 
.A1(n_2018),
.A2(n_2023),
.B(n_2034),
.C(n_2027),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2025),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_2041),
.B(n_2035),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_2051),
.B(n_2028),
.C(n_2021),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_2045),
.B(n_2036),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_2043),
.A2(n_2037),
.B(n_2029),
.Y(n_2056)
);

NAND4xp25_ASAP7_75t_L g2057 ( 
.A(n_2040),
.B(n_2037),
.C(n_2003),
.D(n_2013),
.Y(n_2057)
);

NOR3xp33_ASAP7_75t_L g2058 ( 
.A(n_2043),
.B(n_2038),
.C(n_1957),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_2052),
.B(n_2044),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_2050),
.B(n_2038),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_1755),
.Y(n_2061)
);

NAND2x1_ASAP7_75t_L g2062 ( 
.A(n_2047),
.B(n_1983),
.Y(n_2062)
);

NAND4xp25_ASAP7_75t_L g2063 ( 
.A(n_2046),
.B(n_1983),
.C(n_1981),
.D(n_1951),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_2039),
.B(n_1951),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_SL g2065 ( 
.A(n_2042),
.B(n_1972),
.C(n_1969),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_2048),
.A2(n_1983),
.B(n_1981),
.Y(n_2066)
);

AOI32xp33_ASAP7_75t_L g2067 ( 
.A1(n_2049),
.A2(n_1956),
.A3(n_1979),
.B1(n_1977),
.B2(n_1976),
.Y(n_2067)
);

OAI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_2056),
.A2(n_1982),
.B1(n_1977),
.B2(n_1976),
.C(n_1956),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2055),
.Y(n_2069)
);

NAND3xp33_ASAP7_75t_SL g2070 ( 
.A(n_2060),
.B(n_1979),
.C(n_1982),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2054),
.A2(n_2057),
.B1(n_2058),
.B2(n_2063),
.C(n_2059),
.Y(n_2071)
);

AOI32xp33_ASAP7_75t_L g2072 ( 
.A1(n_2064),
.A2(n_1975),
.A3(n_1974),
.B1(n_1870),
.B2(n_1865),
.Y(n_2072)
);

AOI221x1_ASAP7_75t_L g2073 ( 
.A1(n_2061),
.A2(n_1975),
.B1(n_1974),
.B2(n_1913),
.C(n_1931),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2062),
.Y(n_2074)
);

OR2x2_ASAP7_75t_L g2075 ( 
.A(n_2070),
.B(n_2053),
.Y(n_2075)
);

AOI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_2071),
.A2(n_2066),
.B(n_2065),
.C(n_2067),
.Y(n_2076)
);

AOI211xp5_ASAP7_75t_L g2077 ( 
.A1(n_2068),
.A2(n_1975),
.B(n_1974),
.C(n_1728),
.Y(n_2077)
);

OAI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_2074),
.A2(n_1861),
.B(n_1921),
.C(n_1919),
.Y(n_2078)
);

AOI21xp33_ASAP7_75t_L g2079 ( 
.A1(n_2069),
.A2(n_1914),
.B(n_1901),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2073),
.Y(n_2080)
);

CKINVDCx20_ASAP7_75t_R g2081 ( 
.A(n_2072),
.Y(n_2081)
);

CKINVDCx20_ASAP7_75t_R g2082 ( 
.A(n_2069),
.Y(n_2082)
);

NAND4xp75_ASAP7_75t_L g2083 ( 
.A(n_2080),
.B(n_2079),
.C(n_2082),
.D(n_2076),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2075),
.Y(n_2084)
);

XNOR2xp5_ASAP7_75t_L g2085 ( 
.A(n_2081),
.B(n_1725),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2078),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2077),
.B(n_1882),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_2082),
.A2(n_1881),
.B1(n_1901),
.B2(n_1914),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2080),
.B(n_1916),
.Y(n_2089)
);

AOI322xp5_ASAP7_75t_L g2090 ( 
.A1(n_2084),
.A2(n_1864),
.A3(n_1866),
.B1(n_1867),
.B2(n_1886),
.C1(n_1890),
.C2(n_1872),
.Y(n_2090)
);

NAND3x1_ASAP7_75t_L g2091 ( 
.A(n_2089),
.B(n_1917),
.C(n_1916),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2085),
.Y(n_2092)
);

AOI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_2083),
.A2(n_1881),
.B1(n_1917),
.B2(n_1934),
.Y(n_2093)
);

AOI221xp5_ASAP7_75t_SL g2094 ( 
.A1(n_2086),
.A2(n_1933),
.B1(n_1932),
.B2(n_1929),
.C(n_1919),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2093),
.A2(n_2088),
.B1(n_2089),
.B2(n_2087),
.Y(n_2095)
);

XNOR2x1_ASAP7_75t_SL g2096 ( 
.A(n_2092),
.B(n_1929),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_SL g2097 ( 
.A1(n_2095),
.A2(n_2091),
.B1(n_2094),
.B2(n_1881),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2097),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_SL g2099 ( 
.A1(n_2097),
.A2(n_2096),
.B1(n_2090),
.B2(n_1921),
.Y(n_2099)
);

AOI22x1_ASAP7_75t_L g2100 ( 
.A1(n_2098),
.A2(n_1945),
.B1(n_1946),
.B2(n_1890),
.Y(n_2100)
);

NOR2x1p5_ASAP7_75t_L g2101 ( 
.A(n_2099),
.B(n_1630),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2101),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2100),
.B(n_1886),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2102),
.B(n_1886),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2104),
.A2(n_2103),
.B(n_1946),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2105),
.Y(n_2106)
);

OAI221xp5_ASAP7_75t_R g2107 ( 
.A1(n_2106),
.A2(n_1936),
.B1(n_1945),
.B2(n_1890),
.C(n_1875),
.Y(n_2107)
);

AOI211xp5_ASAP7_75t_L g2108 ( 
.A1(n_2107),
.A2(n_1704),
.B(n_1662),
.C(n_1890),
.Y(n_2108)
);


endmodule