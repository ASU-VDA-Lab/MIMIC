module real_aes_15320_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_87;
wire n_171;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx2_ASAP7_75t_SL g262 ( .A(n_0), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_1), .Y(n_123) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_2), .A2(n_42), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g164 ( .A(n_2), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_3), .B(n_154), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_4), .B(n_273), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_5), .A2(n_529), .B1(n_709), .B2(n_710), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_5), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_6), .A2(n_35), .B1(n_629), .B2(n_630), .Y(n_628) );
INVxp33_ASAP7_75t_SL g644 ( .A(n_6), .Y(n_644) );
AND2x2_ASAP7_75t_L g166 ( .A(n_7), .B(n_134), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_8), .B(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g540 ( .A(n_9), .Y(n_540) );
OAI222xp33_ASAP7_75t_L g659 ( .A1(n_10), .A2(n_48), .B1(n_55), .B2(n_576), .C1(n_660), .C2(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g683 ( .A(n_10), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_11), .A2(n_28), .B1(n_556), .B2(n_560), .Y(n_555) );
INVx1_ASAP7_75t_L g603 ( .A(n_11), .Y(n_603) );
INVx3_ASAP7_75t_L g535 ( .A(n_12), .Y(n_535) );
INVx1_ASAP7_75t_L g742 ( .A(n_13), .Y(n_742) );
INVx1_ASAP7_75t_L g747 ( .A(n_14), .Y(n_747) );
INVx1_ASAP7_75t_L g547 ( .A(n_15), .Y(n_547) );
INVx2_ASAP7_75t_L g553 ( .A(n_15), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_16), .B(n_129), .Y(n_202) );
INVx1_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
BUFx3_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_18), .B(n_133), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_19), .A2(n_64), .B1(n_580), .B2(n_584), .Y(n_579) );
INVxp33_ASAP7_75t_SL g700 ( .A(n_19), .Y(n_700) );
BUFx10_ASAP7_75t_L g722 ( .A(n_20), .Y(n_722) );
INVx1_ASAP7_75t_L g578 ( .A(n_21), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_22), .Y(n_196) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_23), .B(n_114), .C(n_276), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_24), .B(n_239), .Y(n_238) );
INVxp33_ASAP7_75t_L g595 ( .A(n_25), .Y(n_595) );
INVx1_ASAP7_75t_L g620 ( .A(n_25), .Y(n_620) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_25), .Y(n_707) );
INVx1_ASAP7_75t_L g85 ( .A(n_26), .Y(n_85) );
INVx2_ASAP7_75t_L g602 ( .A(n_27), .Y(n_602) );
INVxp33_ASAP7_75t_SL g697 ( .A(n_28), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_29), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g654 ( .A(n_30), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g675 ( .A1(n_30), .A2(n_676), .B(n_678), .C(n_690), .Y(n_675) );
INVxp67_ASAP7_75t_SL g548 ( .A(n_31), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_31), .A2(n_52), .B1(n_611), .B2(n_614), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_32), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g594 ( .A(n_33), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_33), .B(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_33), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_34), .B(n_127), .Y(n_126) );
INVxp33_ASAP7_75t_SL g650 ( .A(n_35), .Y(n_650) );
AND2x4_ASAP7_75t_L g84 ( .A(n_36), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_36), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_37), .B(n_133), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_38), .B(n_230), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_39), .B(n_133), .Y(n_292) );
INVx1_ASAP7_75t_L g546 ( .A(n_40), .Y(n_546) );
INVx1_ASAP7_75t_L g559 ( .A(n_40), .Y(n_559) );
INVx1_ASAP7_75t_L g744 ( .A(n_41), .Y(n_744) );
INVx1_ASAP7_75t_L g163 ( .A(n_42), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_43), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_44), .A2(n_153), .B(n_260), .C(n_263), .Y(n_259) );
INVx1_ASAP7_75t_L g733 ( .A(n_44), .Y(n_733) );
INVx1_ASAP7_75t_L g623 ( .A(n_45), .Y(n_623) );
INVx1_ASAP7_75t_L g110 ( .A(n_46), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_47), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g686 ( .A(n_48), .Y(n_686) );
INVx3_ASAP7_75t_L g193 ( .A(n_49), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_50), .B(n_189), .Y(n_301) );
INVx1_ASAP7_75t_L g205 ( .A(n_51), .Y(n_205) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_52), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_53), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_54), .B(n_118), .Y(n_271) );
INVx1_ASAP7_75t_L g627 ( .A(n_55), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_56), .B(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_57), .A2(n_68), .B1(n_750), .B2(n_751), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_57), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_58), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g254 ( .A(n_59), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_59), .A2(n_254), .B1(n_529), .B2(n_710), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_60), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_61), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_62), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
BUFx3_ASAP7_75t_L g129 ( .A(n_63), .Y(n_129) );
INVx1_ASAP7_75t_L g159 ( .A(n_63), .Y(n_159) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_64), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_65), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g191 ( .A(n_66), .Y(n_191) );
INVx2_ASAP7_75t_L g601 ( .A(n_67), .Y(n_601) );
AND2x2_ASAP7_75t_L g613 ( .A(n_67), .B(n_602), .Y(n_613) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_67), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_68), .B(n_145), .Y(n_244) );
INVx1_ASAP7_75t_L g750 ( .A(n_68), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_69), .B(n_134), .Y(n_247) );
INVx2_ASAP7_75t_L g538 ( .A(n_70), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_71), .B(n_91), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_72), .Y(n_183) );
INVx1_ASAP7_75t_L g178 ( .A(n_73), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_74), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_75), .B(n_189), .Y(n_295) );
INVx1_ASAP7_75t_L g554 ( .A(n_76), .Y(n_554) );
OAI21xp33_ASAP7_75t_SL g694 ( .A1(n_76), .A2(n_695), .B(n_696), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_95), .B(n_518), .Y(n_77) );
BUFx6f_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
NOR2xp33_ASAP7_75t_L g79 ( .A(n_80), .B(n_86), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
AO31x2_ASAP7_75t_L g137 ( .A1(n_81), .A2(n_138), .A3(n_160), .B(n_166), .Y(n_137) );
AO31x2_ASAP7_75t_L g336 ( .A1(n_81), .A2(n_138), .A3(n_160), .B(n_166), .Y(n_336) );
BUFx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
OAI21xp33_ASAP7_75t_L g264 ( .A1(n_83), .A2(n_161), .B(n_258), .Y(n_264) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx2_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVx3_ASAP7_75t_L g181 ( .A(n_84), .Y(n_181) );
BUFx6f_ASAP7_75t_SL g212 ( .A(n_84), .Y(n_212) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_85), .Y(n_525) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_86), .A2(n_524), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AOI22x1_ASAP7_75t_L g139 ( .A1(n_88), .A2(n_140), .B1(n_149), .B2(n_156), .Y(n_139) );
INVx1_ASAP7_75t_L g263 ( .A(n_88), .Y(n_263) );
AOI21x1_ASAP7_75t_L g270 ( .A1(n_88), .A2(n_271), .B(n_272), .Y(n_270) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g121 ( .A(n_89), .Y(n_121) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
INVx2_ASAP7_75t_L g154 ( .A(n_93), .Y(n_154) );
INVx2_ASAP7_75t_L g298 ( .A(n_93), .Y(n_298) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_416), .Y(n_98) );
NOR3xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_338), .C(n_389), .Y(n_99) );
OAI221xp5_ASAP7_75t_SL g100 ( .A1(n_101), .A2(n_232), .B1(n_280), .B2(n_285), .C(n_307), .Y(n_100) );
AOI211xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_167), .B(n_214), .C(n_222), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g513 ( .A(n_103), .B(n_218), .Y(n_513) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_136), .Y(n_103) );
INVx1_ASAP7_75t_L g216 ( .A(n_104), .Y(n_216) );
AND2x2_ASAP7_75t_L g368 ( .A(n_104), .B(n_314), .Y(n_368) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_104), .Y(n_413) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g225 ( .A(n_105), .Y(n_225) );
INVx3_ASAP7_75t_L g316 ( .A(n_105), .Y(n_316) );
AND2x2_ASAP7_75t_L g344 ( .A(n_105), .B(n_227), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_105), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI21x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_111), .B(n_132), .Y(n_106) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_107), .A2(n_199), .B(n_213), .Y(n_198) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_109), .Y(n_230) );
INVx1_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_122), .B(n_130), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_120), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g207 ( .A(n_115), .Y(n_207) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_116), .Y(n_119) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_116), .Y(n_185) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx3_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_119), .Y(n_151) );
INVx2_ASAP7_75t_L g239 ( .A(n_119), .Y(n_239) );
INVx3_ASAP7_75t_L g253 ( .A(n_119), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_120), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_120), .A2(n_244), .B(n_245), .Y(n_243) );
BUFx10_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g276 ( .A(n_121), .Y(n_276) );
O2A1O1Ixp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B(n_126), .C(n_128), .Y(n_122) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_129), .B(n_181), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g190 ( .A(n_129), .B(n_181), .C(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g206 ( .A(n_129), .Y(n_206) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_130), .A2(n_270), .B(n_274), .Y(n_269) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g305 ( .A(n_131), .Y(n_305) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_133), .Y(n_268) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g325 ( .A(n_137), .B(n_284), .Y(n_325) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_139), .A2(n_228), .B(n_231), .Y(n_227) );
OAI22x1_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_143), .B1(n_144), .B2(n_148), .Y(n_140) );
INVxp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g241 ( .A(n_146), .Y(n_241) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_146), .Y(n_256) );
INVx2_ASAP7_75t_L g273 ( .A(n_146), .Y(n_273) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B1(n_153), .B2(n_155), .Y(n_149) );
INVxp67_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVxp67_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21x1_ASAP7_75t_SL g251 ( .A1(n_156), .A2(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_157), .A2(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx3_ASAP7_75t_L g242 ( .A(n_159), .Y(n_242) );
INVxp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_162) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_163), .A2(n_164), .B(n_165), .Y(n_174) );
INVx1_ASAP7_75t_L g231 ( .A(n_166), .Y(n_231) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_168), .A2(n_340), .A3(n_344), .B1(n_345), .B2(n_348), .C1(n_355), .C2(n_363), .Y(n_339) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g363 ( .A(n_170), .B(n_315), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_170), .B(n_315), .Y(n_378) );
AND2x2_ASAP7_75t_L g431 ( .A(n_170), .B(n_344), .Y(n_431) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_197), .Y(n_170) );
INVx3_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_195), .Y(n_171) );
AO21x1_ASAP7_75t_L g353 ( .A1(n_172), .A2(n_175), .B(n_195), .Y(n_353) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g195 ( .A(n_173), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_188), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B1(n_182), .B2(n_186), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
INVx2_ASAP7_75t_L g246 ( .A(n_179), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_181), .B(n_187), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g192 ( .A(n_181), .B(n_187), .C(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
INVx2_ASAP7_75t_L g189 ( .A(n_184), .Y(n_189) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g211 ( .A(n_185), .Y(n_211) );
INVx2_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B1(n_192), .B2(n_194), .Y(n_188) );
INVx1_ASAP7_75t_L g221 ( .A(n_197), .Y(n_221) );
AND2x2_ASAP7_75t_L g226 ( .A(n_197), .B(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g284 ( .A(n_197), .Y(n_284) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_197), .Y(n_373) );
INVx2_ASAP7_75t_L g386 ( .A(n_197), .Y(n_386) );
AND2x2_ASAP7_75t_L g396 ( .A(n_197), .B(n_220), .Y(n_396) );
INVx1_ASAP7_75t_L g457 ( .A(n_197), .Y(n_457) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_208), .B(n_212), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_203), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_207), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_212), .A2(n_237), .B(n_243), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g474 ( .A(n_216), .Y(n_474) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g500 ( .A(n_219), .B(n_335), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g314 ( .A(n_220), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_220), .B(n_316), .Y(n_337) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_224), .B(n_226), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_224), .B(n_422), .Y(n_446) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_225), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g405 ( .A(n_226), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g315 ( .A(n_227), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g424 ( .A(n_227), .Y(n_424) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_228), .A2(n_236), .B(n_247), .Y(n_235) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_228), .A2(n_236), .B(n_247), .Y(n_288) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2x1_ASAP7_75t_SL g303 ( .A(n_229), .B(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g323 ( .A(n_230), .Y(n_323) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_248), .Y(n_232) );
AND2x2_ASAP7_75t_L g330 ( .A(n_233), .B(n_290), .Y(n_330) );
OR2x2_ASAP7_75t_L g497 ( .A(n_233), .B(n_328), .Y(n_497) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g310 ( .A(n_234), .B(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g342 ( .A(n_234), .Y(n_342) );
AND2x2_ASAP7_75t_L g469 ( .A(n_234), .B(n_249), .Y(n_469) );
AND2x4_ASAP7_75t_L g485 ( .A(n_234), .B(n_382), .Y(n_485) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_235), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_240), .B(n_242), .Y(n_237) );
INVx2_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
INVxp67_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
OR2x2_ASAP7_75t_L g346 ( .A(n_248), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g393 ( .A(n_248), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_265), .Y(n_248) );
AND2x4_ASAP7_75t_L g287 ( .A(n_249), .B(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_249), .Y(n_332) );
INVx1_ASAP7_75t_L g358 ( .A(n_249), .Y(n_358) );
AND2x2_ASAP7_75t_L g401 ( .A(n_249), .B(n_321), .Y(n_401) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_257), .B(n_264), .Y(n_250) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x4_ASAP7_75t_L g362 ( .A(n_265), .B(n_290), .Y(n_362) );
INVx1_ASAP7_75t_L g376 ( .A(n_265), .Y(n_376) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_266), .Y(n_306) );
INVx2_ASAP7_75t_L g329 ( .A(n_266), .Y(n_329) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_269), .B(n_279), .Y(n_267) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_269), .A2(n_279), .B(n_322), .Y(n_321) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B(n_278), .Y(n_274) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g443 ( .A(n_283), .B(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g464 ( .A(n_283), .Y(n_464) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_284), .B(n_453), .Y(n_467) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g374 ( .A(n_287), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g437 ( .A(n_287), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g462 ( .A(n_287), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g506 ( .A(n_287), .Y(n_506) );
AND2x2_ASAP7_75t_L g359 ( .A(n_288), .B(n_329), .Y(n_359) );
AND2x4_ASAP7_75t_L g361 ( .A(n_288), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g366 ( .A(n_288), .B(n_319), .Y(n_366) );
AND2x4_ASAP7_75t_L g381 ( .A(n_288), .B(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_306), .Y(n_289) );
INVx2_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
INVx2_ASAP7_75t_L g333 ( .A(n_290), .Y(n_333) );
BUFx2_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
INVx1_ASAP7_75t_L g403 ( .A(n_290), .Y(n_403) );
AND2x2_ASAP7_75t_L g463 ( .A(n_290), .B(n_321), .Y(n_463) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2x1_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OAI21x1_ASAP7_75t_SL g293 ( .A1(n_294), .A2(n_299), .B(n_303), .Y(n_293) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g343 ( .A(n_306), .B(n_311), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_317), .B(n_324), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_310), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g486 ( .A(n_310), .Y(n_486) );
AND2x2_ASAP7_75t_L g498 ( .A(n_310), .B(n_318), .Y(n_498) );
BUFx2_ASAP7_75t_L g438 ( .A(n_311), .Y(n_438) );
INVx1_ASAP7_75t_L g512 ( .A(n_311), .Y(n_512) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_315), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_318), .A2(n_509), .B1(n_511), .B2(n_513), .Y(n_508) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_SL g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OR2x6_ASAP7_75t_L g328 ( .A(n_320), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g382 ( .A(n_320), .Y(n_382) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_331), .B2(n_334), .Y(n_324) );
INVx2_ASAP7_75t_SL g369 ( .A(n_325), .Y(n_369) );
OR2x2_ASAP7_75t_L g398 ( .A(n_325), .B(n_337), .Y(n_398) );
INVx2_ASAP7_75t_L g435 ( .A(n_326), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g483 ( .A(n_328), .B(n_333), .Y(n_483) );
OR2x2_ASAP7_75t_L g516 ( .A(n_328), .B(n_342), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g404 ( .A(n_332), .B(n_359), .Y(n_404) );
INVx1_ASAP7_75t_L g380 ( .A(n_333), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_333), .B(n_357), .Y(n_420) );
OR2x2_ASAP7_75t_L g456 ( .A(n_333), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g453 ( .A(n_335), .Y(n_453) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g354 ( .A(n_336), .Y(n_354) );
INVx1_ASAP7_75t_L g406 ( .A(n_337), .Y(n_406) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_337), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_364), .Y(n_338) );
INVx2_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx2_ASAP7_75t_L g410 ( .A(n_342), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_342), .B(n_362), .Y(n_415) );
AND2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g488 ( .A(n_343), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_344), .Y(n_490) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g468 ( .A(n_347), .B(n_469), .Y(n_468) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_348), .B(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g481 ( .A(n_349), .Y(n_481) );
OR2x6_ASAP7_75t_L g349 ( .A(n_350), .B(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g444 ( .A(n_351), .Y(n_444) );
AND2x2_ASAP7_75t_L g504 ( .A(n_351), .B(n_354), .Y(n_504) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g385 ( .A(n_353), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_353), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_354), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g495 ( .A(n_354), .Y(n_495) );
NAND2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_360), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_357), .Y(n_458) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221x1_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_370), .B2(n_374), .C(n_377), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_400), .B1(n_404), .B2(n_405), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_367), .A2(n_408), .B1(n_411), .B2(n_414), .Y(n_407) );
INVxp67_ASAP7_75t_SL g505 ( .A(n_367), .Y(n_505) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g445 ( .A(n_372), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_375), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_375), .B(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_383), .B2(n_388), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AND2x4_ASAP7_75t_L g448 ( .A(n_380), .B(n_393), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_381), .A2(n_391), .B1(n_394), .B2(n_397), .Y(n_390) );
AND2x2_ASAP7_75t_L g471 ( .A(n_381), .B(n_438), .Y(n_471) );
OR2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g452 ( .A(n_385), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g473 ( .A(n_385), .Y(n_473) );
AND2x2_ASAP7_75t_L g494 ( .A(n_385), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g511 ( .A(n_385), .B(n_512), .Y(n_511) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_390), .B(n_399), .C(n_407), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_396), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_405), .A2(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g510 ( .A(n_413), .Y(n_510) );
INVx1_ASAP7_75t_L g426 ( .A(n_414), .Y(n_426) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_475), .Y(n_416) );
NAND3xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_432), .C(n_449), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g509 ( .A1(n_429), .A2(n_484), .B1(n_495), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g517 ( .A(n_429), .Y(n_517) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_439), .B(n_441), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_445), .B2(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_448), .A2(n_472), .B(n_492), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_458), .B(n_459), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_455), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g480 ( .A(n_457), .Y(n_480) );
NAND3xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_465), .C(n_470), .Y(n_459) );
NAND3xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_462), .C(n_464), .Y(n_460) );
AND2x2_ASAP7_75t_L g492 ( .A(n_463), .B(n_485), .Y(n_492) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .C(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_501), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_482), .B(n_489), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND4xp25_ASAP7_75t_SL g482 ( .A(n_483), .B(n_484), .C(n_486), .D(n_487), .Y(n_482) );
INVx3_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_491), .B(n_493), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B1(n_498), .B2(n_499), .Y(n_493) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_507), .Y(n_501) );
AOI21xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_505), .B(n_506), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_504), .A2(n_513), .B1(n_515), .B2(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OAI211xp5_ASAP7_75t_SL g518 ( .A1(n_519), .A2(n_528), .B(n_711), .C(n_739), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g718 ( .A(n_525), .Y(n_718) );
AND2x2_ASAP7_75t_L g737 ( .A(n_526), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_527), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g710 ( .A(n_529), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_529), .A2(n_710), .B1(n_740), .B2(n_755), .C(n_756), .Y(n_739) );
AND3x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_634), .C(n_674), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_586), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_541), .B1(n_566), .B2(n_570), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_533), .Y(n_532) );
AND2x6_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
OR2x6_ASAP7_75t_L g618 ( .A(n_534), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g568 ( .A(n_535), .Y(n_568) );
AND3x1_ASAP7_75t_L g591 ( .A(n_535), .B(n_592), .C(n_595), .Y(n_591) );
INVx2_ASAP7_75t_L g673 ( .A(n_535), .Y(n_673) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x4_ASAP7_75t_L g569 ( .A(n_537), .B(n_540), .Y(n_569) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_537), .Y(n_671) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g725 ( .A(n_538), .Y(n_725) );
INVx1_ASAP7_75t_L g641 ( .A(n_539), .Y(n_641) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g646 ( .A(n_540), .Y(n_646) );
OR2x2_ASAP7_75t_L g724 ( .A(n_540), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g730 ( .A(n_540), .B(n_725), .Y(n_730) );
OAI221xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_548), .B1(n_549), .B2(n_554), .C(n_555), .Y(n_541) );
INVx4_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g551 ( .A(n_546), .B(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g574 ( .A(n_546), .B(n_547), .Y(n_574) );
INVx1_ASAP7_75t_L g662 ( .A(n_547), .Y(n_662) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g585 ( .A(n_550), .Y(n_585) );
BUFx12f_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g657 ( .A(n_551), .Y(n_657) );
AND2x4_ASAP7_75t_L g564 ( .A(n_552), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g558 ( .A(n_553), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g583 ( .A(n_553), .B(n_565), .Y(n_583) );
BUFx4f_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g643 ( .A(n_558), .Y(n_643) );
INVx2_ASAP7_75t_L g648 ( .A(n_558), .Y(n_648) );
INVx2_ASAP7_75t_L g565 ( .A(n_559), .Y(n_565) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_562), .Y(n_577) );
BUFx6f_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g658 ( .A(n_563), .B(n_641), .Y(n_658) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g666 ( .A(n_565), .Y(n_666) );
CKINVDCx8_ASAP7_75t_R g566 ( .A(n_567), .Y(n_566) );
AND2x6_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B1(n_576), .B2(n_578), .C(n_579), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
CKINVDCx8_ASAP7_75t_R g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_578), .A2(n_679), .B1(n_683), .B2(n_684), .C1(n_686), .C2(n_687), .Y(n_678) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_596), .B1(n_618), .B2(n_621), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_588), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g677 ( .A(n_593), .Y(n_677) );
AND2x4_ASAP7_75t_L g684 ( .A(n_593), .B(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_SL g687 ( .A(n_593), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_603), .B1(n_604), .B2(n_609), .C(n_610), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_599), .Y(n_622) );
OR2x6_ASAP7_75t_L g676 ( .A(n_599), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_SL g695 ( .A(n_599), .B(n_692), .Y(n_695) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g607 ( .A(n_601), .Y(n_607) );
AND2x4_ASAP7_75t_L g616 ( .A(n_601), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g608 ( .A(n_602), .Y(n_608) );
INVx2_ASAP7_75t_L g617 ( .A(n_602), .Y(n_617) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx12f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_606), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x4_ASAP7_75t_L g682 ( .A(n_607), .B(n_608), .Y(n_682) );
BUFx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_612), .Y(n_629) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_613), .Y(n_699) );
INVx4_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx4_ASAP7_75t_L g703 ( .A(n_615), .Y(n_703) );
INVx5_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_616), .Y(n_633) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_617), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_624), .B2(n_627), .C(n_628), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_623), .A2(n_637), .B1(n_644), .B2(n_645), .Y(n_636) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI31xp33_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_658), .A3(n_659), .B(n_667), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_649), .Y(n_635) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
AND2x4_ASAP7_75t_L g652 ( .A(n_640), .B(n_653), .Y(n_652) );
AND2x6_ASAP7_75t_L g655 ( .A(n_640), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AND2x4_ASAP7_75t_L g661 ( .A(n_646), .B(n_662), .Y(n_661) );
AND2x4_ASAP7_75t_L g664 ( .A(n_646), .B(n_665), .Y(n_664) );
INVx5_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_654), .B2(n_655), .Y(n_649) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
CKINVDCx14_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g720 ( .A(n_662), .B(n_721), .C(n_723), .Y(n_720) );
AND2x4_ASAP7_75t_L g727 ( .A(n_662), .B(n_728), .Y(n_727) );
CKINVDCx8_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g708 ( .A(n_673), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_694), .B(n_704), .Y(n_674) );
AND2x2_ASAP7_75t_SL g698 ( .A(n_677), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g691 ( .A(n_682), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
CKINVDCx8_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_R g702 ( .A(n_692), .Y(n_702) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_701), .Y(n_696) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_731), .B1(n_732), .B2(n_734), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx4_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_717), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g738 ( .A(n_718), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_726), .Y(n_719) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_720), .Y(n_759) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx11_ASAP7_75t_R g762 ( .A(n_722), .Y(n_762) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g763 ( .A(n_726), .Y(n_763) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g755 ( .A(n_740), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_746), .B1(n_753), .B2(n_754), .Y(n_740) );
INVx1_ASAP7_75t_L g753 ( .A(n_741), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_742), .Y(n_745) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g754 ( .A(n_746), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_746) );
INVx1_ASAP7_75t_L g752 ( .A(n_747), .Y(n_752) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x6_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
endmodule