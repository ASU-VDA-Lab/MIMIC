module fake_jpeg_11737_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_83),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_72),
.Y(n_77)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_59),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_70),
.B1(n_57),
.B2(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_67),
.B1(n_5),
.B2(n_6),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_22),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_73),
.B1(n_67),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_60),
.B1(n_71),
.B2(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_95),
.B1(n_19),
.B2(n_48),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_56),
.B1(n_58),
.B2(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_68),
.B1(n_66),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_73),
.B1(n_67),
.B2(n_5),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_61),
.B1(n_54),
.B2(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_97),
.B(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_109),
.B1(n_111),
.B2(n_116),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_3),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_84),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_119),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_7),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_4),
.B(n_6),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_134),
.Y(n_145)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_92),
.B(n_36),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_92),
.B(n_8),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_136),
.B(n_9),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_34),
.C(n_47),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_17),
.C(n_46),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_49),
.B(n_45),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_7),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_8),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_144),
.C(n_146),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_153),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_9),
.C(n_10),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_151),
.C(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_120),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_152),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_10),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_128),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_125),
.B(n_124),
.Y(n_159)
);

AO221x1_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_128),
.B1(n_132),
.B2(n_150),
.C(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_130),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_128),
.B1(n_132),
.B2(n_144),
.C(n_147),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_148),
.A3(n_131),
.B1(n_145),
.B2(n_136),
.C1(n_12),
.C2(n_13),
.Y(n_166)
);

NAND2xp67_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_11),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_12),
.Y(n_168)
);


endmodule