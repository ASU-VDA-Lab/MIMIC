module fake_jpeg_2612_n_149 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_149);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_1),
.C(n_4),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_20),
.C(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_8),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_55),
.C(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_31),
.B(n_35),
.C(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_67),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_22),
.C(n_16),
.Y(n_55)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_33),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_16),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_19),
.C(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_4),
.Y(n_92)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_44),
.B(n_40),
.C(n_41),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_83),
.B1(n_93),
.B2(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_30),
.B1(n_34),
.B2(n_44),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_88),
.B1(n_94),
.B2(n_64),
.Y(n_103)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_92),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_19),
.B1(n_23),
.B2(n_48),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_8),
.C(n_10),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_103),
.B1(n_61),
.B2(n_63),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_57),
.B(n_66),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_86),
.B(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_106),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_79),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_79),
.A3(n_91),
.B1(n_77),
.B2(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AO221x1_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_121),
.B1(n_98),
.B2(n_96),
.C(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_111),
.B1(n_99),
.B2(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_104),
.C(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_124),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_122),
.B2(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_128),
.C(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_137),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_142),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_138),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_138),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_145),
.B(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_140),
.B1(n_120),
.B2(n_105),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_104),
.Y(n_149)
);


endmodule