module fake_jpeg_17348_n_356 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_47),
.Y(n_82)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_17),
.B(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_59),
.Y(n_74)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_57),
.Y(n_86)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_12),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_27),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_38),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_14),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_16),
.B1(n_29),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_72),
.A2(n_73),
.B1(n_103),
.B2(n_106),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_29),
.B1(n_25),
.B2(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_75),
.B(n_78),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_80),
.B(n_93),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_21),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_84),
.B(n_108),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_37),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_107),
.B(n_3),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_113),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_41),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_40),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_105)
);

OA22x2_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_20),
.B1(n_4),
.B2(n_7),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_37),
.B1(n_33),
.B2(n_15),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_60),
.B(n_12),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_122),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_50),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_111),
.A2(n_120),
.B(n_31),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_48),
.B(n_26),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_58),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_10),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_61),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_166),
.C(n_152),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_85),
.B1(n_115),
.B2(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_132),
.B1(n_152),
.B2(n_156),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_26),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_SL g176 ( 
.A(n_126),
.B(n_127),
.C(n_137),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_0),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_10),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_20),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_123),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_20),
.B(n_4),
.C(n_5),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_SL g198 ( 
.A(n_131),
.B(n_143),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_103),
.B1(n_105),
.B2(n_118),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_133),
.B(n_148),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_140),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_165),
.B1(n_170),
.B2(n_129),
.Y(n_178)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_149),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_8),
.B1(n_9),
.B2(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_92),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_74),
.B(n_81),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_73),
.A2(n_106),
.B1(n_96),
.B2(n_71),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_79),
.B(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_158),
.B(n_162),
.Y(n_197)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_97),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_89),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_71),
.B1(n_89),
.B2(n_117),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_90),
.A2(n_94),
.B(n_104),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_77),
.A2(n_90),
.B1(n_98),
.B2(n_95),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_98),
.B1(n_126),
.B2(n_128),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_187),
.B1(n_196),
.B2(n_207),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_179),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_178),
.A2(n_190),
.B1(n_193),
.B2(n_204),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_142),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_194),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_126),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_130),
.A2(n_133),
.B1(n_127),
.B2(n_134),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_188),
.B(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_146),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_130),
.B1(n_138),
.B2(n_134),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_167),
.B(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_127),
.A2(n_142),
.B1(n_144),
.B2(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_199),
.B(n_186),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_131),
.B(n_144),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_204),
.B(n_208),
.Y(n_231)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_202),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_166),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_151),
.A2(n_163),
.B1(n_139),
.B2(n_150),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_196),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_208),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_136),
.B1(n_145),
.B2(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_211),
.A2(n_216),
.B1(n_235),
.B2(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_145),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_222),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_215),
.B(n_236),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_178),
.B1(n_190),
.B2(n_198),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_174),
.C(n_187),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_240),
.C(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_194),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_204),
.B1(n_172),
.B2(n_176),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_239),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_226),
.A2(n_217),
.B1(n_213),
.B2(n_240),
.Y(n_268)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_238),
.Y(n_246)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_209),
.B(n_177),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_231),
.B(n_239),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_172),
.A2(n_176),
.B1(n_185),
.B2(n_179),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_181),
.B1(n_182),
.B2(n_184),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_197),
.B(n_180),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_197),
.B(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_171),
.C(n_181),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_173),
.B(n_171),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_241),
.B(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_210),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_250),
.B(n_251),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_228),
.B1(n_225),
.B2(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_268),
.B1(n_212),
.B2(n_234),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_256),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_219),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_223),
.B(n_230),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_258),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_269),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_216),
.B(n_211),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

NAND2x1p5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_213),
.C(n_224),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_272),
.C(n_256),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_241),
.B(n_233),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_254),
.Y(n_295)
);

AOI322xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_220),
.A3(n_234),
.B1(n_212),
.B2(n_232),
.C1(n_229),
.C2(n_227),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_269),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_279),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_252),
.B1(n_267),
.B2(n_263),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_282),
.B1(n_246),
.B2(n_266),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_260),
.B1(n_249),
.B2(n_268),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_286),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_247),
.A2(n_259),
.B1(n_257),
.B2(n_272),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_265),
.C(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_286),
.C(n_246),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_259),
.C(n_251),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_248),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_291),
.B(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_296),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_290),
.Y(n_307)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_311),
.C(n_314),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_250),
.B1(n_266),
.B2(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_245),
.B1(n_261),
.B2(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_303),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_277),
.B1(n_281),
.B2(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_277),
.B(n_280),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_306),
.A2(n_283),
.B(n_275),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_279),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_308),
.B(n_285),
.CI(n_273),
.CON(n_315),
.SN(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_295),
.C(n_290),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_305),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_285),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_296),
.B(n_307),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_319),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_299),
.C(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_300),
.C(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_323),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_305),
.B(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_308),
.C(n_304),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_298),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

NOR2x1_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_313),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_SL g342 ( 
.A(n_330),
.B(n_325),
.C(n_318),
.Y(n_342)
);

INVx11_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_335),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_313),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_333),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_322),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_316),
.B(n_324),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_315),
.B(n_318),
.Y(n_340)
);

NAND4xp25_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_316),
.C(n_315),
.D(n_328),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_339),
.B(n_342),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_340),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_325),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_343),
.B(n_345),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_334),
.B(n_333),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_344),
.A2(n_332),
.B1(n_337),
.B2(n_336),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_341),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_351),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_347),
.A2(n_348),
.B(n_349),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_351),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_348),
.B(n_353),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_329),
.Y(n_356)
);


endmodule