module fake_netlist_6_88_n_1408 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1408);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1408;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_1196;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_161),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_86),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_132),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_383),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_150),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_117),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_282),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_70),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_241),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_193),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_13),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_187),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_212),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_287),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_246),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_46),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_237),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_264),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_375),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_255),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_96),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_214),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_249),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_236),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_265),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_26),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_225),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_40),
.B(n_202),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_297),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_295),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_318),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_66),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_85),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_141),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_208),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_168),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_149),
.B(n_231),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_80),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_185),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_270),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_1),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_260),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_352),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_317),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_76),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_48),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_194),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_41),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_340),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_198),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_238),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_142),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_372),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_322),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_294),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_233),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_205),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_134),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_176),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_204),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_197),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_156),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_116),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_226),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_25),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_235),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_257),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_166),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_114),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_251),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_319),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_334),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_111),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_371),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_62),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_139),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_240),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_19),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_291),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_53),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_L g470 ( 
.A(n_20),
.B(n_224),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_347),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_324),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_342),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_3),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_118),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_64),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_368),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_313),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_54),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_91),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_147),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_363),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_278),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_210),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_195),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_250),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_90),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_85),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_84),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_23),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_221),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_259),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_74),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_56),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_72),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_154),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_273),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_338),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_41),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_6),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_57),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_46),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_65),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_314),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_234),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_62),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_175),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_196),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_339),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_135),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_125),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_345),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_276),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_7),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_305),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_65),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_74),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_113),
.B(n_106),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_106),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_323),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_335),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_243),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_81),
.B(n_370),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_81),
.B(n_290),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_124),
.Y(n_525)
);

BUFx2_ASAP7_75t_SL g526 ( 
.A(n_327),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_207),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_355),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_306),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_5),
.B(n_25),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_310),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_158),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_164),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_357),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_358),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_309),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_40),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_293),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_190),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_110),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_227),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_308),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_184),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_153),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_285),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_244),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_123),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_157),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_23),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_3),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_148),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_55),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_94),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_254),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_97),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_253),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_369),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_256),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_201),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_382),
.Y(n_560)
);

BUFx2_ASAP7_75t_SL g561 ( 
.A(n_312),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_232),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_298),
.B(n_266),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_517),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_517),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_517),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_393),
.B(n_0),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_0),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_517),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_454),
.A2(n_462),
.B1(n_549),
.B2(n_407),
.Y(n_572)
);

AOI22x1_ASAP7_75t_SL g573 ( 
.A1(n_396),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_489),
.B(n_444),
.Y(n_574)
);

OAI22x1_ASAP7_75t_R g575 ( 
.A1(n_418),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_397),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_415),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_386),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_501),
.Y(n_579)
);

BUFx8_ASAP7_75t_SL g580 ( 
.A(n_400),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_397),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_392),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_404),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_406),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_409),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_404),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_404),
.Y(n_588)
);

OA21x2_ASAP7_75t_L g589 ( 
.A1(n_423),
.A2(n_6),
.B(n_7),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_429),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_444),
.B(n_8),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_401),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_412),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_406),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_501),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_393),
.B(n_8),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_390),
.B(n_9),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_9),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_406),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_406),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_437),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_445),
.B(n_10),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_419),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_416),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_453),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_426),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_467),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_390),
.B(n_421),
.Y(n_611)
);

NOR2x1_ASAP7_75t_L g612 ( 
.A(n_398),
.B(n_112),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_445),
.B(n_423),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_434),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_452),
.B(n_11),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_404),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_453),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_435),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_464),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_385),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_398),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_537),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_402),
.Y(n_625)
);

BUFx8_ASAP7_75t_SL g626 ( 
.A(n_433),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_402),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_530),
.A2(n_476),
.B1(n_488),
.B2(n_487),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_495),
.Y(n_632)
);

INVx6_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_408),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_421),
.B(n_14),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_499),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_519),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_493),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_408),
.B(n_15),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_556),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_495),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_556),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_552),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_494),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_592),
.B(n_414),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_564),
.Y(n_650)
);

OR2x2_ASAP7_75t_SL g651 ( 
.A(n_592),
.B(n_574),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_607),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_574),
.A2(n_502),
.B1(n_506),
.B2(n_503),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_611),
.B(n_457),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_611),
.B(n_389),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_571),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_565),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_626),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_642),
.B(n_511),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_590),
.Y(n_661)
);

CKINVDCx8_ASAP7_75t_R g662 ( 
.A(n_569),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_625),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_625),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_568),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_576),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_586),
.B(n_470),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_622),
.B(n_555),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_576),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_621),
.B(n_510),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_581),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_604),
.B(n_514),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_581),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_581),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_591),
.B(n_518),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_595),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_600),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_600),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_600),
.Y(n_680)
);

CKINVDCx6p67_ASAP7_75t_R g681 ( 
.A(n_632),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_601),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_601),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_636),
.B(n_523),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_633),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_645),
.B(n_436),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_606),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_608),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_644),
.B(n_524),
.Y(n_692)
);

INVx8_ASAP7_75t_L g693 ( 
.A(n_595),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_633),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_654),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_670),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_649),
.A2(n_599),
.B1(n_635),
.B2(n_598),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_655),
.B(n_585),
.Y(n_698)
);

INVx8_ASAP7_75t_L g699 ( 
.A(n_649),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_649),
.A2(n_613),
.B1(n_589),
.B2(n_597),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_670),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_649),
.B(n_570),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_672),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_689),
.B(n_602),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_689),
.B(n_585),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_662),
.B(n_630),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_673),
.A2(n_613),
.B1(n_589),
.B2(n_597),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_666),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_652),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_671),
.B(n_603),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_651),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_666),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_673),
.B(n_635),
.C(n_598),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_651),
.B(n_640),
.Y(n_714)
);

NOR2xp67_ASAP7_75t_L g715 ( 
.A(n_688),
.B(n_617),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_660),
.B(n_630),
.C(n_572),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_690),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_694),
.B(n_653),
.Y(n_718)
);

OAI221xp5_ASAP7_75t_L g719 ( 
.A1(n_657),
.A2(n_570),
.B1(n_615),
.B2(n_646),
.C(n_609),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_572),
.C(n_647),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_SL g721 ( 
.A(n_681),
.B(n_441),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_669),
.B(n_615),
.C(n_628),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_661),
.B(n_634),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_672),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_663),
.B(n_634),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_691),
.B(n_595),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_691),
.B(n_619),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_672),
.B(n_619),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_664),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_692),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_668),
.B(n_634),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_678),
.B(n_569),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_682),
.B(n_608),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_657),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_685),
.B(n_687),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_676),
.B(n_643),
.Y(n_736)
);

OAI221xp5_ASAP7_75t_L g737 ( 
.A1(n_650),
.A2(n_646),
.B1(n_609),
.B2(n_641),
.C(n_582),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_682),
.B(n_643),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_656),
.B(n_579),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_656),
.B(n_578),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_686),
.B(n_466),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_648),
.B(n_579),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_648),
.B(n_596),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_659),
.A2(n_641),
.B1(n_478),
.B2(n_560),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_659),
.B(n_580),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_665),
.B(n_623),
.C(n_610),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_665),
.B(n_667),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_667),
.B(n_577),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_674),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_674),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_675),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_679),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_652),
.B(n_529),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_680),
.B(n_538),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_695),
.B(n_658),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_704),
.B(n_681),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_710),
.B(n_545),
.Y(n_757)
);

OAI321xp33_ASAP7_75t_L g758 ( 
.A1(n_713),
.A2(n_623),
.A3(n_610),
.B1(n_594),
.B2(n_614),
.C(n_605),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_711),
.A2(n_452),
.B(n_513),
.C(n_473),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_742),
.B(n_596),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_732),
.A2(n_693),
.B(n_677),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_714),
.B(n_405),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_743),
.B(n_618),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_707),
.A2(n_424),
.B1(n_563),
.B2(n_513),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_749),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_714),
.A2(n_593),
.B(n_624),
.C(n_620),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_697),
.A2(n_473),
.B(n_388),
.C(n_391),
.Y(n_767)
);

O2A1O1Ixp5_ASAP7_75t_L g768 ( 
.A1(n_734),
.A2(n_465),
.B(n_547),
.C(n_403),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_705),
.A2(n_707),
.B(n_747),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_706),
.B(n_540),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_700),
.B(n_413),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_700),
.B(n_734),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_728),
.A2(n_693),
.B(n_677),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_702),
.A2(n_559),
.B1(n_554),
.B2(n_394),
.Y(n_774)
);

O2A1O1Ixp5_ASAP7_75t_L g775 ( 
.A1(n_698),
.A2(n_584),
.B(n_587),
.C(n_583),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_739),
.B(n_627),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_722),
.A2(n_612),
.B(n_395),
.Y(n_777)
);

AOI21x1_ASAP7_75t_L g778 ( 
.A1(n_726),
.A2(n_684),
.B(n_683),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_723),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_749),
.B(n_683),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_702),
.A2(n_716),
.B1(n_720),
.B2(n_718),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_748),
.B(n_631),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_735),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_727),
.A2(n_693),
.B(n_677),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_703),
.B(n_387),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_751),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_754),
.A2(n_616),
.B(n_588),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_708),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_719),
.A2(n_637),
.B(n_639),
.C(n_629),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_696),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_702),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_712),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_730),
.B(n_417),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_746),
.A2(n_410),
.B(n_399),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_741),
.B(n_550),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_699),
.A2(n_420),
.B1(n_422),
.B2(n_411),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_701),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_750),
.B(n_425),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_733),
.A2(n_443),
.B(n_439),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_699),
.A2(n_428),
.B1(n_430),
.B2(n_427),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_724),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_744),
.B(n_431),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_737),
.B(n_553),
.Y(n_805)
);

NOR2x1_ASAP7_75t_L g806 ( 
.A(n_745),
.B(n_526),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_740),
.A2(n_449),
.B(n_447),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_752),
.B(n_456),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_729),
.B(n_721),
.Y(n_809)
);

NOR2x1_ASAP7_75t_R g810 ( 
.A(n_709),
.B(n_432),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_699),
.A2(n_460),
.B1(n_461),
.B2(n_458),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_740),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_731),
.B(n_736),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_725),
.B(n_438),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_725),
.B(n_472),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_715),
.A2(n_638),
.B(n_482),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_695),
.B(n_440),
.Y(n_818)
);

AND2x6_ASAP7_75t_L g819 ( 
.A(n_711),
.B(n_475),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_695),
.B(n_442),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_695),
.B(n_561),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_732),
.A2(n_484),
.B(n_483),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_695),
.B(n_446),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_707),
.B(n_486),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_732),
.A2(n_507),
.B(n_492),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_695),
.B(n_448),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_702),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_704),
.B(n_638),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_702),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_709),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_729),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_742),
.B(n_521),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_704),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_707),
.B(n_527),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_709),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_707),
.B(n_535),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_700),
.A2(n_548),
.B(n_546),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_695),
.B(n_450),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_749),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_732),
.A2(n_557),
.B(n_455),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_695),
.B(n_451),
.Y(n_841)
);

NOR2x1p5_ASAP7_75t_SL g842 ( 
.A(n_696),
.B(n_459),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_711),
.A2(n_468),
.B1(n_471),
.B2(n_463),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_704),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_749),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_749),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_481),
.C(n_477),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_695),
.A2(n_575),
.B(n_491),
.C(n_496),
.Y(n_848)
);

AOI21xp33_ASAP7_75t_L g849 ( 
.A1(n_695),
.A2(n_497),
.B(n_485),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_695),
.B(n_498),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_749),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_695),
.B(n_504),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_695),
.B(n_505),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_707),
.B(n_512),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_695),
.B(n_515),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_SL g856 ( 
.A1(n_772),
.A2(n_522),
.B(n_520),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_757),
.B(n_525),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_844),
.B(n_528),
.Y(n_858)
);

AOI21x1_ASAP7_75t_SL g859 ( 
.A1(n_824),
.A2(n_573),
.B(n_532),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_782),
.A2(n_533),
.B1(n_534),
.B2(n_531),
.Y(n_860)
);

OAI21xp33_ASAP7_75t_SL g861 ( 
.A1(n_834),
.A2(n_16),
.B(n_17),
.Y(n_861)
);

O2A1O1Ixp5_ASAP7_75t_L g862 ( 
.A1(n_764),
.A2(n_837),
.B(n_777),
.C(n_807),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_831),
.B(n_115),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_844),
.B(n_821),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_780),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_812),
.B(n_536),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_783),
.B(n_539),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_778),
.A2(n_542),
.B(n_541),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_769),
.A2(n_544),
.B(n_543),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_760),
.B(n_551),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_833),
.B(n_558),
.Y(n_871)
);

AO31x2_ASAP7_75t_L g872 ( 
.A1(n_767),
.A2(n_836),
.A3(n_759),
.B(n_774),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_831),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_R g874 ( 
.A(n_756),
.B(n_562),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_781),
.B(n_18),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_816),
.B(n_18),
.Y(n_876)
);

OA21x2_ASAP7_75t_L g877 ( 
.A1(n_768),
.A2(n_120),
.B(n_119),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_831),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_820),
.B(n_19),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_854),
.A2(n_122),
.B(n_121),
.Y(n_880)
);

OA21x2_ASAP7_75t_L g881 ( 
.A1(n_775),
.A2(n_127),
.B(n_126),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_845),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_761),
.A2(n_384),
.B(n_129),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_851),
.B(n_128),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_821),
.B(n_130),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_784),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_771),
.A2(n_773),
.B(n_785),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_826),
.B(n_20),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_770),
.B(n_850),
.Y(n_889)
);

AND2x6_ASAP7_75t_L g890 ( 
.A(n_813),
.B(n_131),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_837),
.A2(n_136),
.B(n_137),
.C(n_133),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_853),
.B(n_21),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_805),
.A2(n_24),
.B(n_21),
.C(n_22),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_762),
.A2(n_140),
.B(n_138),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_763),
.B(n_22),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_776),
.B(n_24),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_755),
.B(n_26),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_830),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_791),
.A2(n_803),
.B(n_799),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_832),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_777),
.A2(n_144),
.B(n_143),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_797),
.A2(n_27),
.B(n_28),
.Y(n_903)
);

AO21x2_ASAP7_75t_L g904 ( 
.A1(n_807),
.A2(n_146),
.B(n_145),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_796),
.A2(n_152),
.B(n_151),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_793),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_815),
.A2(n_159),
.B(n_155),
.Y(n_907)
);

OAI21x1_ASAP7_75t_SL g908 ( 
.A1(n_796),
.A2(n_162),
.B(n_160),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_792),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_779),
.A2(n_165),
.B1(n_167),
.B2(n_163),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_795),
.B(n_29),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_SL g912 ( 
.A1(n_786),
.A2(n_170),
.B(n_169),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_806),
.B(n_171),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_839),
.B(n_172),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_832),
.B(n_30),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_846),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_840),
.A2(n_174),
.B(n_173),
.Y(n_917)
);

OAI22x1_ASAP7_75t_L g918 ( 
.A1(n_827),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_918)
);

NOR2x1_ASAP7_75t_L g919 ( 
.A(n_818),
.B(n_823),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_788),
.A2(n_178),
.B(n_177),
.Y(n_920)
);

AO31x2_ASAP7_75t_L g921 ( 
.A1(n_822),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_829),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_838),
.B(n_34),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_814),
.A2(n_180),
.B(n_179),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_847),
.B(n_181),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_835),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_787),
.A2(n_183),
.B(n_182),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_819),
.B(n_35),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_849),
.B(n_186),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_800),
.A2(n_189),
.B(n_188),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_819),
.B(n_35),
.Y(n_931)
);

NAND2x1_ASAP7_75t_L g932 ( 
.A(n_819),
.B(n_808),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_841),
.A2(n_36),
.B(n_37),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_852),
.B(n_36),
.Y(n_934)
);

INVx3_ASAP7_75t_SL g935 ( 
.A(n_794),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_825),
.A2(n_192),
.B(n_191),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_855),
.B(n_37),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_802),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_819),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_804),
.A2(n_200),
.B(n_199),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_809),
.B(n_38),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_766),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_843),
.B(n_38),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_798),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_801),
.A2(n_206),
.B(n_203),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_790),
.B(n_39),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_811),
.A2(n_380),
.B(n_211),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_810),
.Y(n_948)
);

AO31x2_ASAP7_75t_L g949 ( 
.A1(n_842),
.A2(n_43),
.A3(n_39),
.B(n_42),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_817),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_758),
.A2(n_213),
.B(n_209),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_758),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_848),
.A2(n_216),
.B(n_215),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_769),
.A2(n_218),
.B(n_217),
.Y(n_954)
);

CKINVDCx8_ASAP7_75t_R g955 ( 
.A(n_830),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_830),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_769),
.A2(n_220),
.B(n_219),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_828),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_830),
.B(n_222),
.Y(n_959)
);

OAI22x1_ASAP7_75t_L g960 ( 
.A1(n_770),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_757),
.B(n_45),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_765),
.B(n_223),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_780),
.Y(n_963)
);

O2A1O1Ixp5_ASAP7_75t_L g964 ( 
.A1(n_764),
.A2(n_277),
.B(n_379),
.C(n_378),
.Y(n_964)
);

AOI21xp33_ASAP7_75t_L g965 ( 
.A1(n_757),
.A2(n_47),
.B(n_48),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_831),
.Y(n_966)
);

AND3x4_ASAP7_75t_L g967 ( 
.A(n_816),
.B(n_49),
.C(n_50),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_844),
.B(n_51),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_772),
.A2(n_281),
.B1(n_377),
.B2(n_376),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_828),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_844),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_831),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_769),
.A2(n_229),
.B(n_228),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_769),
.A2(n_239),
.B(n_230),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_778),
.A2(n_245),
.B(n_242),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_757),
.B(n_52),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_769),
.A2(n_248),
.B(n_247),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_831),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_L g979 ( 
.A1(n_757),
.A2(n_55),
.B(n_56),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_757),
.B(n_57),
.Y(n_980)
);

AND3x2_ASAP7_75t_L g981 ( 
.A(n_757),
.B(n_58),
.C(n_59),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_757),
.B(n_58),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_757),
.A2(n_288),
.B1(n_374),
.B2(n_373),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_769),
.A2(n_258),
.B(n_252),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_769),
.A2(n_262),
.B(n_261),
.Y(n_985)
);

AO31x2_ASAP7_75t_L g986 ( 
.A1(n_764),
.A2(n_59),
.A3(n_60),
.B(n_61),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_SL g987 ( 
.A(n_830),
.B(n_263),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_769),
.A2(n_268),
.B(n_267),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_831),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_757),
.B(n_60),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_757),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_991)
);

OAI21x1_ASAP7_75t_SL g992 ( 
.A1(n_837),
.A2(n_271),
.B(n_269),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_844),
.B(n_63),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_830),
.B(n_272),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_757),
.B(n_66),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_765),
.B(n_274),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_757),
.A2(n_299),
.B1(n_366),
.B2(n_365),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_765),
.B(n_275),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_757),
.A2(n_296),
.B1(n_364),
.B2(n_362),
.Y(n_999)
);

AO21x2_ASAP7_75t_L g1000 ( 
.A1(n_957),
.A2(n_292),
.B(n_360),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_901),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_966),
.B(n_279),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_906),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_898),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_899),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_971),
.B(n_67),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_909),
.Y(n_1007)
);

CKINVDCx11_ASAP7_75t_R g1008 ( 
.A(n_955),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_889),
.A2(n_961),
.B1(n_943),
.B2(n_937),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_934),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1010)
);

AND2x6_ASAP7_75t_L g1011 ( 
.A(n_939),
.B(n_280),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_878),
.Y(n_1012)
);

AOI22x1_ASAP7_75t_L g1013 ( 
.A1(n_973),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1013)
);

AO21x2_ASAP7_75t_L g1014 ( 
.A1(n_977),
.A2(n_300),
.B(n_359),
.Y(n_1014)
);

AO21x2_ASAP7_75t_L g1015 ( 
.A1(n_868),
.A2(n_289),
.B(n_356),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_886),
.B(n_71),
.Y(n_1016)
);

AO21x1_ASAP7_75t_L g1017 ( 
.A1(n_905),
.A2(n_888),
.B(n_879),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_865),
.Y(n_1018)
);

BUFx2_ASAP7_75t_SL g1019 ( 
.A(n_886),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_864),
.B(n_71),
.Y(n_1020)
);

OR2x6_ASAP7_75t_L g1021 ( 
.A(n_876),
.B(n_72),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_963),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_892),
.A2(n_302),
.B(n_354),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_870),
.B(n_73),
.Y(n_1024)
);

OA21x2_ASAP7_75t_L g1025 ( 
.A1(n_902),
.A2(n_301),
.B(n_353),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_878),
.Y(n_1026)
);

AO21x2_ASAP7_75t_L g1027 ( 
.A1(n_992),
.A2(n_286),
.B(n_349),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_956),
.Y(n_1028)
);

NAND2x1p5_ASAP7_75t_L g1029 ( 
.A(n_972),
.B(n_283),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_R g1030 ( 
.A(n_926),
.B(n_73),
.Y(n_1030)
);

CKINVDCx6p67_ASAP7_75t_R g1031 ( 
.A(n_935),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_882),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_972),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_920),
.A2(n_284),
.B(n_348),
.Y(n_1034)
);

OAI221xp5_ASAP7_75t_SL g1035 ( 
.A1(n_976),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.C(n_78),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_858),
.B(n_75),
.Y(n_1036)
);

INVx6_ASAP7_75t_L g1037 ( 
.A(n_972),
.Y(n_1037)
);

AO21x2_ASAP7_75t_L g1038 ( 
.A1(n_908),
.A2(n_367),
.B(n_346),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_897),
.B(n_77),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_980),
.B(n_78),
.C(n_79),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_884),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_866),
.B(n_79),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_916),
.B(n_344),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_968),
.B(n_80),
.Y(n_1044)
);

BUFx8_ASAP7_75t_SL g1045 ( 
.A(n_948),
.Y(n_1045)
);

OA21x2_ASAP7_75t_L g1046 ( 
.A1(n_964),
.A2(n_343),
.B(n_341),
.Y(n_1046)
);

BUFx2_ASAP7_75t_SL g1047 ( 
.A(n_873),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_962),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_874),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_SL g1050 ( 
.A1(n_951),
.A2(n_337),
.B(n_336),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_872),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_958),
.B(n_82),
.Y(n_1052)
);

OA21x2_ASAP7_75t_L g1053 ( 
.A1(n_891),
.A2(n_333),
.B(n_332),
.Y(n_1053)
);

AO21x2_ASAP7_75t_L g1054 ( 
.A1(n_917),
.A2(n_331),
.B(n_329),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_869),
.A2(n_328),
.B(n_326),
.Y(n_1055)
);

AO21x2_ASAP7_75t_L g1056 ( 
.A1(n_936),
.A2(n_325),
.B(n_321),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_978),
.B(n_320),
.Y(n_1057)
);

BUFx8_ASAP7_75t_L g1058 ( 
.A(n_922),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_989),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_883),
.A2(n_316),
.B(n_315),
.Y(n_1060)
);

CKINVDCx11_ASAP7_75t_R g1061 ( 
.A(n_938),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_982),
.A2(n_311),
.B1(n_307),
.B2(n_304),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_993),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_876),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_990),
.B(n_83),
.C(n_84),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_970),
.B(n_303),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_872),
.Y(n_1067)
);

BUFx2_ASAP7_75t_SL g1068 ( 
.A(n_959),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_962),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_995),
.A2(n_83),
.B(n_86),
.C(n_87),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_954),
.A2(n_87),
.B(n_88),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_996),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_932),
.A2(n_88),
.B(n_89),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_996),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_974),
.A2(n_89),
.B(n_90),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_923),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_984),
.A2(n_92),
.B(n_93),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_965),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_941),
.B(n_95),
.Y(n_1079)
);

AO21x2_ASAP7_75t_L g1080 ( 
.A1(n_985),
.A2(n_98),
.B(n_99),
.Y(n_1080)
);

OR2x6_ASAP7_75t_L g1081 ( 
.A(n_998),
.B(n_99),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_872),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_100),
.B(n_101),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_986),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_986),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_975),
.A2(n_102),
.B(n_103),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_890),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_947),
.A2(n_104),
.B(n_105),
.Y(n_1088)
);

NAND3xp33_ASAP7_75t_L g1089 ( 
.A(n_871),
.B(n_903),
.C(n_860),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_944),
.B(n_933),
.C(n_919),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_986),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_927),
.A2(n_104),
.B(n_105),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_875),
.A2(n_107),
.B(n_108),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_994),
.B(n_863),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_894),
.A2(n_107),
.B(n_108),
.Y(n_1095)
);

BUFx2_ASAP7_75t_R g1096 ( 
.A(n_928),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_867),
.B(n_109),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_857),
.B(n_896),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_880),
.A2(n_929),
.B(n_885),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_950),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_895),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_915),
.B(n_111),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_914),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_940),
.A2(n_953),
.B(n_911),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_931),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_946),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_952),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_925),
.A2(n_907),
.B(n_930),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_979),
.A2(n_890),
.B1(n_960),
.B2(n_967),
.Y(n_1109)
);

BUFx8_ASAP7_75t_SL g1110 ( 
.A(n_859),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_981),
.Y(n_1111)
);

INVxp67_ASAP7_75t_SL g1112 ( 
.A(n_987),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_856),
.B(n_991),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_913),
.B(n_893),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_969),
.A2(n_861),
.B(n_924),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_949),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_904),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_949),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_SL g1119 ( 
.A(n_910),
.B(n_881),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_999),
.B(n_997),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_983),
.B(n_877),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_877),
.Y(n_1122)
);

CKINVDCx16_ASAP7_75t_R g1123 ( 
.A(n_918),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_921),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_945),
.A2(n_912),
.B(n_921),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_966),
.B(n_900),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_898),
.Y(n_1127)
);

AO21x2_ASAP7_75t_L g1128 ( 
.A1(n_887),
.A2(n_973),
.B(n_957),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_862),
.A2(n_769),
.B(n_772),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_898),
.Y(n_1130)
);

CKINVDCx16_ASAP7_75t_R g1131 ( 
.A(n_898),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_961),
.A2(n_764),
.A3(n_767),
.B(n_759),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_862),
.A2(n_973),
.B(n_957),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_971),
.B(n_757),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1032),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1009),
.A2(n_1107),
.B1(n_1109),
.B2(n_1022),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1074),
.B(n_1072),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1019),
.B(n_1069),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1001),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1129),
.A2(n_1118),
.B(n_1116),
.Y(n_1140)
);

CKINVDCx8_ASAP7_75t_R g1141 ( 
.A(n_1131),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1018),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1058),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1028),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1018),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1003),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1078),
.A2(n_1039),
.B1(n_1093),
.B2(n_1013),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1107),
.B(n_1098),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1007),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1058),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1026),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1013),
.A2(n_1010),
.B1(n_1089),
.B2(n_1042),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1041),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1100),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_1017),
.A2(n_1128),
.B(n_1118),
.Y(n_1155)
);

OAI221xp5_ASAP7_75t_L g1156 ( 
.A1(n_1035),
.A2(n_1076),
.B1(n_1020),
.B2(n_1077),
.C(n_1134),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_SL g1157 ( 
.A(n_1049),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1059),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1106),
.Y(n_1159)
);

AOI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1108),
.A2(n_1005),
.B(n_1099),
.Y(n_1160)
);

OAI221xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1021),
.A2(n_1070),
.B1(n_1081),
.B2(n_1016),
.C(n_1065),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1090),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1101),
.B(n_1041),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1040),
.A2(n_1120),
.B1(n_1114),
.B2(n_1095),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1008),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1048),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1051),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1051),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1048),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1067),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1026),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_1123),
.A2(n_1021),
.B1(n_1081),
.B2(n_1112),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1026),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1084),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1063),
.Y(n_1176)
);

AO21x1_ASAP7_75t_L g1177 ( 
.A1(n_1115),
.A2(n_1113),
.B(n_1114),
.Y(n_1177)
);

INVxp33_ASAP7_75t_L g1178 ( 
.A(n_1036),
.Y(n_1178)
);

BUFx2_ASAP7_75t_SL g1179 ( 
.A(n_1004),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1023),
.A2(n_1079),
.B1(n_1097),
.B2(n_1024),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1044),
.B(n_1033),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1091),
.Y(n_1183)
);

OAI222xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1111),
.A2(n_1030),
.B1(n_1123),
.B2(n_1016),
.C1(n_1096),
.C2(n_1061),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_1127),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1006),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1091),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1102),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1133),
.A2(n_1075),
.B(n_1071),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1002),
.Y(n_1190)
);

INVx8_ASAP7_75t_L g1191 ( 
.A(n_1011),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1037),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1124),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1066),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1031),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1126),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1133),
.A2(n_1000),
.B1(n_1025),
.B2(n_1034),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1037),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1103),
.B(n_1047),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1119),
.A2(n_1125),
.B(n_1000),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1064),
.B(n_1087),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1130),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1052),
.B(n_1105),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1083),
.Y(n_1204)
);

AO21x1_ASAP7_75t_SL g1205 ( 
.A1(n_1110),
.A2(n_1050),
.B(n_1094),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1012),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1012),
.B(n_1068),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1080),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1057),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1011),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1011),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_1011),
.Y(n_1213)
);

AOI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1104),
.A2(n_1025),
.B(n_1046),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1132),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1043),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1086),
.Y(n_1217)
);

BUFx4f_ASAP7_75t_SL g1218 ( 
.A(n_1131),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1132),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1132),
.B(n_1014),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1029),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1094),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1073),
.Y(n_1223)
);

BUFx4f_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1034),
.A2(n_1054),
.B(n_1056),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1142),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1156),
.A2(n_1147),
.B1(n_1152),
.B2(n_1136),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1203),
.B(n_1038),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1192),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1186),
.B(n_1027),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1145),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1148),
.B(n_1062),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1165),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1213),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1178),
.B(n_1092),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1135),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1148),
.B(n_1117),
.Y(n_1237)
);

CKINVDCx6p67_ASAP7_75t_R g1238 ( 
.A(n_1150),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1156),
.A2(n_1117),
.B1(n_1121),
.B2(n_1088),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1207),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1136),
.B(n_1055),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1193),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1188),
.B(n_1015),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1163),
.B(n_1060),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1211),
.Y(n_1245)
);

INVx4_ASAP7_75t_R g1246 ( 
.A(n_1157),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1167),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1182),
.B(n_1053),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1159),
.B(n_1122),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1140),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1168),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1149),
.Y(n_1252)
);

BUFx2_ASAP7_75t_L g1253 ( 
.A(n_1173),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1170),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1151),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1161),
.B(n_1194),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1139),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1176),
.B(n_1137),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1181),
.B(n_1137),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1154),
.B(n_1146),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1173),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1192),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1172),
.B(n_1196),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1192),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1152),
.A2(n_1177),
.B1(n_1164),
.B2(n_1162),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1190),
.B(n_1164),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1189),
.A2(n_1214),
.B(n_1204),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1222),
.B(n_1216),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1153),
.B(n_1166),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1215),
.A2(n_1219),
.B1(n_1191),
.B2(n_1205),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1221),
.A2(n_1218),
.B1(n_1195),
.B2(n_1201),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1161),
.B(n_1169),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1198),
.B(n_1169),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1157),
.A2(n_1213),
.B1(n_1199),
.B2(n_1138),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1171),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1158),
.Y(n_1276)
);

OAI221xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1184),
.A2(n_1197),
.B1(n_1223),
.B2(n_1138),
.C(n_1199),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1174),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1175),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1191),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1227),
.A2(n_1141),
.B1(n_1138),
.B2(n_1218),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1234),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1259),
.B(n_1180),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1256),
.B(n_1210),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1258),
.Y(n_1285)
);

NOR2x1_ASAP7_75t_L g1286 ( 
.A(n_1274),
.B(n_1144),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1256),
.B(n_1187),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1252),
.B(n_1183),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1247),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1247),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1250),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1251),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1235),
.B(n_1155),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1251),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1254),
.Y(n_1295)
);

OAI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1227),
.A2(n_1201),
.B1(n_1143),
.B2(n_1179),
.C(n_1202),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1265),
.A2(n_1271),
.B(n_1239),
.Y(n_1297)
);

OAI21xp33_ASAP7_75t_L g1298 ( 
.A1(n_1265),
.A2(n_1208),
.B(n_1220),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1233),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1228),
.B(n_1224),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1226),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1280),
.B(n_1212),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1269),
.B(n_1209),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1231),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1278),
.B(n_1224),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1232),
.A2(n_1191),
.B1(n_1212),
.B2(n_1225),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1260),
.B(n_1240),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1240),
.B(n_1237),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1236),
.B(n_1200),
.Y(n_1309)
);

NOR2xp67_ASAP7_75t_SL g1310 ( 
.A(n_1233),
.B(n_1212),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1268),
.B(n_1249),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1277),
.A2(n_1195),
.B1(n_1165),
.B2(n_1206),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1230),
.B(n_1200),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1272),
.A2(n_1197),
.B1(n_1184),
.B2(n_1217),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1279),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1244),
.B(n_1225),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1263),
.B(n_1160),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1289),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1290),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1311),
.B(n_1242),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1292),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1293),
.B(n_1243),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1293),
.B(n_1267),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1294),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1313),
.B(n_1267),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1313),
.B(n_1248),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1295),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1308),
.B(n_1257),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1305),
.B(n_1309),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1316),
.B(n_1317),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1297),
.B(n_1266),
.C(n_1241),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1285),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1307),
.B(n_1261),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1301),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1300),
.B(n_1279),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1304),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1282),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1283),
.B(n_1253),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1338),
.B(n_1300),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1334),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1330),
.B(n_1309),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1329),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1329),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1320),
.B(n_1305),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1336),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1321),
.Y(n_1346)
);

NAND2x1_ASAP7_75t_L g1347 ( 
.A(n_1337),
.B(n_1315),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1323),
.B(n_1291),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1331),
.A2(n_1296),
.B1(n_1284),
.B2(n_1281),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1318),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1337),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1319),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1322),
.B(n_1304),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1324),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1327),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1344),
.B(n_1323),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1342),
.B(n_1329),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1340),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1343),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1348),
.Y(n_1360)
);

OAI311xp33_ASAP7_75t_L g1361 ( 
.A1(n_1346),
.A2(n_1298),
.A3(n_1287),
.B1(n_1306),
.C1(n_1270),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1345),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1345),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1350),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1349),
.B(n_1286),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1347),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1341),
.B(n_1326),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1341),
.B(n_1325),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1357),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1356),
.B(n_1353),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1365),
.B(n_1364),
.C(n_1314),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1358),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1367),
.B(n_1299),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1359),
.A2(n_1312),
.B1(n_1310),
.B2(n_1302),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1357),
.A2(n_1302),
.B1(n_1332),
.B2(n_1335),
.Y(n_1375)
);

NAND4xp25_ASAP7_75t_L g1376 ( 
.A(n_1360),
.B(n_1333),
.C(n_1303),
.D(n_1288),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1373),
.B(n_1299),
.Y(n_1377)
);

OA22x2_ASAP7_75t_L g1378 ( 
.A1(n_1374),
.A2(n_1375),
.B1(n_1369),
.B2(n_1360),
.Y(n_1378)
);

OAI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1371),
.A2(n_1339),
.B1(n_1366),
.B2(n_1354),
.C(n_1355),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1376),
.B(n_1185),
.Y(n_1380)
);

NOR3xp33_ASAP7_75t_L g1381 ( 
.A(n_1372),
.B(n_1366),
.C(n_1328),
.Y(n_1381)
);

OAI211xp5_ASAP7_75t_L g1382 ( 
.A1(n_1379),
.A2(n_1380),
.B(n_1381),
.C(n_1378),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1377),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1381),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1381),
.B(n_1370),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_1380),
.B(n_1276),
.C(n_1229),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1381),
.B(n_1306),
.C(n_1352),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_L g1388 ( 
.A(n_1382),
.B(n_1229),
.C(n_1245),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1384),
.B(n_1362),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1383),
.B(n_1367),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1390),
.Y(n_1391)
);

NAND4xp75_ASAP7_75t_L g1392 ( 
.A(n_1389),
.B(n_1385),
.C(n_1185),
.D(n_1246),
.Y(n_1392)
);

INVxp33_ASAP7_75t_L g1393 ( 
.A(n_1392),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1393),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1394),
.A2(n_1388),
.B(n_1391),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1394),
.A2(n_1386),
.B1(n_1387),
.B2(n_1238),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1395),
.B(n_1362),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1396),
.Y(n_1398)
);

OAI211xp5_ASAP7_75t_L g1399 ( 
.A1(n_1398),
.A2(n_1238),
.B(n_1262),
.C(n_1264),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1397),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1400),
.A2(n_1351),
.B1(n_1264),
.B2(n_1262),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1399),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1402),
.A2(n_1351),
.B1(n_1368),
.B2(n_1229),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1401),
.A2(n_1368),
.B1(n_1363),
.B2(n_1270),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1403),
.A2(n_1273),
.B(n_1361),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1404),
.A2(n_1280),
.B(n_1255),
.Y(n_1406)
);

OR2x6_ASAP7_75t_L g1407 ( 
.A(n_1406),
.B(n_1275),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1407),
.A2(n_1405),
.B1(n_1275),
.B2(n_1255),
.Y(n_1408)
);


endmodule