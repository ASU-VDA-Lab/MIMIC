module fake_jpeg_28671_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_47),
.Y(n_93)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g96 ( 
.A(n_50),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_15),
.C(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_55),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g103 ( 
.A(n_52),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_15),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_56),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_70),
.Y(n_95)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_21),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_64),
.Y(n_112)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_0),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_18),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_24),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_83),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_85),
.Y(n_122)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_87),
.B(n_113),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_28),
.B1(n_42),
.B2(n_33),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_90),
.A2(n_94),
.B1(n_105),
.B2(n_118),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_28),
.B1(n_20),
.B2(n_43),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_92),
.A2(n_99),
.B1(n_109),
.B2(n_130),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_36),
.B1(n_20),
.B2(n_43),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_30),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_98),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_32),
.B(n_70),
.C(n_41),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_100),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_18),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_125),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_43),
.B1(n_30),
.B2(n_40),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_65),
.A2(n_30),
.B1(n_43),
.B2(n_40),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_44),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_52),
.B(n_29),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_104),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_63),
.A2(n_40),
.B1(n_29),
.B2(n_26),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_82),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_146),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_49),
.B(n_3),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_136),
.A2(n_165),
.B(n_5),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

BUFx2_ASAP7_75t_SL g143 ( 
.A(n_103),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_25),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_149),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_25),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_39),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_151),
.B(n_168),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_39),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_39),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_161),
.Y(n_197)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_74),
.B1(n_31),
.B2(n_52),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_160),
.A2(n_112),
.B1(n_115),
.B2(n_93),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_74),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_163),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_31),
.B1(n_50),
.B2(n_4),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_167),
.Y(n_209)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_170),
.Y(n_181)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_177),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_172),
.A2(n_123),
.B1(n_131),
.B2(n_120),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_2),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_178),
.Y(n_195)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_89),
.B(n_3),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_50),
.B1(n_4),
.B2(n_5),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_93),
.B1(n_120),
.B2(n_117),
.Y(n_208)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_98),
.B(n_3),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_108),
.C(n_127),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_110),
.B1(n_111),
.B2(n_86),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_202),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_98),
.B1(n_111),
.B2(n_86),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_122),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_184),
.B(n_139),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_115),
.B(n_112),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_200),
.B(n_210),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_92),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_177),
.C(n_157),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_213),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_131),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_117),
.B1(n_131),
.B2(n_108),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_208),
.A2(n_159),
.B1(n_170),
.B2(n_140),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_123),
.B1(n_6),
.B2(n_7),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_173),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_138),
.B(n_7),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_7),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_142),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_156),
.B1(n_167),
.B2(n_154),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_240),
.C(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_228),
.B1(n_232),
.B2(n_252),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_141),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_226),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_180),
.B1(n_179),
.B2(n_158),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_134),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_237),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_163),
.B1(n_153),
.B2(n_145),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_234),
.A2(n_196),
.B(n_198),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_236),
.B(n_241),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_171),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_210),
.A2(n_195),
.B(n_189),
.Y(n_239)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_239),
.A2(n_216),
.B(n_194),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_135),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_247),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_246),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_137),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_258),
.B1(n_186),
.B2(n_205),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_166),
.C(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_218),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_12),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_251),
.B(n_254),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_164),
.B1(n_12),
.B2(n_13),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_218),
.Y(n_253)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_253),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_12),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_202),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_255),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_208),
.A2(n_13),
.B1(n_184),
.B2(n_221),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_194),
.B1(n_205),
.B2(n_193),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_186),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_257),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_190),
.B1(n_220),
.B2(n_199),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_262),
.B(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_185),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_185),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_281),
.C(n_240),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_267),
.A2(n_268),
.B1(n_273),
.B2(n_276),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_255),
.A2(n_193),
.B1(n_219),
.B2(n_198),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_216),
.C(n_222),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_284),
.B(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_219),
.B1(n_222),
.B2(n_203),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_244),
.A2(n_219),
.B1(n_196),
.B2(n_194),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_234),
.B(n_254),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_203),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_245),
.A2(n_211),
.B(n_216),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_204),
.B1(n_211),
.B2(n_229),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_288),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_231),
.B(n_204),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_245),
.B1(n_232),
.B2(n_228),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_290),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_245),
.A2(n_236),
.B(n_257),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_294),
.B(n_307),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_235),
.B(n_239),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_296),
.B(n_300),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_245),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_313),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_225),
.Y(n_299)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_262),
.A2(n_252),
.B1(n_246),
.B2(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_265),
.B(n_227),
.Y(n_301)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_265),
.B(n_249),
.Y(n_306)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_278),
.A2(n_234),
.B(n_237),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_243),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_310),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_240),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_306),
.Y(n_327)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_250),
.B1(n_238),
.B2(n_242),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_319),
.B1(n_320),
.B2(n_283),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_270),
.B(n_249),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_315),
.Y(n_344)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_316),
.B(n_288),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_274),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_261),
.C(n_266),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_324),
.B(n_327),
.C(n_330),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_281),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_301),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_293),
.A2(n_291),
.B1(n_276),
.B2(n_287),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_338),
.B1(n_339),
.B2(n_304),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_292),
.C(n_290),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_299),
.B(n_233),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_279),
.C(n_294),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_284),
.C(n_269),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_336),
.C(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_264),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_297),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_289),
.B1(n_269),
.B2(n_260),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_263),
.B1(n_224),
.B2(n_272),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_296),
.B(n_258),
.C(n_233),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_341),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_302),
.B1(n_263),
.B2(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_349),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_335),
.B1(n_337),
.B2(n_342),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_350),
.B(n_357),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_322),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_317),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_354),
.Y(n_365)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_327),
.B(n_313),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_361),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_305),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_362),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_333),
.A2(n_296),
.B1(n_311),
.B2(n_305),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_360),
.A2(n_339),
.B1(n_332),
.B2(n_328),
.Y(n_373)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_332),
.B(n_296),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_308),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_364),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_324),
.C(n_330),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_379),
.C(n_357),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_370),
.A2(n_360),
.B1(n_350),
.B2(n_320),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_340),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_374),
.B(n_351),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_347),
.A2(n_304),
.B1(n_344),
.B2(n_334),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_375),
.B(n_346),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_352),
.A2(n_345),
.B(n_362),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_377),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_326),
.C(n_307),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_381),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_355),
.B1(n_267),
.B2(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

NOR3xp33_ASAP7_75t_SL g385 ( 
.A(n_369),
.B(n_279),
.C(n_303),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_370),
.B1(n_285),
.B2(n_273),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_387),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_315),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_389),
.B(n_390),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_374),
.B(n_359),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_368),
.B(n_251),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_382),
.A2(n_377),
.B(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_379),
.C(n_366),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_401),
.C(n_391),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_384),
.A2(n_367),
.B(n_378),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_397),
.A2(n_388),
.B(n_385),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_380),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_373),
.C(n_375),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_404),
.Y(n_413)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_403),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_392),
.B(n_387),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_407),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_310),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_398),
.A2(n_401),
.B1(n_399),
.B2(n_395),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_409),
.B(n_268),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_397),
.A2(n_371),
.B1(n_318),
.B2(n_319),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_396),
.C(n_405),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_410),
.B(n_412),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_403),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_415),
.B(n_417),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_407),
.C(n_371),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_414),
.Y(n_419)
);

AOI33xp33_ASAP7_75t_L g420 ( 
.A1(n_419),
.A2(n_248),
.A3(n_253),
.B1(n_280),
.B2(n_411),
.B3(n_418),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_280),
.Y(n_421)
);


endmodule