module fake_jpeg_12096_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_14),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_46),
.B(n_58),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_29),
.B1(n_39),
.B2(n_38),
.Y(n_86)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_64),
.Y(n_89)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_59),
.Y(n_97)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_4),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_21),
.B(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_32),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_65),
.B1(n_71),
.B2(n_56),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_13),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_33),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_5),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_80),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_10),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_69),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_37),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_12),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_11),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_84),
.A2(n_86),
.B1(n_45),
.B2(n_107),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_35),
.B1(n_41),
.B2(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_91),
.A2(n_93),
.B1(n_109),
.B2(n_111),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_41),
.B1(n_35),
.B2(n_31),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_39),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_70),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_45),
.B(n_77),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_117),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_25),
.B(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_118),
.Y(n_124)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_113),
.B1(n_102),
.B2(n_81),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_60),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_43),
.B(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_61),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_130),
.C(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_127),
.B(n_128),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_73),
.Y(n_128)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_79),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_145),
.B(n_130),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_98),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_84),
.A2(n_93),
.B1(n_91),
.B2(n_96),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_88),
.B1(n_103),
.B2(n_92),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_82),
.B1(n_100),
.B2(n_83),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_106),
.B1(n_81),
.B2(n_90),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_156),
.B(n_157),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_90),
.B1(n_106),
.B2(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_98),
.B(n_89),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_98),
.B(n_89),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_170),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_123),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_130),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_137),
.B1(n_124),
.B2(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_182),
.C(n_155),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_123),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_184),
.A2(n_196),
.B(n_178),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_143),
.B1(n_124),
.B2(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_186),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_133),
.B1(n_126),
.B2(n_134),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.C(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_156),
.B1(n_142),
.B2(n_134),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_136),
.B1(n_158),
.B2(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_201),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_213),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_162),
.C(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_161),
.C(n_175),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_184),
.A2(n_190),
.B(n_167),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

AOI221xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_161),
.B1(n_172),
.B2(n_163),
.C(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_220),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_207),
.B(n_211),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_205),
.A2(n_186),
.B1(n_196),
.B2(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_209),
.Y(n_220)
);

BUFx12f_ASAP7_75t_SL g221 ( 
.A(n_212),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_175),
.C(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_173),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_167),
.B1(n_172),
.B2(n_191),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_182),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_204),
.B(n_208),
.C(n_211),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_225),
.A2(n_227),
.B(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_216),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_235),
.B(n_226),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_223),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_216),
.B(n_222),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_218),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.C(n_240),
.Y(n_243)
);

OAI31xp33_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_221),
.A3(n_224),
.B(n_223),
.Y(n_238)
);

AOI311xp33_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_239),
.A3(n_234),
.B(n_177),
.C(n_209),
.Y(n_241)
);

OAI321xp33_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_210),
.A3(n_174),
.B1(n_171),
.B2(n_147),
.C(n_169),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_214),
.A3(n_202),
.B1(n_210),
.B2(n_197),
.C1(n_159),
.C2(n_187),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_242),
.B(n_214),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.B(n_171),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_243),
.Y(n_247)
);


endmodule