module fake_jpeg_22013_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_17),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_43),
.Y(n_44)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_19),
.B1(n_21),
.B2(n_32),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_49),
.B1(n_55),
.B2(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_42),
.B1(n_23),
.B2(n_17),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_73),
.B1(n_51),
.B2(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_80),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_72),
.B1(n_36),
.B2(n_44),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_23),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_36),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_67),
.B1(n_73),
.B2(n_69),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_0),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_62),
.B1(n_52),
.B2(n_58),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_13),
.C(n_15),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_98),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_94),
.B(n_97),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_52),
.B1(n_35),
.B2(n_39),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_1),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_23),
.B1(n_37),
.B2(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_102),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_101),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_119),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_69),
.C(n_76),
.Y(n_108)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_114),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_69),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_84),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_72),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_70),
.Y(n_120)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_82),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_127),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_98),
.B(n_100),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_135),
.B(n_139),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_96),
.C(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_113),
.B(n_112),
.C(n_103),
.D(n_105),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_92),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_18),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_78),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_18),
.B(n_30),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_110),
.B1(n_105),
.B2(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_110),
.C(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_129),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_135),
.Y(n_156)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_159),
.B(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_151),
.C(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_164),
.C(n_30),
.Y(n_176)
);

AO221x1_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_79),
.B1(n_45),
.B2(n_34),
.C(n_4),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_129),
.B(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_135),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_30),
.B(n_18),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_133),
.C(n_139),
.Y(n_164)
);

XOR2x1_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_111),
.B1(n_79),
.B2(n_12),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_111),
.B1(n_145),
.B2(n_79),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_154),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_162),
.B1(n_167),
.B2(n_18),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_172),
.B(n_1),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_2),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_159),
.C(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_30),
.C(n_18),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_164),
.C(n_161),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_163),
.B1(n_160),
.B2(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_183),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_167),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_184),
.A2(n_170),
.A3(n_171),
.B1(n_175),
.B2(n_173),
.C1(n_11),
.C2(n_7),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_3),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_4),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_4),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_194),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_179),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_195),
.B(n_186),
.C(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_184),
.C(n_182),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_198),
.A2(n_5),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_197),
.C2(n_165),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_5),
.B(n_6),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_8),
.C(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_9),
.Y(n_203)
);


endmodule