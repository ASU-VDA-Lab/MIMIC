module fake_netlist_5_2172_n_1984 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_1984);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1984;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_69),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_177),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_29),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_99),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_137),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_36),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_97),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_48),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_101),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_53),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_0),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_22),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_53),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_91),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_94),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_145),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_110),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_17),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_25),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_60),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_78),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_49),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_148),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_168),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_109),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_131),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_39),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_112),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_12),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_28),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_180),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_93),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_15),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_66),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_65),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_165),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_96),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_8),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_140),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_31),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_82),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_167),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_198),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_81),
.Y(n_287)
);

BUFx8_ASAP7_75t_SL g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_57),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_103),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_13),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_74),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_169),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_121),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_133),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_58),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_79),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_76),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_179),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_150),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_8),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_138),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_50),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_120),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_1),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_21),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_28),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_1),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_18),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_39),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_172),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_44),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_51),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_71),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_68),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_46),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_26),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_161),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_139),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_31),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_61),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_84),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_126),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_19),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_186),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_182),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_155),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_36),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_108),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_152),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_14),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_158),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_196),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_54),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_142),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_183),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_75),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_189),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_30),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_62),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_95),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_49),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_55),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_115),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_50),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_20),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_16),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_176),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_190),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_85),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_123),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_149),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_6),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_153),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_45),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_188),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_162),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_11),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_197),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_24),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_72),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_102),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_89),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_117),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_64),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_63),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_144),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_125),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_200),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_15),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_194),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_23),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_42),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_65),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_111),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_136),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_86),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_83),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_98),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_37),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_43),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_20),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_41),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_156),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_129),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_127),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_118),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_88),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_40),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_77),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_55),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_10),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_21),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_130),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_61),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_184),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_288),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_305),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_219),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_294),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_312),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_273),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_294),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_318),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_255),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_359),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_250),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_250),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_271),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_329),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_205),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_259),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_226),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_250),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_262),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_240),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_269),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_282),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_274),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_269),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_331),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_279),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_270),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_269),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_281),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_292),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_275),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_278),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_269),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_283),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_269),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_286),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_286),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_219),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_296),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_284),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_285),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_289),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_286),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_392),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_210),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_286),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_263),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_299),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_286),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_300),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_353),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_303),
.Y(n_462)
);

BUFx2_ASAP7_75t_SL g463 ( 
.A(n_227),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_301),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_302),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_254),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_350),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_352),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_392),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_353),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_212),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_216),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_297),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_355),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_222),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_401),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_306),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_356),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_225),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_247),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_260),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_357),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_335),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_221),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_358),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_394),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_361),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_362),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_363),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_290),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_327),
.B(n_0),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_221),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_370),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_210),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_316),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_321),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_229),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_333),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_229),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_231),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_231),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_366),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_242),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_343),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_242),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_327),
.B(n_2),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_249),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_233),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_365),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_384),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_233),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_419),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_426),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_437),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_258),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_468),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_409),
.B(n_228),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_R g523 ( 
.A(n_441),
.B(n_372),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_496),
.B(n_258),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_430),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_433),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_266),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_266),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_442),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_412),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_444),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_368),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_445),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_417),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_418),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_410),
.B(n_368),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_418),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_450),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_451),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_447),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_452),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_453),
.Y(n_548)
);

AND2x6_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_364),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_458),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_464),
.Y(n_554)
);

NOR2x1_ASAP7_75t_L g555 ( 
.A(n_462),
.B(n_364),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_473),
.B(n_364),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

AND2x6_ASAP7_75t_L g561 ( 
.A(n_495),
.B(n_235),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_479),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_481),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_485),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_487),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_494),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_422),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_489),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_423),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_410),
.B(n_287),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_499),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_500),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_425),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_448),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_448),
.B(n_287),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_411),
.B(n_235),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_414),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_491),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_413),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_416),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_431),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_435),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_435),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_480),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_463),
.B(n_393),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_492),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_424),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_421),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_424),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_427),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_415),
.B(n_393),
.Y(n_598)
);

INVx6_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_506),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_415),
.B(n_457),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_599),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_522),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_523),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_427),
.Y(n_606)
);

AO22x2_ASAP7_75t_L g607 ( 
.A1(n_536),
.A2(n_224),
.B1(n_236),
.B2(n_218),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

INVx6_ASAP7_75t_L g609 ( 
.A(n_579),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_455),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_555),
.B(n_324),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_521),
.A2(n_434),
.B1(n_416),
.B2(n_432),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_520),
.B(n_432),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_549),
.A2(n_224),
.B1(n_236),
.B2(n_218),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_562),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_563),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_542),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_470),
.Y(n_618)
);

INVx6_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_524),
.B(n_436),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_585),
.B(n_439),
.C(n_436),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

AND2x2_ASAP7_75t_SL g624 ( 
.A(n_579),
.B(n_324),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_566),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_591),
.B(n_455),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_528),
.B(n_439),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_522),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_599),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_531),
.B(n_549),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_440),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_590),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_592),
.B(n_440),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_542),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_577),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_581),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_590),
.B(n_334),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_449),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_590),
.B(n_472),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_549),
.A2(n_251),
.B1(n_291),
.B2(n_267),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_530),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_517),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_457),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_530),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_594),
.B(n_449),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_596),
.A2(n_501),
.B1(n_503),
.B2(n_498),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_549),
.A2(n_251),
.B1(n_291),
.B2(n_267),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_549),
.B(n_460),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_597),
.A2(n_460),
.B1(n_466),
.B2(n_465),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_465),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_574),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_534),
.Y(n_655)
);

OAI22x1_ASAP7_75t_L g656 ( 
.A1(n_595),
.A2(n_501),
.B1(n_503),
.B2(n_498),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_599),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_541),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_334),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_518),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_536),
.B(n_466),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_541),
.B(n_469),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_534),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_548),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_588),
.B(n_354),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_525),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_601),
.A2(n_493),
.B1(n_478),
.B2(n_482),
.Y(n_667)
);

AND3x2_ASAP7_75t_L g668 ( 
.A(n_586),
.B(n_375),
.C(n_317),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_469),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_588),
.B(n_354),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_601),
.B(n_471),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_526),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_588),
.B(n_454),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_561),
.A2(n_317),
.B1(n_391),
.B2(n_375),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_572),
.B(n_471),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_527),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_537),
.B(n_478),
.Y(n_678)
);

BUFx4f_ASAP7_75t_L g679 ( 
.A(n_599),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_573),
.B(n_482),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_569),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_545),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_550),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_600),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_574),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_574),
.B(n_360),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_574),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_571),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_574),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_546),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

INVx4_ASAP7_75t_SL g692 ( 
.A(n_557),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_548),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_561),
.A2(n_391),
.B1(n_378),
.B2(n_379),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_561),
.B(n_486),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_552),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_554),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_573),
.Y(n_698)
);

BUFx4f_ASAP7_75t_L g699 ( 
.A(n_557),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_556),
.B(n_486),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_519),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_539),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_559),
.B(n_406),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_558),
.B(n_493),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_573),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_539),
.B(n_497),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_546),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_575),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_575),
.B(n_209),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_575),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_540),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_540),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_559),
.B(n_360),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_560),
.B(n_497),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_560),
.B(n_507),
.C(n_504),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_557),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_564),
.B(n_504),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_582),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_582),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_576),
.B(n_380),
.C(n_276),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_557),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_580),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_519),
.B(n_507),
.Y(n_725)
);

AO22x2_ASAP7_75t_L g726 ( 
.A1(n_557),
.A2(n_378),
.B1(n_379),
.B2(n_234),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_532),
.B(n_235),
.Y(n_727)
);

BUFx4f_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_580),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_532),
.B(n_509),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_571),
.Y(n_731)
);

CKINVDCx6p67_ASAP7_75t_R g732 ( 
.A(n_587),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_580),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_580),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_535),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_535),
.B(n_509),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_580),
.B(n_207),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_543),
.B(n_235),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_543),
.B(n_268),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_544),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_544),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_587),
.B(n_246),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_533),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_547),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_547),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_533),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_553),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_553),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_565),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_565),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_567),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_567),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_570),
.B(n_235),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_658),
.B(n_511),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_624),
.B(n_675),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_614),
.B(n_399),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_624),
.B(n_369),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_643),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_643),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_665),
.A2(n_385),
.B(n_304),
.C(n_345),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_646),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_675),
.B(n_214),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_698),
.B(n_220),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_604),
.B(n_511),
.Y(n_764)
);

BUFx12f_ASAP7_75t_L g765 ( 
.A(n_701),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_648),
.B(n_490),
.C(n_570),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_SL g767 ( 
.A(n_722),
.B(n_408),
.C(n_584),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_613),
.B(n_389),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_620),
.B(n_277),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_698),
.B(n_230),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_632),
.B(n_206),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_609),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_628),
.B(n_584),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_610),
.B(n_208),
.C(n_206),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_646),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_708),
.B(n_232),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_708),
.B(n_614),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_642),
.A2(n_337),
.B1(n_349),
.B2(n_376),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_642),
.B(n_238),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_L g781 ( 
.A1(n_627),
.A2(n_645),
.B1(n_650),
.B2(n_631),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_679),
.B(n_211),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_609),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_655),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_609),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_714),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_661),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_649),
.B(n_243),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_661),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_295),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_649),
.B(n_399),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_674),
.A2(n_265),
.B1(n_399),
.B2(n_407),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_680),
.B(n_248),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_702),
.B(n_257),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_719),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_663),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_605),
.B(n_593),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_679),
.B(n_211),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_605),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_705),
.B(n_264),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_674),
.A2(n_399),
.B1(n_339),
.B2(n_405),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_626),
.B(n_398),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_619),
.Y(n_803)
);

NOR2xp67_ASAP7_75t_L g804 ( 
.A(n_681),
.B(n_593),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_633),
.B(n_213),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_710),
.B(n_280),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_659),
.B(n_293),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_659),
.B(n_298),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_652),
.B(n_399),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_659),
.B(n_313),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_662),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_671),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_619),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_626),
.B(n_213),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_717),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_619),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_645),
.B(n_657),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_603),
.B(n_215),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_615),
.Y(n_819)
);

OAI221xp5_ASAP7_75t_L g820 ( 
.A1(n_706),
.A2(n_703),
.B1(n_637),
.B2(n_636),
.C(n_616),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_717),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_625),
.Y(n_822)
);

BUFx5_ASAP7_75t_L g823 ( 
.A(n_724),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_663),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_603),
.B(n_215),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_711),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_603),
.B(n_217),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_703),
.A2(n_342),
.B1(n_336),
.B2(n_348),
.C(n_351),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_659),
.B(n_367),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_608),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_694),
.A2(n_371),
.B1(n_374),
.B2(n_377),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_654),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_653),
.A2(n_395),
.B1(n_237),
.B2(n_239),
.Y(n_834)
);

NOR2x1p5_ASAP7_75t_L g835 ( 
.A(n_673),
.B(n_408),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_373),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_688),
.B(n_746),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_645),
.B(n_600),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_716),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_716),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_665),
.A2(n_538),
.B(n_223),
.C(n_323),
.Y(n_841)
);

INVxp67_ASAP7_75t_L g842 ( 
.A(n_678),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_606),
.A2(n_326),
.B1(n_404),
.B2(n_403),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_712),
.B(n_223),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_611),
.B(n_638),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_647),
.B(n_237),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_690),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_622),
.B(n_239),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_635),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_699),
.A2(n_328),
.B(n_256),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_611),
.B(n_241),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_635),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_721),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_700),
.B(n_241),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_721),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_611),
.B(n_245),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_611),
.B(n_245),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_720),
.Y(n_858)
);

AND2x2_ASAP7_75t_SL g859 ( 
.A(n_694),
.B(n_227),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_611),
.B(n_256),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_678),
.A2(n_332),
.B1(n_272),
.B2(n_307),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_629),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_644),
.B(n_272),
.Y(n_863)
);

OAI22x1_ASAP7_75t_R g864 ( 
.A1(n_744),
.A2(n_538),
.B1(n_404),
.B2(n_403),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_664),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_660),
.B(n_307),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_SL g867 ( 
.A(n_748),
.B(n_227),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_667),
.B(n_310),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_669),
.A2(n_332),
.B(n_310),
.C(n_397),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_664),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_735),
.B(n_749),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_739),
.B(n_320),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_749),
.B(n_244),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_666),
.B(n_320),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_693),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_607),
.A2(n_402),
.B1(n_400),
.B2(n_249),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_651),
.B(n_323),
.Y(n_877)
);

BUFx6f_ASAP7_75t_SL g878 ( 
.A(n_684),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_672),
.B(n_328),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_676),
.Y(n_880)
);

NOR2x1p5_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_253),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_701),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_607),
.A2(n_402),
.B1(n_400),
.B2(n_253),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_677),
.B(n_341),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_682),
.B(n_341),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_683),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_693),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_731),
.Y(n_888)
);

AND2x6_ASAP7_75t_SL g889 ( 
.A(n_742),
.B(n_745),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_691),
.B(n_344),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_718),
.A2(n_397),
.B(n_396),
.Y(n_891)
);

AOI221xp5_ASAP7_75t_L g892 ( 
.A1(n_722),
.A2(n_309),
.B1(n_311),
.B2(n_314),
.C(n_315),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_684),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_R g894 ( 
.A(n_740),
.B(n_396),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_607),
.A2(n_382),
.B1(n_308),
.B2(n_309),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_696),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_704),
.B(n_344),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_715),
.B(n_346),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_748),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_726),
.A2(n_709),
.B1(n_733),
.B2(n_729),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_697),
.B(n_346),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_727),
.B(n_347),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_654),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_709),
.B(n_347),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_748),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_727),
.B(n_381),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_709),
.B(n_381),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_738),
.B(n_386),
.Y(n_908)
);

OAI22xp33_ASAP7_75t_L g909 ( 
.A1(n_618),
.A2(n_326),
.B1(n_314),
.B2(n_315),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_652),
.B(n_386),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_725),
.B(n_330),
.C(n_319),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_741),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_SL g913 ( 
.A(n_748),
.B(n_244),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_652),
.B(n_387),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_670),
.B(n_387),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_618),
.B(n_394),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_778),
.A2(n_718),
.B(n_695),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_826),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_842),
.B(n_612),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_755),
.B(n_670),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_769),
.B(n_639),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_757),
.A2(n_723),
.B(n_833),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_833),
.A2(n_723),
.B(n_652),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_845),
.A2(n_686),
.B(n_737),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_763),
.A2(n_776),
.B(n_770),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_769),
.B(n_726),
.Y(n_926)
);

O2A1O1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_790),
.A2(n_738),
.B(n_753),
.C(n_713),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_790),
.A2(n_736),
.B1(n_730),
.B2(n_753),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_802),
.A2(n_752),
.B1(n_751),
.B2(n_747),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_802),
.A2(n_728),
.B(n_686),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_815),
.B(n_734),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_814),
.A2(n_734),
.B(n_713),
.C(n_750),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_768),
.B(n_726),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_815),
.Y(n_934)
);

AOI21x1_ASAP7_75t_L g935 ( 
.A1(n_807),
.A2(n_641),
.B(n_618),
.Y(n_935)
);

INVx4_ASAP7_75t_L g936 ( 
.A(n_815),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_808),
.A2(n_641),
.B(n_656),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_903),
.A2(n_685),
.B(n_689),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_903),
.A2(n_685),
.B(n_689),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_793),
.A2(n_654),
.B(n_687),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_787),
.B(n_750),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_762),
.A2(n_621),
.B(n_623),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_810),
.A2(n_641),
.B(n_602),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_814),
.B(n_740),
.C(n_741),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_830),
.A2(n_654),
.B(n_687),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_836),
.A2(n_687),
.B(n_617),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_772),
.A2(n_687),
.B(n_617),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_783),
.A2(n_602),
.B(n_623),
.Y(n_948)
);

AO22x1_ASAP7_75t_L g949 ( 
.A1(n_848),
.A2(n_743),
.B1(n_382),
.B2(n_340),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_785),
.A2(n_813),
.B(n_803),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_828),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_768),
.B(n_621),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_758),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_900),
.A2(n_788),
.B(n_780),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_816),
.A2(n_847),
.B(n_791),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_754),
.B(n_743),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_869),
.A2(n_742),
.B(n_668),
.C(n_244),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_795),
.B(n_690),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_764),
.B(n_742),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_839),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_786),
.B(n_690),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_912),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_707),
.B1(n_690),
.B2(n_634),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_809),
.A2(n_634),
.B(n_707),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_799),
.B(n_388),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_847),
.A2(n_634),
.B(n_707),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_840),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_789),
.B(n_707),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_779),
.B(n_388),
.C(n_390),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_758),
.Y(n_970)
);

BUFx12f_ASAP7_75t_L g971 ( 
.A(n_765),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_900),
.A2(n_390),
.B(n_692),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_853),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_779),
.A2(n_308),
.B1(n_311),
.B2(n_319),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_759),
.A2(n_692),
.B(n_634),
.Y(n_975)
);

INVx3_ASAP7_75t_SL g976 ( 
.A(n_882),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_815),
.B(n_692),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_855),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_854),
.B(n_322),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_854),
.B(n_322),
.Y(n_980)
);

AO22x1_ASAP7_75t_L g981 ( 
.A1(n_848),
.A2(n_383),
.B1(n_340),
.B2(n_330),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_811),
.B(n_252),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_756),
.A2(n_383),
.B(n_141),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_891),
.A2(n_252),
.B(n_338),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_865),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_902),
.A2(n_261),
.B(n_394),
.C(n_4),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_821),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_756),
.A2(n_204),
.B(n_201),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_837),
.B(n_2),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_791),
.A2(n_193),
.B(n_175),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_821),
.B(n_170),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_801),
.A2(n_166),
.B(n_160),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_821),
.B(n_105),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_905),
.B(n_154),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_817),
.B(n_3),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_849),
.B(n_151),
.Y(n_996)
);

OAI321xp33_ASAP7_75t_L g997 ( 
.A1(n_843),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_888),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_821),
.B(n_146),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_801),
.A2(n_134),
.B(n_122),
.Y(n_1000)
);

NAND2x1p5_ASAP7_75t_L g1001 ( 
.A(n_899),
.B(n_119),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_849),
.B(n_852),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_794),
.A2(n_114),
.B(n_113),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_761),
.A2(n_92),
.B(n_90),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_775),
.A2(n_87),
.B(n_80),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_902),
.A2(n_906),
.B(n_908),
.C(n_841),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_870),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_781),
.A2(n_904),
.B(n_907),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_852),
.B(n_70),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_870),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_875),
.B(n_67),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_906),
.A2(n_9),
.B(n_10),
.C(n_13),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_846),
.B(n_17),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_875),
.B(n_23),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_820),
.A2(n_908),
.B1(n_819),
.B2(n_822),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_887),
.B(n_27),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_773),
.B(n_30),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_32),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_862),
.B(n_32),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_867),
.B(n_33),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_887),
.A2(n_33),
.B(n_34),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_823),
.B(n_34),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_832),
.A2(n_35),
.B(n_37),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_851),
.A2(n_38),
.B(n_40),
.C(n_41),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_777),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_823),
.B(n_42),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_832),
.A2(n_43),
.B(n_45),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_823),
.B(n_46),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_777),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_823),
.B(n_47),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_784),
.A2(n_824),
.B(n_796),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_SL g1032 ( 
.A1(n_910),
.A2(n_47),
.B(n_52),
.C(n_54),
.Y(n_1032)
);

AOI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_859),
.A2(n_58),
.B(n_59),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_859),
.A2(n_760),
.B(n_774),
.C(n_831),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_823),
.B(n_59),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_880),
.A2(n_60),
.B1(n_896),
.B2(n_886),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_823),
.B(n_796),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_838),
.B(n_805),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_858),
.A2(n_915),
.B(n_861),
.C(n_800),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_792),
.A2(n_895),
.B1(n_876),
.B2(n_883),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_868),
.B(n_877),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_824),
.B(n_792),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_806),
.B(n_844),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_L g1044 ( 
.A(n_893),
.B(n_797),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_863),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_809),
.A2(n_914),
.B(n_910),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_862),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_899),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_866),
.B(n_874),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_871),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_879),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_884),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_885),
.B(n_901),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_771),
.A2(n_890),
.B(n_857),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_856),
.A2(n_860),
.B(n_850),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_897),
.B(n_876),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_871),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_871),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_916),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_835),
.B(n_911),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_782),
.A2(n_798),
.B(n_827),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_873),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_894),
.B(n_878),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_SL g1064 ( 
.A(n_804),
.B(n_878),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_898),
.A2(n_818),
.B(n_825),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_873),
.B(n_881),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_913),
.A2(n_829),
.B(n_873),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_892),
.A2(n_895),
.B(n_883),
.C(n_766),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_909),
.B(n_894),
.Y(n_1070)
);

CKINVDCx8_ASAP7_75t_R g1071 ( 
.A(n_864),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_767),
.A2(n_802),
.B(n_790),
.C(n_755),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_912),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_762),
.A2(n_755),
.B(n_802),
.C(n_790),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_842),
.B(n_787),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_815),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_790),
.A2(n_802),
.B(n_755),
.C(n_762),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_842),
.B(n_787),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_778),
.A2(n_630),
.B(n_631),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_888),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_859),
.A2(n_802),
.B1(n_790),
.B2(n_755),
.Y(n_1085)
);

BUFx8_ASAP7_75t_L g1086 ( 
.A(n_878),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_755),
.B(n_769),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_778),
.A2(n_630),
.B(n_614),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1083),
.A2(n_1077),
.B(n_1076),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_SL g1092 ( 
.A1(n_919),
.A2(n_980),
.B(n_979),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1088),
.B(n_1079),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1072),
.B(n_984),
.C(n_928),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1080),
.A2(n_1087),
.B(n_1081),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1045),
.B(n_1051),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_955),
.A2(n_1031),
.B(n_945),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1075),
.B(n_1082),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_962),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_934),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_SL g1102 ( 
.A(n_971),
.Y(n_1102)
);

AOI21xp33_ASAP7_75t_L g1103 ( 
.A1(n_1040),
.A2(n_1074),
.B(n_1041),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1089),
.A2(n_920),
.B(n_954),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_924),
.A2(n_940),
.B(n_1037),
.Y(n_1105)
);

OAI22x1_ASAP7_75t_L g1106 ( 
.A1(n_969),
.A2(n_929),
.B1(n_1017),
.B2(n_941),
.Y(n_1106)
);

NAND2x1_ASAP7_75t_L g1107 ( 
.A(n_934),
.B(n_936),
.Y(n_1107)
);

NOR2x1_ASAP7_75t_L g1108 ( 
.A(n_944),
.B(n_1044),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1037),
.A2(n_966),
.B(n_948),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_SL g1110 ( 
.A1(n_1022),
.A2(n_1028),
.B(n_1026),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_920),
.B(n_1049),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_917),
.A2(n_922),
.B(n_942),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1008),
.A2(n_943),
.B(n_925),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1006),
.A2(n_933),
.B(n_926),
.Y(n_1114)
);

NAND2x1_ASAP7_75t_L g1115 ( 
.A(n_936),
.B(n_987),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1053),
.B(n_1052),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_976),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_1040),
.A2(n_1056),
.B(n_927),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_938),
.A2(n_939),
.B(n_947),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1084),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1048),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_950),
.A2(n_1055),
.B(n_999),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1013),
.A2(n_1068),
.B(n_1018),
.C(n_921),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_993),
.A2(n_999),
.B(n_1046),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1043),
.B(n_968),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_993),
.A2(n_1011),
.B(n_977),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1011),
.A2(n_923),
.B(n_1054),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_968),
.B(n_921),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_933),
.A2(n_926),
.B(n_1033),
.Y(n_1129)
);

INVx6_ASAP7_75t_L g1130 ( 
.A(n_1086),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_930),
.A2(n_1042),
.B(n_952),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1022),
.A2(n_1035),
.B(n_1030),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_1073),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1039),
.A2(n_961),
.B(n_958),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1029),
.A2(n_918),
.B(n_951),
.Y(n_1135)
);

BUFx8_ASAP7_75t_SL g1136 ( 
.A(n_1060),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_956),
.B(n_1059),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1015),
.B(n_958),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_961),
.A2(n_931),
.B(n_1061),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_1064),
.B(n_1071),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1047),
.B(n_960),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1067),
.A2(n_1034),
.B(n_1033),
.C(n_1065),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_987),
.A2(n_1078),
.B(n_1005),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_931),
.A2(n_1078),
.B(n_932),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1019),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1070),
.A2(n_1030),
.B1(n_1026),
.B2(n_1028),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1070),
.B(n_1050),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_967),
.B(n_973),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_SL g1150 ( 
.A1(n_1035),
.A2(n_1027),
.B(n_1023),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1048),
.B(n_1058),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_985),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1060),
.A2(n_1002),
.B1(n_1038),
.B2(n_995),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_978),
.B(n_1010),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_1058),
.B(n_1050),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_989),
.B(n_1019),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1007),
.B(n_1025),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1004),
.A2(n_972),
.B(n_963),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_953),
.B(n_970),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_992),
.A2(n_1000),
.B(n_996),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1014),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1016),
.B(n_1036),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1062),
.B(n_1057),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1009),
.A2(n_983),
.B(n_988),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_SL g1165 ( 
.A(n_935),
.B(n_937),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_990),
.A2(n_991),
.B(n_1003),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_991),
.A2(n_982),
.B(n_1001),
.Y(n_1167)
);

INVx8_ASAP7_75t_L g1168 ( 
.A(n_1066),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1062),
.B(n_1066),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1001),
.A2(n_1020),
.B(n_957),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_959),
.B(n_949),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1012),
.A2(n_986),
.B(n_997),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_965),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1021),
.A2(n_974),
.A3(n_1032),
.B(n_1024),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1069),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_981),
.B(n_974),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_994),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1076),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_1086),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1085),
.A2(n_980),
.B1(n_979),
.B2(n_790),
.Y(n_1181)
);

BUFx12f_ASAP7_75t_L g1182 ( 
.A(n_1086),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1085),
.A2(n_1040),
.B1(n_1088),
.B2(n_1068),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_928),
.B(n_1072),
.Y(n_1188)
);

O2A1O1Ixp5_ASAP7_75t_L g1189 ( 
.A1(n_1074),
.A2(n_984),
.B(n_1006),
.C(n_980),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1191)
);

INVx8_ASAP7_75t_L g1192 ( 
.A(n_1019),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1079),
.A2(n_1072),
.B(n_1074),
.C(n_980),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1075),
.B(n_787),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_918),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1085),
.A2(n_1040),
.B1(n_1088),
.B2(n_1068),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1075),
.B(n_787),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1084),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_928),
.B(n_1072),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1006),
.A2(n_1008),
.A3(n_1034),
.B(n_932),
.Y(n_1207)
);

OAI22x1_ASAP7_75t_L g1208 ( 
.A1(n_928),
.A2(n_919),
.B1(n_969),
.B2(n_522),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1084),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1210)
);

OAI22x1_ASAP7_75t_L g1211 ( 
.A1(n_928),
.A2(n_919),
.B1(n_969),
.B2(n_522),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1048),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_934),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1029),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1079),
.A2(n_1072),
.B(n_1074),
.C(n_980),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1083),
.A2(n_699),
.B(n_718),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1029),
.Y(n_1218)
);

AOI211xp5_ASAP7_75t_L g1219 ( 
.A1(n_919),
.A2(n_802),
.B(n_790),
.C(n_1040),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1220)
);

AO32x2_ASAP7_75t_L g1221 ( 
.A1(n_1040),
.A2(n_834),
.A3(n_974),
.B1(n_1058),
.B2(n_936),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_918),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_962),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1088),
.B(n_1085),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1029),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1075),
.B(n_812),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_962),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_928),
.B(n_1072),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_975),
.A2(n_964),
.B(n_946),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1057),
.B(n_849),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_928),
.B(n_1072),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_918),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1111),
.B(n_1125),
.Y(n_1235)
);

NOR2x1_ASAP7_75t_SL g1236 ( 
.A(n_1161),
.B(n_1148),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1181),
.A2(n_1095),
.B1(n_1211),
.B2(n_1208),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_1117),
.B(n_1204),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1186),
.A2(n_1202),
.B1(n_1106),
.B2(n_1176),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_L g1240 ( 
.A(n_1209),
.B(n_1097),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1101),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1149),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1120),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1101),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1154),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1219),
.A2(n_1092),
.B1(n_1123),
.B2(n_1111),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1189),
.A2(n_1158),
.B(n_1142),
.C(n_1193),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1154),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1227),
.B(n_1099),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1200),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1116),
.B(n_1097),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1222),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1090),
.B(n_1180),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1224),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1137),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1090),
.B(n_1180),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1199),
.A2(n_1203),
.B1(n_1186),
.B2(n_1202),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1116),
.A2(n_1220),
.B1(n_1225),
.B2(n_1183),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1156),
.B(n_1146),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1153),
.B(n_1171),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1091),
.A2(n_1112),
.B(n_1096),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1100),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1234),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1184),
.A2(n_1187),
.B1(n_1201),
.B2(n_1212),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1182),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1121),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1157),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1157),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1133),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1214),
.Y(n_1273)
);

AO21x1_ASAP7_75t_L g1274 ( 
.A1(n_1188),
.A2(n_1233),
.B(n_1230),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1141),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1229),
.B(n_1187),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1094),
.A2(n_1231),
.B(n_1228),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1201),
.A2(n_1206),
.B1(n_1210),
.B2(n_1212),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1121),
.B(n_1213),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1206),
.B(n_1210),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1118),
.A2(n_1104),
.B(n_1216),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1168),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1213),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1213),
.B(n_1163),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1175),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1192),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1176),
.A2(n_1130),
.B1(n_1173),
.B2(n_1179),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1192),
.B(n_1168),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1138),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1177),
.B(n_1114),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1114),
.B(n_1221),
.Y(n_1292)
);

BUFx12f_ASAP7_75t_L g1293 ( 
.A(n_1130),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1221),
.B(n_1140),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1221),
.B(n_1155),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1192),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1128),
.B(n_1093),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1215),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1168),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1218),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1205),
.A2(n_1172),
.B1(n_1103),
.B2(n_1129),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1162),
.B(n_1147),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1130),
.B(n_1151),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1226),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1155),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1151),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1162),
.A2(n_1108),
.B1(n_1170),
.B2(n_1147),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1214),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1102),
.Y(n_1310)
);

AOI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1103),
.A2(n_1172),
.B(n_1118),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1136),
.Y(n_1312)
);

INVx5_ASAP7_75t_L g1313 ( 
.A(n_1144),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_L g1314 ( 
.A1(n_1178),
.A2(n_1113),
.B(n_1132),
.C(n_1131),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1185),
.A2(n_1190),
.B(n_1196),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1165),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1129),
.B(n_1174),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1134),
.A2(n_1160),
.B(n_1167),
.C(n_1178),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1107),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1115),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1174),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1135),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1110),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1174),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1207),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1139),
.B(n_1152),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1124),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1207),
.B(n_1145),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1126),
.B(n_1122),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1105),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1109),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1119),
.Y(n_1332)
);

NAND2x1_ASAP7_75t_L g1333 ( 
.A(n_1150),
.B(n_1166),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1127),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1194),
.B(n_1223),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1191),
.A2(n_1197),
.B(n_1198),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1098),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_SL g1338 ( 
.A(n_1164),
.B(n_1217),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1092),
.A2(n_802),
.B(n_790),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1121),
.Y(n_1340)
);

NOR2x1_ASAP7_75t_R g1341 ( 
.A(n_1130),
.B(n_605),
.Y(n_1341)
);

AND2x2_ASAP7_75t_SL g1342 ( 
.A(n_1181),
.B(n_1085),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1149),
.Y(n_1344)
);

INVx8_ASAP7_75t_L g1345 ( 
.A(n_1168),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1092),
.B(n_787),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1149),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1092),
.A2(n_1219),
.B(n_1181),
.C(n_1072),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1219),
.A2(n_980),
.B(n_979),
.C(n_790),
.Y(n_1350)
);

NAND2x1p5_ASAP7_75t_L g1351 ( 
.A(n_1101),
.B(n_934),
.Y(n_1351)
);

NOR2x1_ASAP7_75t_L g1352 ( 
.A(n_1117),
.B(n_740),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1091),
.A2(n_1112),
.B(n_1096),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1224),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1092),
.B(n_787),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1227),
.B(n_1099),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1204),
.B(n_748),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1224),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1149),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1149),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1091),
.A2(n_1112),
.B(n_1096),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1120),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1101),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1149),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1100),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1117),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1121),
.Y(n_1369)
);

OR2x6_ASAP7_75t_L g1370 ( 
.A(n_1192),
.B(n_1168),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1117),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1094),
.A2(n_1195),
.B(n_1194),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1181),
.A2(n_1040),
.B1(n_980),
.B2(n_979),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1120),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1149),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1169),
.B(n_1232),
.Y(n_1376)
);

BUFx2_ASAP7_75t_SL g1377 ( 
.A(n_1117),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1094),
.A2(n_1195),
.B(n_1194),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1091),
.A2(n_1112),
.B(n_1096),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1092),
.B(n_787),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1120),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1120),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1100),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1121),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1181),
.A2(n_1040),
.B1(n_980),
.B2(n_979),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1091),
.A2(n_1112),
.B(n_1096),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1111),
.B(n_1125),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1092),
.A2(n_1219),
.B(n_1123),
.C(n_1079),
.Y(n_1388)
);

INVx3_ASAP7_75t_SL g1389 ( 
.A(n_1130),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1120),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1339),
.A2(n_1342),
.B1(n_1373),
.B2(n_1385),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1258),
.B(n_1294),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1237),
.A2(n_1261),
.B1(n_1247),
.B2(n_1380),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1247),
.A2(n_1346),
.B1(n_1356),
.B2(n_1239),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1265),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1313),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1288),
.A2(n_1303),
.B1(n_1291),
.B2(n_1250),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1303),
.A2(n_1357),
.B1(n_1281),
.B2(n_1263),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1251),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1371),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1296),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1324),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1313),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1313),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1369),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1368),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1253),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1270),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1369),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1252),
.B(n_1290),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1271),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1262),
.A2(n_1362),
.B(n_1354),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1242),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1272),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1246),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1349),
.B(n_1290),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1321),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1277),
.A2(n_1378),
.B(n_1372),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1235),
.B(n_1387),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1344),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1348),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1360),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1289),
.B(n_1370),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1350),
.A2(n_1388),
.B(n_1308),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1249),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1313),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1359),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1361),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1335),
.A2(n_1333),
.B(n_1336),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1366),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1274),
.A2(n_1302),
.B1(n_1311),
.B2(n_1276),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1335),
.A2(n_1315),
.B(n_1336),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1375),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1235),
.A2(n_1387),
.B1(n_1298),
.B2(n_1256),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1311),
.A2(n_1281),
.B1(n_1259),
.B2(n_1266),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1369),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1256),
.B(n_1275),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1359),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1292),
.B(n_1254),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1345),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1243),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1254),
.B(n_1257),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1322),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1322),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1322),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1367),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1314),
.A2(n_1248),
.B(n_1354),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1355),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1389),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1293),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1259),
.A2(n_1278),
.B1(n_1266),
.B2(n_1323),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1240),
.A2(n_1286),
.B1(n_1383),
.B2(n_1298),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1286),
.A2(n_1383),
.B1(n_1388),
.B2(n_1280),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1257),
.A2(n_1264),
.B1(n_1280),
.B2(n_1282),
.Y(n_1454)
);

AO21x1_ASAP7_75t_SL g1455 ( 
.A1(n_1328),
.A2(n_1264),
.B(n_1329),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_SL g1456 ( 
.A(n_1374),
.Y(n_1456)
);

AO21x1_ASAP7_75t_L g1457 ( 
.A1(n_1326),
.A2(n_1278),
.B(n_1328),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1299),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1301),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1260),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1314),
.A2(n_1386),
.B(n_1379),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1352),
.A2(n_1364),
.B1(n_1343),
.B2(n_1347),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1244),
.A2(n_1268),
.B1(n_1376),
.B2(n_1347),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1289),
.B(n_1370),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1295),
.B(n_1317),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1381),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1267),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1312),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1305),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1330),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1382),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1310),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1236),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1255),
.Y(n_1474)
);

BUFx8_ASAP7_75t_L g1475 ( 
.A(n_1287),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1241),
.B(n_1309),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1241),
.B(n_1309),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1327),
.B(n_1331),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1244),
.A2(n_1343),
.B1(n_1353),
.B2(n_1268),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1238),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1353),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1245),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1345),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1334),
.A2(n_1332),
.B(n_1337),
.Y(n_1484)
);

CKINVDCx11_ASAP7_75t_R g1485 ( 
.A(n_1340),
.Y(n_1485)
);

NAND2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1327),
.B(n_1331),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1273),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1304),
.A2(n_1358),
.B1(n_1370),
.B2(n_1289),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1273),
.B(n_1365),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1340),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1364),
.A2(n_1376),
.B1(n_1285),
.B2(n_1377),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1337),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1307),
.B(n_1306),
.Y(n_1493)
);

NAND2x1_ASAP7_75t_L g1494 ( 
.A(n_1332),
.B(n_1334),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1285),
.Y(n_1495)
);

AO21x1_ASAP7_75t_SL g1496 ( 
.A1(n_1297),
.A2(n_1338),
.B(n_1318),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1345),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1306),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_SL g1499 ( 
.A(n_1279),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1363),
.B(n_1390),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1283),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1306),
.B(n_1304),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1304),
.A2(n_1300),
.B1(n_1269),
.B2(n_1284),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1351),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1351),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1384),
.Y(n_1506)
);

AOI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1320),
.A2(n_1316),
.B(n_1279),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1341),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1316),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1319),
.A2(n_1269),
.B(n_1284),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1319),
.Y(n_1511)
);

INVx6_ASAP7_75t_L g1512 ( 
.A(n_1369),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1272),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1371),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1267),
.Y(n_1515)
);

BUFx10_ASAP7_75t_L g1516 ( 
.A(n_1368),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1339),
.A2(n_1342),
.B1(n_1181),
.B2(n_1373),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1371),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1369),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1277),
.A2(n_1378),
.B(n_1372),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1339),
.A2(n_1342),
.B1(n_1181),
.B2(n_1373),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1325),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1339),
.A2(n_1092),
.B1(n_1181),
.B2(n_532),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1321),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1457),
.A2(n_1402),
.A3(n_1412),
.B(n_1522),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1475),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1457),
.A2(n_1424),
.B(n_1432),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1465),
.B(n_1439),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1502),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1470),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1465),
.B(n_1439),
.Y(n_1532)
);

BUFx4f_ASAP7_75t_SL g1533 ( 
.A(n_1467),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1441),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1492),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1454),
.B(n_1392),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1514),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1400),
.B(n_1518),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1441),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1392),
.B(n_1442),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1427),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1438),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1443),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1448),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1442),
.B(n_1416),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1429),
.B(n_1478),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1502),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1416),
.B(n_1435),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1453),
.B(n_1451),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1407),
.B(n_1415),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1446),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1425),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1408),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1414),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_SL g1555 ( 
.A1(n_1423),
.A2(n_1464),
.B(n_1436),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1391),
.A2(n_1521),
.B(n_1517),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1407),
.B(n_1455),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1400),
.B(n_1518),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1411),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1474),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1434),
.B(n_1447),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1455),
.B(n_1395),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1401),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1484),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1418),
.A2(n_1520),
.B(n_1431),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1512),
.Y(n_1566)
);

AOI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1494),
.A2(n_1507),
.B(n_1473),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1494),
.A2(n_1478),
.B(n_1486),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1394),
.B(n_1393),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1437),
.B(n_1413),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1444),
.B(n_1445),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1513),
.Y(n_1572)
);

AO21x2_ASAP7_75t_L g1573 ( 
.A1(n_1507),
.A2(n_1509),
.B(n_1399),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1420),
.B(n_1421),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1423),
.A2(n_1464),
.B(n_1409),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1461),
.B(n_1460),
.Y(n_1576)
);

BUFx3_ASAP7_75t_L g1577 ( 
.A(n_1466),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1422),
.B(n_1428),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1444),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1523),
.B(n_1452),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1397),
.B(n_1398),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1493),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1481),
.B(n_1458),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1466),
.Y(n_1585)
);

INVxp33_ASAP7_75t_L g1586 ( 
.A(n_1514),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1459),
.B(n_1469),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1417),
.B(n_1524),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1495),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1512),
.Y(n_1590)
);

AO21x2_ASAP7_75t_L g1591 ( 
.A1(n_1488),
.A2(n_1482),
.B(n_1487),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1511),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1406),
.B(n_1480),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1511),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1476),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1476),
.B(n_1489),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1500),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1477),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1491),
.B(n_1477),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1504),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1549),
.A2(n_1462),
.B1(n_1508),
.B2(n_1463),
.C(n_1479),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1527),
.B(n_1496),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1524),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1569),
.A2(n_1464),
.B1(n_1423),
.B2(n_1501),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1540),
.B(n_1417),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1546),
.B(n_1396),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1527),
.B(n_1489),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1546),
.B(n_1396),
.Y(n_1610)
);

INVx5_ASAP7_75t_L g1611 ( 
.A(n_1546),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1576),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1546),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1540),
.B(n_1403),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1576),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1564),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1557),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1536),
.B(n_1403),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1531),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1564),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1531),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1573),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1557),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1546),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1571),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1556),
.A2(n_1503),
.B(n_1426),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1535),
.B(n_1426),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1532),
.B(n_1404),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1573),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1532),
.B(n_1404),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1562),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1525),
.B(n_1404),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1525),
.B(n_1498),
.Y(n_1633)
);

AND2x2_ASAP7_75t_SL g1634 ( 
.A(n_1549),
.B(n_1436),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1562),
.B(n_1504),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1561),
.B(n_1505),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1525),
.B(n_1505),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1525),
.Y(n_1638)
);

INVx4_ASAP7_75t_R g1639 ( 
.A(n_1534),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1582),
.A2(n_1468),
.B1(n_1449),
.B2(n_1516),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_SL g1641 ( 
.A(n_1561),
.B(n_1436),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1528),
.B(n_1510),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1528),
.B(n_1510),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1607),
.B(n_1544),
.Y(n_1644)
);

NAND3xp33_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1530),
.C(n_1548),
.Y(n_1645)
);

NOR3xp33_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1537),
.C(n_1599),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1541),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1640),
.A2(n_1548),
.B(n_1586),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1614),
.B(n_1542),
.Y(n_1649)
);

NOR3xp33_ASAP7_75t_L g1650 ( 
.A(n_1626),
.B(n_1597),
.C(n_1588),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1640),
.A2(n_1588),
.B1(n_1572),
.B2(n_1570),
.C(n_1560),
.Y(n_1651)
);

AND2x2_ASAP7_75t_SL g1652 ( 
.A(n_1634),
.B(n_1545),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1631),
.B(n_1596),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1605),
.B(n_1554),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1634),
.A2(n_1529),
.B1(n_1547),
.B2(n_1526),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1601),
.A2(n_1567),
.B(n_1580),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1626),
.A2(n_1593),
.B(n_1558),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1623),
.B(n_1583),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1605),
.B(n_1595),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1606),
.A2(n_1584),
.B(n_1574),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1634),
.A2(n_1529),
.B1(n_1547),
.B2(n_1526),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1634),
.A2(n_1526),
.B1(n_1533),
.B2(n_1468),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1595),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1565),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_SL g1665 ( 
.A1(n_1606),
.A2(n_1538),
.B(n_1551),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1628),
.B(n_1598),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_L g1668 ( 
.A(n_1629),
.B(n_1589),
.C(n_1587),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1618),
.A2(n_1555),
.B1(n_1575),
.B2(n_1585),
.C(n_1577),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1602),
.B(n_1555),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1641),
.A2(n_1575),
.B(n_1600),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1618),
.B(n_1592),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1604),
.A2(n_1440),
.B(n_1578),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1641),
.A2(n_1499),
.B(n_1409),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1642),
.B(n_1565),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1601),
.B(n_1622),
.C(n_1629),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1622),
.A2(n_1577),
.B1(n_1539),
.B2(n_1585),
.C(n_1526),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1642),
.B(n_1565),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1643),
.B(n_1579),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1594),
.Y(n_1681)
);

AOI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1633),
.A2(n_1612),
.B1(n_1637),
.B2(n_1632),
.C(n_1615),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1543),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1635),
.B(n_1550),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1624),
.A2(n_1480),
.B1(n_1590),
.B2(n_1566),
.C(n_1483),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1633),
.B(n_1559),
.C(n_1563),
.D(n_1552),
.Y(n_1686)
);

NAND3xp33_ASAP7_75t_SL g1687 ( 
.A(n_1633),
.B(n_1406),
.C(n_1501),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1635),
.A2(n_1591),
.B1(n_1449),
.B2(n_1499),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1617),
.B(n_1543),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1635),
.B(n_1550),
.Y(n_1690)
);

NAND3xp33_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1559),
.C(n_1563),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1635),
.B(n_1552),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1625),
.B(n_1516),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1604),
.A2(n_1440),
.B(n_1567),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1619),
.B(n_1553),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1621),
.B(n_1553),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1673),
.B(n_1612),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1696),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1681),
.B(n_1615),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1697),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1680),
.B(n_1609),
.Y(n_1702)
);

NAND4xp25_ASAP7_75t_L g1703 ( 
.A(n_1646),
.B(n_1627),
.C(n_1636),
.D(n_1609),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1683),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1695),
.B(n_1621),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1650),
.B(n_1638),
.C(n_1627),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1693),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1687),
.A2(n_1625),
.B1(n_1610),
.B2(n_1608),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1683),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1691),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1692),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1663),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1656),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1656),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1671),
.B(n_1602),
.Y(n_1715)
);

AND2x4_ASAP7_75t_SL g1716 ( 
.A(n_1689),
.B(n_1608),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1656),
.Y(n_1717)
);

BUFx2_ASAP7_75t_SL g1718 ( 
.A(n_1664),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1656),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1689),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1653),
.B(n_1652),
.Y(n_1721)
);

NAND2x1_ASAP7_75t_L g1722 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1649),
.B(n_1616),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1682),
.B(n_1616),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1666),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1652),
.B(n_1658),
.Y(n_1726)
);

NAND2x1_ASAP7_75t_L g1727 ( 
.A(n_1675),
.B(n_1639),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1667),
.B(n_1613),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1669),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1684),
.Y(n_1730)
);

INVxp67_ASAP7_75t_SL g1731 ( 
.A(n_1677),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1647),
.B(n_1616),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1664),
.B(n_1611),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1690),
.B(n_1620),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1644),
.B(n_1620),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1668),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1662),
.B(n_1608),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1711),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1699),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1721),
.B(n_1671),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1711),
.B(n_1654),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1706),
.A2(n_1648),
.B(n_1657),
.C(n_1645),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1699),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1701),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1705),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1701),
.B(n_1659),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1705),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1713),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1731),
.B(n_1660),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1704),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1710),
.B(n_1724),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1704),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1716),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1721),
.B(n_1676),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1710),
.B(n_1679),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1735),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1712),
.B(n_1660),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1735),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

INVx3_ASAP7_75t_R g1761 ( 
.A(n_1715),
.Y(n_1761)
);

NOR2xp67_ASAP7_75t_L g1762 ( 
.A(n_1706),
.B(n_1672),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1726),
.B(n_1679),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1723),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1723),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1714),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1726),
.B(n_1611),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1712),
.B(n_1725),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1724),
.B(n_1686),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1722),
.B(n_1611),
.Y(n_1770)
);

NOR2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1722),
.B(n_1645),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1714),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1718),
.B(n_1611),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1729),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1734),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1714),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1709),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1707),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1732),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1709),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1700),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1748),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1779),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1739),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1748),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1749),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1740),
.B(n_1767),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1756),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1743),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1744),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1738),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1771),
.A2(n_1737),
.B1(n_1703),
.B2(n_1708),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1758),
.B(n_1736),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1769),
.B(n_1736),
.Y(n_1796)
);

OAI311xp33_ASAP7_75t_L g1797 ( 
.A1(n_1742),
.A2(n_1703),
.A3(n_1665),
.B1(n_1651),
.C1(n_1688),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1753),
.B(n_1715),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1698),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1751),
.B(n_1729),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1751),
.B(n_1762),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1730),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1738),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1755),
.B(n_1698),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1753),
.B(n_1715),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1740),
.B(n_1718),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1756),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1760),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1750),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1750),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1755),
.B(n_1702),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1752),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1752),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1760),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1778),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1716),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1741),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1781),
.B(n_1728),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1778),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1763),
.B(n_1716),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1782),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1745),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1766),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1770),
.B(n_1727),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1746),
.B(n_1728),
.Y(n_1825)
);

INVxp67_ASAP7_75t_L g1826 ( 
.A(n_1745),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1747),
.B(n_1702),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1747),
.B(n_1685),
.C(n_1668),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1782),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1803),
.Y(n_1830)
);

AND2x2_ASAP7_75t_SL g1831 ( 
.A(n_1801),
.B(n_1737),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1788),
.B(n_1817),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1806),
.B(n_1783),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1795),
.B(n_1764),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1803),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1785),
.B(n_1467),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1796),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1796),
.B(n_1765),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1784),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1806),
.B(n_1789),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1819),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1789),
.B(n_1783),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1819),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1829),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1824),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1794),
.A2(n_1737),
.B1(n_1759),
.B2(n_1757),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1799),
.B(n_1775),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1829),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1828),
.A2(n_1777),
.B1(n_1715),
.B2(n_1770),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1799),
.B(n_1768),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1822),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1798),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1804),
.B(n_1776),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1816),
.B(n_1770),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1797),
.A2(n_1727),
.B(n_1773),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1824),
.B(n_1773),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1804),
.B(n_1766),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1784),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1793),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1802),
.A2(n_1670),
.B1(n_1678),
.B2(n_1661),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1787),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_SL g1863 ( 
.A1(n_1816),
.A2(n_1611),
.B1(n_1763),
.B2(n_1733),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1776),
.Y(n_1864)
);

AOI22x1_ASAP7_75t_L g1865 ( 
.A1(n_1826),
.A2(n_1515),
.B1(n_1450),
.B2(n_1506),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1787),
.Y(n_1866)
);

CKINVDCx16_ASAP7_75t_R g1867 ( 
.A(n_1824),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1786),
.B(n_1754),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1836),
.B(n_1515),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1841),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1852),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1837),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1841),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1831),
.B(n_1798),
.Y(n_1874)
);

XNOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1865),
.B(n_1824),
.Y(n_1875)
);

OAI31xp33_ASAP7_75t_SL g1876 ( 
.A1(n_1856),
.A2(n_1805),
.A3(n_1798),
.B(n_1820),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1867),
.B(n_1832),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1846),
.A2(n_1820),
.B1(n_1805),
.B2(n_1825),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1843),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1843),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_L g1881 ( 
.A1(n_1851),
.A2(n_1805),
.B(n_1791),
.C(n_1792),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1831),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1844),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1851),
.B(n_1818),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1849),
.A2(n_1811),
.B1(n_1674),
.B2(n_1827),
.Y(n_1885)
);

OAI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1845),
.A2(n_1810),
.B(n_1809),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1838),
.B(n_1811),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_SL g1888 ( 
.A1(n_1845),
.A2(n_1761),
.B(n_1821),
.C(n_1815),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1847),
.B(n_1812),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1861),
.A2(n_1655),
.B1(n_1694),
.B2(n_1717),
.C(n_1719),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1844),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1840),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1833),
.B(n_1754),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1845),
.B(n_1813),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1840),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1848),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1848),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1892),
.B(n_1833),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1874),
.A2(n_1857),
.B1(n_1855),
.B2(n_1842),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1877),
.B(n_1834),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1877),
.B(n_1853),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_SL g1902 ( 
.A(n_1882),
.B(n_1865),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1894),
.B(n_1857),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1874),
.A2(n_1860),
.B1(n_1835),
.B2(n_1830),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1871),
.B(n_1842),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1870),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1873),
.Y(n_1907)
);

INVxp67_ASAP7_75t_SL g1908 ( 
.A(n_1875),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_L g1909 ( 
.A(n_1872),
.B(n_1850),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1895),
.B(n_1855),
.Y(n_1910)
);

INVxp33_ASAP7_75t_L g1911 ( 
.A(n_1869),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1893),
.B(n_1847),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1887),
.B(n_1868),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1876),
.B(n_1857),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1879),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1889),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_L g1917 ( 
.A(n_1869),
.B(n_1839),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1880),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1883),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1886),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1898),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1909),
.A2(n_1888),
.B(n_1890),
.Y(n_1922)
);

NOR4xp25_ASAP7_75t_L g1923 ( 
.A(n_1909),
.B(n_1888),
.C(n_1896),
.D(n_1891),
.Y(n_1923)
);

AOI211xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1908),
.A2(n_1881),
.B(n_1878),
.C(n_1884),
.Y(n_1924)
);

XOR2xp5_ASAP7_75t_L g1925 ( 
.A(n_1911),
.B(n_1885),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_SL g1926 ( 
.A(n_1902),
.B(n_1863),
.C(n_1850),
.Y(n_1926)
);

XOR2xp5_ASAP7_75t_L g1927 ( 
.A(n_1911),
.B(n_1899),
.Y(n_1927)
);

NOR3xp33_ASAP7_75t_L g1928 ( 
.A(n_1901),
.B(n_1920),
.C(n_1900),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_SL g1929 ( 
.A1(n_1901),
.A2(n_1897),
.B(n_1853),
.Y(n_1929)
);

NOR3xp33_ASAP7_75t_L g1930 ( 
.A(n_1900),
.B(n_1450),
.C(n_1471),
.Y(n_1930)
);

O2A1O1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1904),
.A2(n_1866),
.B(n_1862),
.C(n_1859),
.Y(n_1931)
);

NOR3x1_ASAP7_75t_L g1932 ( 
.A(n_1905),
.B(n_1858),
.C(n_1854),
.Y(n_1932)
);

NAND3xp33_ASAP7_75t_L g1933 ( 
.A(n_1904),
.B(n_1859),
.C(n_1839),
.Y(n_1933)
);

OAI21xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1914),
.A2(n_1858),
.B(n_1854),
.Y(n_1934)
);

AOI221xp5_ASAP7_75t_L g1935 ( 
.A1(n_1923),
.A2(n_1916),
.B1(n_1910),
.B2(n_1919),
.C(n_1918),
.Y(n_1935)
);

OAI21xp33_ASAP7_75t_L g1936 ( 
.A1(n_1934),
.A2(n_1917),
.B(n_1912),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1921),
.Y(n_1937)
);

OAI211xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1924),
.A2(n_1913),
.B(n_1907),
.C(n_1906),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1922),
.A2(n_1903),
.B(n_1915),
.Y(n_1939)
);

NAND4xp75_ASAP7_75t_L g1940 ( 
.A(n_1932),
.B(n_1903),
.C(n_1866),
.D(n_1862),
.Y(n_1940)
);

AO22x1_ASAP7_75t_L g1941 ( 
.A1(n_1928),
.A2(n_1903),
.B1(n_1475),
.B2(n_1807),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1927),
.B(n_1864),
.Y(n_1942)
);

NOR2x1_ASAP7_75t_L g1943 ( 
.A(n_1933),
.B(n_1925),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1931),
.Y(n_1944)
);

NAND3xp33_ASAP7_75t_L g1945 ( 
.A(n_1929),
.B(n_1930),
.C(n_1926),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1921),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1922),
.A2(n_1864),
.B1(n_1720),
.B2(n_1814),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1936),
.A2(n_1807),
.B(n_1790),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1937),
.Y(n_1949)
);

OAI21xp33_ASAP7_75t_SL g1950 ( 
.A1(n_1940),
.A2(n_1808),
.B(n_1790),
.Y(n_1950)
);

NAND3xp33_ASAP7_75t_L g1951 ( 
.A(n_1935),
.B(n_1471),
.C(n_1808),
.Y(n_1951)
);

NOR3xp33_ASAP7_75t_L g1952 ( 
.A(n_1945),
.B(n_1490),
.C(n_1485),
.Y(n_1952)
);

NAND2x2_ASAP7_75t_L g1953 ( 
.A(n_1942),
.B(n_1497),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1939),
.B(n_1814),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_L g1955 ( 
.A(n_1944),
.B(n_1823),
.C(n_1490),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1949),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1954),
.B(n_1946),
.Y(n_1957)
);

NOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1951),
.B(n_1943),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1955),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1948),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1950),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1953),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1957),
.Y(n_1963)
);

INVx5_ASAP7_75t_L g1964 ( 
.A(n_1959),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1956),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1962),
.B(n_1952),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_L g1967 ( 
.A(n_1958),
.B(n_1938),
.C(n_1941),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1961),
.B(n_1947),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1964),
.Y(n_1969)
);

XOR2xp5_ASAP7_75t_L g1970 ( 
.A(n_1966),
.B(n_1959),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1964),
.A2(n_1960),
.B1(n_1823),
.B2(n_1772),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1963),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1969),
.Y(n_1973)
);

XNOR2xp5_ASAP7_75t_L g1974 ( 
.A(n_1973),
.B(n_1970),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1974),
.Y(n_1975)
);

AOI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1974),
.A2(n_1972),
.B(n_1968),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1976),
.A2(n_1965),
.B(n_1971),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1975),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1978),
.B(n_1967),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_SL g1980 ( 
.A1(n_1977),
.A2(n_1472),
.B(n_1456),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1980),
.A2(n_1516),
.B(n_1440),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1981),
.Y(n_1982)
);

OAI221xp5_ASAP7_75t_R g1983 ( 
.A1(n_1982),
.A2(n_1979),
.B1(n_1761),
.B2(n_1485),
.C(n_1772),
.Y(n_1983)
);

AOI211xp5_ASAP7_75t_L g1984 ( 
.A1(n_1983),
.A2(n_1440),
.B(n_1405),
.C(n_1519),
.Y(n_1984)
);


endmodule