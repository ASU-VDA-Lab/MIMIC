module real_jpeg_22763_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_216;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_35),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_143)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_25),
.B1(n_33),
.B2(n_36),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_7),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_112)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_8),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_44),
.B1(n_61),
.B2(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_44),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_9),
.B(n_53),
.C(n_66),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_9),
.B(n_67),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_33),
.C(n_49),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_21),
.C(n_39),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_9),
.B(n_42),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_115),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_11),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_119),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_118),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_99),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_16),
.B(n_99),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_72),
.C(n_84),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_17),
.B(n_72),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_18),
.B(n_58),
.C(n_70),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_19),
.A2(n_30),
.B1(n_31),
.B2(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_20),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_20),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_21),
.B(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_23),
.A2(n_78),
.B(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_28),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_30),
.A2(n_31),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_30),
.A2(n_31),
.B1(n_169),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_31),
.B(n_163),
.C(n_169),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_31),
.B(n_141),
.C(n_200),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_33),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_43),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_37),
.A2(n_42),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_37),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_81),
.B(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_41),
.A2(n_82),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_41),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_43),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_46),
.A2(n_70),
.B1(n_130),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_46),
.A2(n_70),
.B1(n_91),
.B2(n_126),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_46),
.B(n_91),
.C(n_207),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_54),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_56)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_51),
.Y(n_53)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_53),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_53),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_57),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_71),
.B1(n_113),
.B2(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_58),
.B(n_113),
.C(n_136),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_129),
.C(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_79),
.B1(n_80),
.B2(n_83),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_83),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_80),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_75),
.B(n_144),
.Y(n_174)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_84),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.C(n_96),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_85),
.A2(n_86),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_87),
.A2(n_91),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_89),
.A2(n_143),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_91),
.A2(n_126),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_91),
.B(n_186),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_93),
.A2(n_96),
.B1(n_129),
.B2(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_93),
.Y(n_226)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_96),
.A2(n_129),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_117),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_113),
.B(n_116),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_113),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_156),
.C(n_158),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_113),
.A2(n_146),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_232),
.B(n_236),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_159),
.B(n_218),
.C(n_231),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_148),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_148),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_135),
.B2(n_147),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_125),
.B(n_134),
.C(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_140),
.A2(n_141),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_192),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_150),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_158),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_217),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_178),
.B(n_216),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_175),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_162),
.B(n_175),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_163),
.A2(n_164),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_209),
.B(n_215),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_203),
.B(n_208),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_195),
.B(n_202),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_187),
.B(n_194),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_191),
.B(n_193),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_197),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_200),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_220),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_230),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_228),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_228),
.C(n_230),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);


endmodule