module fake_jpeg_30750_n_146 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_68),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_1),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_53),
.B(n_58),
.C(n_62),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_55),
.B(n_5),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_51),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_47),
.B1(n_50),
.B2(n_48),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_24),
.B1(n_41),
.B2(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_56),
.Y(n_90)
);

OR2x4_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_47),
.Y(n_85)
);

OR2x4_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_94),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_8),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_1),
.CI(n_3),
.CON(n_92),
.SN(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_9),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_54),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_55),
.B1(n_22),
.B2(n_23),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_102),
.B(n_7),
.Y(n_104)
);

OR2x4_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_4),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_80),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_20),
.B(n_36),
.C(n_35),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_115),
.B(n_16),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_8),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_31),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_119),
.Y(n_122)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_11),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_43),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_17),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_127),
.B1(n_130),
.B2(n_132),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_131),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_18),
.B1(n_19),
.B2(n_26),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_33),
.B1(n_34),
.B2(n_105),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_128),
.C(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_115),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B1(n_131),
.B2(n_110),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_123),
.B(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_108),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_127),
.A3(n_137),
.B1(n_121),
.B2(n_133),
.C1(n_126),
.C2(n_134),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_122),
.C(n_118),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_111),
.Y(n_146)
);


endmodule