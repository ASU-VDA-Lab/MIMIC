module fake_jpeg_28534_n_436 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_436);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_436;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_56),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_58),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_59),
.Y(n_149)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_61),
.A2(n_35),
.B(n_38),
.C(n_41),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_63),
.B(n_80),
.Y(n_121)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_71),
.B(n_79),
.Y(n_151)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_77),
.Y(n_120)
);

INVx11_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_1),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_31),
.B(n_2),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_96),
.Y(n_136)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_15),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_19),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_22),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_47),
.B1(n_26),
.B2(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_101),
.A2(n_103),
.B1(n_113),
.B2(n_122),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_26),
.B1(n_33),
.B2(n_40),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_109),
.B(n_126),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_95),
.B1(n_91),
.B2(n_93),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_58),
.A2(n_2),
.B(n_3),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_51),
.A2(n_26),
.B1(n_33),
.B2(n_40),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_59),
.B(n_52),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_30),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_73),
.B1(n_78),
.B2(n_82),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_131),
.B1(n_141),
.B2(n_118),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_65),
.A2(n_26),
.B1(n_33),
.B2(n_40),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_65),
.A2(n_33),
.B1(n_42),
.B2(n_41),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_55),
.A2(n_35),
.B1(n_42),
.B2(n_38),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_148),
.B1(n_67),
.B2(n_92),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_64),
.A2(n_37),
.B1(n_34),
.B2(n_32),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_37),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_171),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_120),
.B(n_22),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_172),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_163),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g229 ( 
.A1(n_164),
.A2(n_169),
.B(n_173),
.Y(n_229)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

OR2x2_ASAP7_75t_SL g169 ( 
.A(n_124),
.B(n_54),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_198),
.B1(n_149),
.B2(n_119),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_30),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_34),
.C(n_90),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_66),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_116),
.B(n_97),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_181),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_3),
.B(n_4),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_134),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_19),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_183),
.Y(n_233)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_100),
.B(n_87),
.Y(n_185)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_19),
.Y(n_187)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_191),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_110),
.B(n_89),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_196),
.C(n_194),
.Y(n_215)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_123),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_112),
.B(n_53),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_194),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_86),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_199),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_106),
.A2(n_50),
.B1(n_46),
.B2(n_36),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_46),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_143),
.A2(n_46),
.B(n_36),
.C(n_6),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_200),
.A2(n_142),
.B(n_36),
.C(n_46),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_221),
.B(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_169),
.A2(n_122),
.B1(n_103),
.B2(n_141),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_218),
.B1(n_225),
.B2(n_196),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_230),
.B1(n_108),
.B2(n_147),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_129),
.B1(n_131),
.B2(n_115),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_173),
.A2(n_149),
.B(n_144),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_146),
.B1(n_107),
.B2(n_153),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_162),
.A2(n_146),
.B1(n_154),
.B2(n_117),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_162),
.A2(n_106),
.B1(n_117),
.B2(n_115),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_231),
.B(n_235),
.Y(n_240)
);

OAI32xp33_ASAP7_75t_L g232 ( 
.A1(n_159),
.A2(n_142),
.A3(n_154),
.B1(n_123),
.B2(n_36),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_189),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_171),
.B(n_142),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_157),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_147),
.C(n_108),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_238),
.A2(n_229),
.B1(n_215),
.B2(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_242),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_177),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_185),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_255),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_252),
.B1(n_263),
.B2(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_200),
.C(n_189),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_209),
.B(n_231),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_221),
.A2(n_191),
.B1(n_158),
.B2(n_183),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_261),
.B1(n_265),
.B2(n_266),
.Y(n_287)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_180),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_259),
.Y(n_286)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_196),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_190),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_242),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_210),
.A2(n_160),
.B1(n_178),
.B2(n_132),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_184),
.B1(n_168),
.B2(n_195),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_188),
.B(n_186),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_216),
.B(n_223),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_123),
.B1(n_165),
.B2(n_163),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_195),
.B1(n_7),
.B2(n_8),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_224),
.A2(n_195),
.B1(n_167),
.B2(n_46),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_269),
.A2(n_273),
.B(n_264),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_275),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_295),
.B1(n_287),
.B2(n_267),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_223),
.B(n_216),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_235),
.Y(n_275)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_232),
.A3(n_222),
.B1(n_201),
.B2(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_255),
.B(n_201),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_278),
.B(n_262),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_243),
.A2(n_222),
.B(n_211),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_281),
.A2(n_292),
.B(n_254),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_205),
.C(n_233),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_294),
.C(n_259),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_240),
.A2(n_252),
.B1(n_250),
.B2(n_242),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_285),
.A2(n_291),
.B1(n_277),
.B2(n_253),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_256),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_240),
.A2(n_217),
.B1(n_233),
.B2(n_205),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_208),
.B(n_207),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_207),
.C(n_236),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_238),
.A2(n_230),
.B1(n_217),
.B2(n_236),
.Y(n_295)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_301),
.B(n_304),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_308),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_300),
.A2(n_303),
.B1(n_316),
.B2(n_320),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_264),
.B(n_260),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_306),
.B1(n_295),
.B2(n_293),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_287),
.A2(n_263),
.B1(n_266),
.B2(n_265),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_253),
.B(n_266),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_317),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_261),
.B1(n_265),
.B2(n_246),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_311),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_257),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_310),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_282),
.C(n_294),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_275),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_273),
.A2(n_261),
.B(n_241),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_272),
.A2(n_228),
.B1(n_226),
.B2(n_208),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_226),
.B(n_204),
.C(n_220),
.D(n_227),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_228),
.Y(n_318)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_319),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_228),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_322),
.A2(n_325),
.B1(n_326),
.B2(n_333),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_285),
.B1(n_277),
.B2(n_268),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_306),
.A2(n_277),
.B1(n_276),
.B2(n_271),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_331),
.C(n_334),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_281),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_271),
.B1(n_291),
.B2(n_269),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_313),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_291),
.B1(n_269),
.B2(n_270),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_335),
.A2(n_338),
.B1(n_314),
.B2(n_316),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_300),
.A2(n_292),
.B1(n_284),
.B2(n_289),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_282),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_286),
.C(n_318),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_307),
.A2(n_278),
.B(n_274),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_310),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_294),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_297),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_358),
.C(n_360),
.Y(n_370)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_341),
.Y(n_347)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_337),
.Y(n_349)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_332),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_350),
.B(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_308),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_354),
.A2(n_329),
.B1(n_338),
.B2(n_335),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_345),
.A2(n_312),
.B1(n_304),
.B2(n_303),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_356),
.A2(n_366),
.B1(n_336),
.B2(n_317),
.Y(n_374)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_286),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_296),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_301),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_342),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_362),
.A2(n_364),
.B1(n_365),
.B2(n_333),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_310),
.B(n_320),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_363),
.A2(n_227),
.B(n_7),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_284),
.C(n_289),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_319),
.C(n_315),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_327),
.A2(n_311),
.B1(n_309),
.B2(n_317),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_8),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_326),
.B1(n_325),
.B2(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_369),
.B(n_374),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_373),
.A2(n_376),
.B1(n_346),
.B2(n_167),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_331),
.B1(n_336),
.B2(n_343),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_343),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_6),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_366),
.A2(n_220),
.B1(n_167),
.B2(n_36),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_383),
.A2(n_354),
.B1(n_361),
.B2(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_388),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_387),
.A2(n_372),
.B1(n_381),
.B2(n_382),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_358),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_355),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_390),
.B(n_393),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_365),
.B(n_364),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_355),
.C(n_360),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_394),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_8),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_395),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_396),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_374),
.B(n_380),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_397),
.A2(n_407),
.B(n_378),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_396),
.B(n_375),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_403),
.Y(n_416)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_384),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_393),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_405),
.B(n_387),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_372),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_383),
.B1(n_371),
.B2(n_382),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_R g409 ( 
.A(n_404),
.B(n_389),
.Y(n_409)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_409),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_410),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_398),
.A2(n_392),
.B(n_381),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_412),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_400),
.A2(n_397),
.B(n_406),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_414),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_390),
.C(n_389),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_8),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_378),
.B1(n_369),
.B2(n_11),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_417),
.B(n_399),
.C(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_416),
.A2(n_401),
.B(n_10),
.C(n_11),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_420),
.B(n_13),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_417),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_425),
.A2(n_421),
.B1(n_418),
.B2(n_414),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_423),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_426),
.A2(n_422),
.B(n_420),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_13),
.B(n_19),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_430),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g433 ( 
.A(n_431),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_432),
.B(n_427),
.C(n_13),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_434),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_435),
.B(n_433),
.Y(n_436)
);


endmodule