module fake_jpeg_20385_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_30),
.B1(n_16),
.B2(n_27),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_23),
.B1(n_16),
.B2(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_49),
.B(n_21),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_22),
.B1(n_36),
.B2(n_41),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_83),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_40),
.B1(n_39),
.B2(n_41),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_72),
.B1(n_82),
.B2(n_88),
.Y(n_91)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_73),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_35),
.B1(n_38),
.B2(n_31),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_37),
.A3(n_38),
.B1(n_31),
.B2(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_70),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_33),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_77),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_33),
.C(n_18),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_79),
.C(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_56),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_30),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_29),
.C(n_25),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_58),
.B1(n_55),
.B2(n_47),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_95),
.B1(n_101),
.B2(n_103),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_53),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_69),
.B(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_58),
.B1(n_57),
.B2(n_53),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_105),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_57),
.B1(n_28),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_28),
.B1(n_25),
.B2(n_15),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_15),
.B1(n_29),
.B2(n_5),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_108),
.B(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_117),
.B(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_80),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_118),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_98),
.B(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_69),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_129),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_79),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_123),
.C(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_79),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_128),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_88),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_73),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_64),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_130),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_140),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_135),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_102),
.B1(n_89),
.B2(n_97),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_91),
.B1(n_98),
.B2(n_100),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_91),
.B1(n_100),
.B2(n_105),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_103),
.C(n_95),
.Y(n_141)
);

XOR2x2_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_143),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_101),
.C(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_151),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_113),
.A3(n_119),
.B1(n_125),
.B2(n_121),
.C1(n_122),
.C2(n_127),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_127),
.A3(n_129),
.B1(n_12),
.B2(n_14),
.C1(n_10),
.C2(n_13),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_137),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_104),
.B(n_67),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_138),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_132),
.C(n_156),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_135),
.B1(n_141),
.B2(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_155),
.B1(n_150),
.B2(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_157),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_169),
.C(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_146),
.B1(n_131),
.B2(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_158),
.B1(n_164),
.B2(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_159),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_174),
.A3(n_175),
.B1(n_176),
.B2(n_177),
.C1(n_168),
.C2(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_159),
.C(n_162),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_14),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_179),
.B(n_180),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_167),
.B1(n_168),
.B2(n_86),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_12),
.A3(n_75),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_8),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_4),
.B(n_5),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_181),
.B(n_7),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_6),
.B(n_7),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_75),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_7),
.Y(n_187)
);


endmodule