module fake_jpeg_8375_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_32),
.B1(n_25),
.B2(n_27),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_30),
.B(n_35),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_50),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_32),
.B1(n_27),
.B2(n_20),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_21),
.B1(n_18),
.B2(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_26),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_25),
.C(n_30),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_28),
.B1(n_39),
.B2(n_17),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_69),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_28),
.B1(n_39),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_66),
.A2(n_73),
.B1(n_76),
.B2(n_86),
.Y(n_119)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_28),
.B1(n_40),
.B2(n_33),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_85),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_40),
.B1(n_22),
.B2(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_26),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_14),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_88),
.B1(n_23),
.B2(n_38),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_35),
.B1(n_24),
.B2(n_21),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_90),
.B1(n_91),
.B2(n_23),
.Y(n_113)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_60),
.B(n_38),
.CI(n_37),
.CON(n_85),
.SN(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_40),
.B1(n_22),
.B2(n_31),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_92),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_63),
.B1(n_50),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_44),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_93),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_102),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_62),
.B1(n_53),
.B2(n_49),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_105),
.B1(n_120),
.B2(n_121),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_82),
.A2(n_52),
.B(n_29),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_115),
.B(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_49),
.B1(n_61),
.B2(n_41),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_49),
.B1(n_61),
.B2(n_34),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_113),
.B1(n_122),
.B2(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_41),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_118),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_0),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_1),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_11),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_41),
.C(n_38),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_37),
.C(n_34),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_41),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_41),
.B1(n_23),
.B2(n_38),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_1),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_128),
.A2(n_132),
.B1(n_133),
.B2(n_71),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_78),
.B(n_94),
.C(n_83),
.D(n_95),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_119),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_141),
.B(n_155),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_8),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_95),
.B1(n_93),
.B2(n_69),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_88),
.B1(n_70),
.B2(n_89),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_38),
.CI(n_37),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_105),
.A2(n_84),
.B1(n_70),
.B2(n_37),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_106),
.B1(n_123),
.B2(n_34),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_117),
.C(n_122),
.Y(n_156)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_142),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_12),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_37),
.B1(n_34),
.B2(n_59),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_182)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_34),
.B1(n_48),
.B2(n_71),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_103),
.B1(n_120),
.B2(n_108),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_152),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_165),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_108),
.B(n_124),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_166),
.B(n_175),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_180),
.B1(n_182),
.B2(n_185),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_164),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_102),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_119),
.B(n_110),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_178),
.B1(n_143),
.B2(n_149),
.Y(n_204)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_99),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_99),
.B1(n_112),
.B2(n_115),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_115),
.C(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_152),
.B(n_138),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_4),
.B(n_5),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_128),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_136),
.B(n_134),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_192),
.A2(n_206),
.B(n_216),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_126),
.B1(n_134),
.B2(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_196),
.B1(n_204),
.B2(n_209),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_143),
.B1(n_136),
.B2(n_149),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_201),
.B(n_205),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_149),
.B(n_131),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_186),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_208),
.B(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_215),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_177),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_226),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_163),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_222),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_165),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_156),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_231),
.C(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_211),
.A2(n_157),
.B(n_166),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_232),
.B1(n_190),
.B2(n_209),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_240),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_162),
.B(n_164),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_172),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_182),
.B1(n_168),
.B2(n_159),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_195),
.B(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_170),
.B(n_158),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_179),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_176),
.B(n_6),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_213),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_202),
.C(n_194),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_249),
.C(n_227),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_202),
.B1(n_190),
.B2(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_203),
.C(n_206),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_225),
.A2(n_203),
.B1(n_207),
.B2(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_207),
.B1(n_176),
.B2(n_7),
.Y(n_256)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_230),
.B(n_240),
.C(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_239),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_263),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_222),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_266),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_231),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_223),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_244),
.B(n_252),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_274),
.C(n_275),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_223),
.C(n_233),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_225),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_281),
.B(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_255),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_286),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_244),
.B(n_257),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_218),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_250),
.B(n_251),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_246),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_257),
.B(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_242),
.Y(n_293)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_292),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_277),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_276),
.B(n_254),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_278),
.A3(n_237),
.B1(n_283),
.B2(n_266),
.C1(n_11),
.C2(n_12),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_268),
.B1(n_218),
.B2(n_275),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

OAI221xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_256),
.B1(n_279),
.B2(n_278),
.C(n_285),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_299),
.A2(n_301),
.B(n_303),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_5),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_305),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_6),
.B(n_7),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_298),
.C(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_310),
.C(n_311),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_309),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_290),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_300),
.B(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.C(n_309),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_14),
.B1(n_15),
.B2(n_312),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule