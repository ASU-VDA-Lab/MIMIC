module fake_jpeg_1073_n_176 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_58),
.Y(n_71)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_47),
.B1(n_54),
.B2(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_80),
.B1(n_63),
.B2(n_61),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_54),
.B1(n_46),
.B2(n_57),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_46),
.B1(n_45),
.B2(n_49),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_51),
.B1(n_56),
.B2(n_50),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_2),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_94),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_95),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_2),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_75),
.B1(n_63),
.B2(n_73),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_106),
.B1(n_110),
.B2(n_43),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_83),
.C(n_93),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_52),
.C(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_64),
.B1(n_66),
.B2(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_66),
.B1(n_56),
.B2(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_115),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_82),
.B1(n_92),
.B2(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_64),
.B1(n_56),
.B2(n_50),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_120),
.B1(n_129),
.B2(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_48),
.B1(n_53),
.B2(n_52),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_53),
.B1(n_48),
.B2(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_6),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_8),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_21),
.B1(n_41),
.B2(n_38),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_107),
.Y(n_130)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_19),
.B(n_37),
.C(n_35),
.D(n_34),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_129),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_134),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_110),
.B(n_29),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_140),
.Y(n_158)
);

AOI221xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_104),
.B(n_9),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_31),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_117),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_26),
.B(n_23),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_10),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_10),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_149),
.C(n_137),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_147),
.C(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_164),
.C(n_159),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_150),
.C(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_165),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_143),
.B1(n_141),
.B2(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_158),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_143),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_146),
.A3(n_142),
.B1(n_14),
.B2(n_15),
.C1(n_17),
.C2(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_166),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_167),
.B(n_154),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_154),
.C(n_11),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_17),
.Y(n_176)
);


endmodule