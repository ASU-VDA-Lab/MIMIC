module fake_jpeg_30476_n_74 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_37),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_1),
.CI(n_2),
.CON(n_48),
.SN(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_32),
.B(n_28),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_45),
.B(n_6),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_32),
.B(n_28),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_26),
.B1(n_31),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_26),
.B2(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_26),
.B1(n_14),
.B2(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_5),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.C(n_44),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_60)
);

AO21x1_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_2),
.B(n_4),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_11),
.B(n_12),
.Y(n_59)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_57),
.CI(n_21),
.CON(n_65),
.SN(n_65)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_5),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_19),
.B(n_20),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_17),
.C(n_7),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_6),
.B(n_10),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_59),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.C(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_25),
.C(n_62),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.C(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_67),
.Y(n_74)
);


endmodule