module fake_aes_9585_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_2), .B(n_9), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_14), .B(n_0), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
OA21x2_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_13), .B(n_15), .Y(n_20) );
NAND2x1p5_ASAP7_75t_L g21 ( .A(n_17), .B(n_11), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_22), .B1(n_16), .B2(n_20), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
NOR2x1_ASAP7_75t_SL g30 ( .A(n_26), .B(n_22), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_11), .Y(n_31) );
NOR3xp33_ASAP7_75t_L g32 ( .A(n_28), .B(n_17), .C(n_16), .Y(n_32) );
O2A1O1Ixp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_0), .B(n_3), .C(n_4), .Y(n_33) );
INVx4_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_31), .B(n_3), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_33), .B1(n_30), .B2(n_8), .Y(n_36) );
AOI22xp33_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_35), .B1(n_7), .B2(n_10), .Y(n_37) );
endmodule