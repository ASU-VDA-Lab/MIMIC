module fake_jpeg_24587_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_49),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_20),
.B1(n_25),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_29),
.B1(n_33),
.B2(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_58),
.A2(n_38),
.B1(n_28),
.B2(n_17),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_31),
.B1(n_18),
.B2(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_31),
.B1(n_18),
.B2(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_20),
.B1(n_33),
.B2(n_23),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_22),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_76),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_20),
.B1(n_33),
.B2(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_75),
.B1(n_82),
.B2(n_38),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_23),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_22),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_29),
.B1(n_37),
.B2(n_21),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_92),
.B1(n_85),
.B2(n_93),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_21),
.B1(n_27),
.B2(n_22),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_19),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_89),
.Y(n_129)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_27),
.B1(n_39),
.B2(n_19),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_65),
.B(n_39),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_97),
.B(n_111),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_58),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_122),
.B1(n_74),
.B2(n_68),
.Y(n_132)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_113),
.B1(n_125),
.B2(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_105),
.Y(n_158)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_36),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_114),
.B1(n_118),
.B2(n_87),
.Y(n_141)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_59),
.B(n_71),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_32),
.B1(n_30),
.B2(n_38),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_73),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g123 ( 
.A(n_58),
.B(n_32),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_73),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_58),
.A2(n_38),
.B(n_28),
.C(n_17),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_55),
.B(n_84),
.C(n_17),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_88),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_132),
.B1(n_138),
.B2(n_143),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_123),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_131),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_152),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_62),
.B(n_74),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_148),
.C(n_160),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_63),
.B1(n_70),
.B2(n_87),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_142),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_161),
.B1(n_163),
.B2(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_89),
.B1(n_28),
.B2(n_17),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_3),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_102),
.B(n_80),
.CI(n_1),
.CON(n_146),
.SN(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_154),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_80),
.C(n_81),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_124),
.A3(n_112),
.B1(n_115),
.B2(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_98),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_81),
.A3(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_11),
.Y(n_186)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_0),
.Y(n_153)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_99),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_0),
.C(n_1),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_110),
.B(n_1),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_167),
.B1(n_176),
.B2(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_124),
.B1(n_113),
.B2(n_108),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_120),
.C(n_96),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_160),
.C(n_162),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_149),
.A2(n_121),
.B1(n_117),
.B2(n_119),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_110),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_106),
.B1(n_100),
.B2(n_95),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_194),
.B(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_126),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_156),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_186),
.B1(n_146),
.B2(n_134),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_132),
.A2(n_117),
.B1(n_101),
.B2(n_103),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_198),
.B1(n_199),
.B2(n_143),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_104),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_196),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_103),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_4),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_136),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_206),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_207),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_205),
.B1(n_208),
.B2(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_138),
.B1(n_145),
.B2(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_173),
.B(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_211),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_145),
.B(n_146),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_224),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_135),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.C(n_223),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_171),
.C(n_169),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_157),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_137),
.C(n_136),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_165),
.A2(n_137),
.B1(n_161),
.B2(n_163),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_147),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_186),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_172),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_245),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_238),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_194),
.CI(n_203),
.CON(n_267),
.SN(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_250),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_226),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_173),
.B(n_191),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_166),
.C(n_176),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_202),
.C(n_227),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_202),
.A2(n_167),
.B1(n_197),
.B2(n_177),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_205),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_255),
.C(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_218),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_258),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_214),
.C(n_215),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_239),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_195),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_249),
.B(n_211),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_230),
.B1(n_177),
.B2(n_246),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_261),
.B1(n_270),
.B2(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_213),
.C(n_216),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_247),
.B1(n_250),
.B2(n_236),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_221),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_266),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_211),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_199),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_166),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_262),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_201),
.B1(n_178),
.B2(n_168),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_248),
.C(n_243),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_275),
.C(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_242),
.B1(n_231),
.B2(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_282),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_245),
.C(n_241),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_286),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_229),
.B1(n_239),
.B2(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_213),
.C(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_178),
.B(n_168),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_265),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_180),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_184),
.B1(n_182),
.B2(n_198),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_269),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_194),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_287),
.C(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_296),
.C(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_277),
.B(n_147),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_275),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_271),
.C(n_272),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_309),
.C(n_288),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_305),
.B(n_294),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_294),
.A2(n_184),
.B1(n_278),
.B2(n_285),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_271),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_279),
.C(n_286),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_252),
.CI(n_8),
.CON(n_322),
.SN(n_322)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_279),
.C(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_297),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_304),
.A2(n_290),
.B(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_289),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_299),
.B1(n_283),
.B2(n_292),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_252),
.B(n_10),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_311),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_8),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_310),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_321),
.B(n_9),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_8),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_323),
.B(n_321),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_325),
.B(n_9),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_330),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_9),
.Y(n_332)
);


endmodule