module fake_netlist_6_4816_n_248 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_39, n_60, n_59, n_32, n_4, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_31, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_248);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_60;
input n_59;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_31;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_248;

wire n_91;
wire n_119;
wire n_146;
wire n_163;
wire n_235;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_113;
wire n_63;
wire n_223;
wire n_73;
wire n_148;
wire n_199;
wire n_138;
wire n_161;
wire n_208;
wire n_226;
wire n_68;
wire n_228;
wire n_166;
wire n_184;
wire n_212;
wire n_158;
wire n_217;
wire n_210;
wire n_216;
wire n_83;
wire n_206;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_168;
wire n_153;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_189;
wire n_85;
wire n_66;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_213;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_155;
wire n_62;
wire n_219;
wire n_75;
wire n_109;
wire n_150;
wire n_233;
wire n_122;
wire n_205;
wire n_140;
wire n_218;
wire n_70;
wire n_120;
wire n_234;
wire n_214;
wire n_67;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_244;
wire n_181;
wire n_76;
wire n_182;
wire n_124;
wire n_238;
wire n_239;
wire n_126;
wire n_202;
wire n_94;
wire n_108;
wire n_97;
wire n_116;
wire n_211;
wire n_64;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_65;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_200;
wire n_196;
wire n_165;
wire n_139;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_243;
wire n_107;
wire n_71;
wire n_74;
wire n_229;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_201;
wire n_103;
wire n_111;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_69;
wire n_128;
wire n_241;
wire n_79;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_221;

INVx1_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx2_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_6),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_0),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_0),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_4),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_7),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_68),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_72),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_77),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_79),
.C(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_77),
.Y(n_149)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_89),
.Y(n_150)
);

OR2x6_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_96),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_109),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_122),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_116),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_132),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

BUFx4f_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_117),
.Y(n_171)
);

OR2x6_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_157),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_117),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_101),
.C(n_97),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_136),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_139),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_150),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_163),
.Y(n_201)
);

AND2x4_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_161),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_88),
.B1(n_78),
.B2(n_76),
.Y(n_203)
);

CKINVDCx6p67_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_143),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_84),
.B(n_82),
.C(n_156),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_143),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_168),
.Y(n_208)
);

OAI221xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_186),
.B1(n_183),
.B2(n_189),
.C(n_123),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_183),
.B1(n_181),
.B2(n_147),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_197),
.A2(n_174),
.B1(n_176),
.B2(n_180),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g216 ( 
.A(n_200),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_176),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_180),
.B(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

AO21x2_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_206),
.B(n_207),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_196),
.B1(n_204),
.B2(n_159),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

AOI211x1_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_228)
);

AOI221xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_229)
);

OAI33xp33_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_221),
.A3(n_227),
.B1(n_226),
.B2(n_223),
.B3(n_222),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_216),
.Y(n_232)
);

OAI33xp33_ASAP7_75t_L g233 ( 
.A1(n_228),
.A2(n_22),
.A3(n_23),
.B1(n_26),
.B2(n_27),
.B3(n_28),
.Y(n_233)
);

OA211x2_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_29),
.B(n_30),
.C(n_32),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_35),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_235),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_241),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_234),
.B1(n_233),
.B2(n_230),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_47),
.B(n_49),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_60),
.B(n_58),
.Y(n_248)
);


endmodule