module fake_jpeg_15662_n_384 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_384);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_384;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_14),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_1),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_54),
.B(n_25),
.Y(n_111)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_65),
.B(n_82),
.Y(n_143)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx2_ASAP7_75t_SL g146 ( 
.A(n_66),
.Y(n_146)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_40),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_91),
.B1(n_102),
.B2(n_33),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_38),
.A2(n_17),
.B1(n_23),
.B2(n_31),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_106),
.B1(n_63),
.B2(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_23),
.B1(n_34),
.B2(n_29),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_85),
.B1(n_94),
.B2(n_107),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_44),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_101),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_21),
.B1(n_18),
.B2(n_36),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_99),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_29),
.B1(n_19),
.B2(n_31),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_21),
.B1(n_15),
.B2(n_3),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_21),
.B1(n_25),
.B2(n_33),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_32),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_108),
.B(n_13),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_32),
.C(n_26),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_33),
.C(n_3),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_124),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_141),
.B1(n_144),
.B2(n_87),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_66),
.A2(n_52),
.B1(n_32),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_117),
.A2(n_150),
.B1(n_159),
.B2(n_113),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_129),
.Y(n_166)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_98),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_137),
.B1(n_100),
.B2(n_97),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_73),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_127),
.B(n_131),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_149),
.B1(n_69),
.B2(n_70),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_59),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_32),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_142),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_73),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_73),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_133),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_32),
.B(n_33),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_134),
.B(n_138),
.C(n_135),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_1),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_165),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_85),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_75),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_78),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_145),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_154),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_7),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_68),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_74),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_105),
.B1(n_110),
.B2(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_83),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_84),
.A2(n_12),
.B1(n_13),
.B2(n_114),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_167),
.Y(n_247)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_169),
.B(n_181),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_170),
.B(n_175),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_190),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_119),
.B(n_88),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_207),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_204),
.B(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_200),
.B1(n_202),
.B2(n_206),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_203),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_69),
.B1(n_70),
.B2(n_105),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_192),
.A2(n_194),
.B1(n_197),
.B2(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_129),
.B(n_110),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_196),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_126),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_139),
.B1(n_158),
.B2(n_130),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_132),
.C(n_140),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_139),
.A2(n_157),
.B1(n_136),
.B2(n_121),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_135),
.A2(n_148),
.B1(n_156),
.B2(n_121),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_143),
.A2(n_148),
.B1(n_146),
.B2(n_122),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_134),
.B(n_137),
.Y(n_204)
);

OR2x2_ASAP7_75t_SL g205 ( 
.A(n_137),
.B(n_143),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_115),
.A2(n_124),
.B1(n_120),
.B2(n_163),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_140),
.A2(n_133),
.B1(n_127),
.B2(n_131),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_211),
.A2(n_145),
.B1(n_118),
.B2(n_153),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_214),
.B(n_218),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_215),
.B(n_235),
.C(n_229),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_145),
.B(n_153),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_216),
.A2(n_220),
.B(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_161),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_204),
.B(n_210),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_231),
.B1(n_235),
.B2(n_252),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_118),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_166),
.B(n_175),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_166),
.B(n_205),
.C(n_199),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_178),
.B1(n_191),
.B2(n_194),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_202),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_239),
.Y(n_268)
);

AO21x2_ASAP7_75t_L g237 ( 
.A1(n_169),
.A2(n_211),
.B(n_178),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_237),
.A2(n_223),
.B1(n_219),
.B2(n_213),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_188),
.B(n_170),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_174),
.B(n_185),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_243),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_242),
.B(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_189),
.Y(n_243)
);

NAND2x1_ASAP7_75t_SL g244 ( 
.A(n_173),
.B(n_209),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_249),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_179),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_246),
.B(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_181),
.B(n_182),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_230),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_183),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_176),
.B1(n_247),
.B2(n_236),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_274),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_239),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_176),
.B(n_216),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_255),
.A2(n_262),
.B(n_264),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_176),
.B1(n_238),
.B2(n_241),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_272),
.C(n_282),
.Y(n_307)
);

A2O1A1O1Ixp25_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_241),
.B(n_237),
.C(n_227),
.D(n_222),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_240),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_242),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_215),
.B(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_226),
.B1(n_221),
.B2(n_248),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_224),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_284),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_214),
.B(n_213),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_260),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_245),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_232),
.B1(n_246),
.B2(n_253),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_219),
.B(n_212),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_287),
.A2(n_290),
.B(n_291),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_223),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_289),
.C(n_310),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_222),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_256),
.A2(n_212),
.B(n_228),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

XOR2x1_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_295),
.B(n_301),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_255),
.A2(n_264),
.B(n_257),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_297),
.A2(n_298),
.B(n_299),
.Y(n_332)
);

XNOR2x2_ASAP7_75t_SL g298 ( 
.A(n_261),
.B(n_268),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_280),
.B(n_279),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_311),
.Y(n_320)
);

XOR2x2_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_276),
.B(n_266),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_276),
.B1(n_281),
.B2(n_277),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_270),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_267),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_266),
.B(n_279),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_277),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_269),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_313),
.B(n_293),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_291),
.B1(n_325),
.B2(n_318),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_288),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_309),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_331),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_306),
.A2(n_301),
.B1(n_291),
.B2(n_295),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_324),
.A2(n_334),
.B1(n_287),
.B2(n_297),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_301),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_286),
.B(n_299),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_304),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_326),
.B(n_328),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_329),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_303),
.B(n_302),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_307),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_307),
.C(n_289),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_306),
.A2(n_292),
.B1(n_308),
.B2(n_304),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_335),
.A2(n_321),
.B1(n_332),
.B2(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_341),
.B(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_344),
.A2(n_345),
.B1(n_346),
.B2(n_350),
.Y(n_356)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_324),
.A2(n_296),
.B(n_312),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_348),
.B(n_349),
.C(n_351),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_296),
.C(n_294),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_325),
.A2(n_298),
.B1(n_318),
.B2(n_322),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_298),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_337),
.A2(n_322),
.B1(n_330),
.B2(n_327),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_354),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_SL g354 ( 
.A1(n_345),
.A2(n_332),
.B(n_326),
.C(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_349),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_348),
.C(n_351),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_340),
.A2(n_317),
.B1(n_315),
.B2(n_319),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_363),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_350),
.A2(n_315),
.B1(n_336),
.B2(n_335),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_369),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_362),
.A2(n_347),
.B(n_339),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_362),
.B(n_354),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_338),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_359),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_357),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_372),
.A2(n_346),
.B(n_354),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_373),
.B(n_374),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_343),
.B1(n_360),
.B2(n_358),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_365),
.B(n_367),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_375),
.A2(n_354),
.B(n_357),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_356),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_379),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_380),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_381),
.A2(n_376),
.B(n_366),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_352),
.C(n_341),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_352),
.Y(n_384)
);


endmodule