module real_aes_7667_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_746;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_753;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_1), .A2(n_140), .B(n_144), .C(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_2), .A2(n_174), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g516 ( .A(n_3), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_4), .B(n_241), .Y(n_260) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_5), .A2(n_174), .B(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g215 ( .A(n_7), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_8), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_8), .B(n_42), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_9), .A2(n_173), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_10), .B(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g486 ( .A(n_11), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_12), .B(n_255), .Y(n_540) );
INVx1_ASAP7_75t_L g160 ( .A(n_13), .Y(n_160) );
INVx1_ASAP7_75t_L g552 ( .A(n_14), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_15), .A2(n_150), .B(n_237), .C(n_239), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_16), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_17), .B(n_504), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_18), .B(n_174), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_19), .B(n_186), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_20), .A2(n_255), .B(n_270), .C(n_272), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_21), .B(n_241), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_22), .B(n_152), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_23), .A2(n_182), .B(n_239), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_24), .B(n_152), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_25), .Y(n_191) );
INVx1_ASAP7_75t_L g148 ( .A(n_26), .Y(n_148) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_28), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_29), .B(n_152), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_30), .A2(n_31), .B1(n_750), .B2(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_30), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_31), .Y(n_750) );
INVx1_ASAP7_75t_L g180 ( .A(n_32), .Y(n_180) );
INVx1_ASAP7_75t_L g495 ( .A(n_33), .Y(n_495) );
INVx2_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_35), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_36), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
INVxp67_ASAP7_75t_L g181 ( .A(n_37), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_38), .A2(n_144), .B(n_147), .C(n_155), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_39), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_40), .A2(n_140), .B(n_144), .C(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_41), .A2(n_105), .B1(n_115), .B2(n_757), .Y(n_104) );
INVx1_ASAP7_75t_L g114 ( .A(n_42), .Y(n_114) );
INVx1_ASAP7_75t_L g494 ( .A(n_43), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_44), .A2(n_199), .B(n_213), .C(n_214), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_45), .B(n_152), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_46), .A2(n_747), .B1(n_753), .B2(n_754), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_46), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_47), .A2(n_748), .B1(n_749), .B2(n_752), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_47), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_48), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_49), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_50), .B(n_456), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_51), .A2(n_460), .B1(n_466), .B2(n_755), .Y(n_465) );
INVx1_ASAP7_75t_L g268 ( .A(n_52), .Y(n_268) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_53), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_54), .B(n_174), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_55), .A2(n_144), .B1(n_272), .B2(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_56), .A2(n_71), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_56), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_57), .Y(n_513) );
CKINVDCx14_ASAP7_75t_R g211 ( .A(n_58), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_59), .A2(n_213), .B(n_258), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_60), .Y(n_568) );
INVx1_ASAP7_75t_L g483 ( .A(n_61), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_62), .A2(n_91), .B1(n_454), .B2(n_455), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_62), .Y(n_455) );
INVx1_ASAP7_75t_L g141 ( .A(n_63), .Y(n_141) );
INVx1_ASAP7_75t_L g159 ( .A(n_64), .Y(n_159) );
INVx1_ASAP7_75t_SL g257 ( .A(n_65), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_67), .B(n_241), .Y(n_274) );
INVx1_ASAP7_75t_L g194 ( .A(n_68), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_SL g503 ( .A1(n_69), .A2(n_258), .B(n_504), .C(n_505), .Y(n_503) );
INVxp67_ASAP7_75t_L g506 ( .A(n_70), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_71), .Y(n_125) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_73), .A2(n_174), .B(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_74), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_75), .A2(n_174), .B(n_234), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_76), .Y(n_498) );
INVx1_ASAP7_75t_L g562 ( .A(n_77), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_78), .A2(n_173), .B(n_175), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_79), .Y(n_142) );
INVx1_ASAP7_75t_L g235 ( .A(n_80), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_81), .A2(n_140), .B(n_144), .C(n_564), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_82), .A2(n_174), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g238 ( .A(n_83), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_84), .B(n_149), .Y(n_529) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
INVx1_ASAP7_75t_L g226 ( .A(n_86), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_87), .B(n_504), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_88), .A2(n_140), .B(n_144), .C(n_515), .Y(n_514) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_89), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g459 ( .A(n_89), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g469 ( .A(n_89), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_90), .A2(n_144), .B(n_193), .C(n_201), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_91), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_92), .B(n_156), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_93), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_94), .A2(n_140), .B(n_144), .C(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_95), .Y(n_544) );
INVx1_ASAP7_75t_L g502 ( .A(n_96), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_97), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_98), .B(n_149), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_99), .B(n_164), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_100), .B(n_164), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g271 ( .A(n_102), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_103), .A2(n_174), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_SL g758 ( .A(n_105), .Y(n_758) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g461 ( .A(n_108), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AO21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_464), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g756 ( .A(n_118), .Y(n_756) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_456), .B(n_463), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_127), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_SL g531 ( .A(n_124), .B(n_163), .Y(n_531) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
XOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_453), .Y(n_127) );
INVx2_ASAP7_75t_L g470 ( .A(n_128), .Y(n_470) );
OR4x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_343), .C(n_390), .D(n_430), .Y(n_128) );
NAND3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_289), .C(n_318), .Y(n_129) );
AOI211xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_204), .B(n_242), .C(n_282), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_131), .A2(n_302), .B(n_319), .C(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_166), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_133), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_SL g285 ( .A(n_133), .Y(n_285) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_133), .Y(n_297) );
AND2x4_ASAP7_75t_L g301 ( .A(n_133), .B(n_249), .Y(n_301) );
AND2x2_ASAP7_75t_L g312 ( .A(n_133), .B(n_189), .Y(n_312) );
OR2x2_ASAP7_75t_L g336 ( .A(n_133), .B(n_245), .Y(n_336) );
AND2x2_ASAP7_75t_L g349 ( .A(n_133), .B(n_250), .Y(n_349) );
AND2x2_ASAP7_75t_L g389 ( .A(n_133), .B(n_375), .Y(n_389) );
AND2x2_ASAP7_75t_L g396 ( .A(n_133), .B(n_359), .Y(n_396) );
AND2x2_ASAP7_75t_L g426 ( .A(n_133), .B(n_167), .Y(n_426) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_161), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_143), .C(n_156), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_135), .A2(n_191), .B(n_192), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_135), .A2(n_223), .B(n_224), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_135), .A2(n_184), .B1(n_492), .B2(n_496), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_135), .A2(n_513), .B(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g561 ( .A1(n_135), .A2(n_562), .B(n_563), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g174 ( .A(n_136), .B(n_140), .Y(n_174) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g273 ( .A(n_138), .Y(n_273) );
INVx1_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
INVx1_ASAP7_75t_L g504 ( .A(n_139), .Y(n_504) );
BUFx3_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
INVx4_ASAP7_75t_SL g184 ( .A(n_140), .Y(n_184) );
INVx5_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g200 ( .A(n_145), .Y(n_200) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_145), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_151), .C(n_153), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g179 ( .A1(n_149), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_149), .A2(n_516), .B(n_517), .C(n_518), .Y(n_515) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_150), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_150), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_150), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
INVx4_ASAP7_75t_L g255 ( .A(n_152), .Y(n_255) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_154), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_156), .A2(n_209), .B(n_216), .Y(n_208) );
INVx1_ASAP7_75t_L g221 ( .A(n_156), .Y(n_221) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_156), .A2(n_547), .B(n_553), .Y(n_546) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_157), .B(n_158), .Y(n_156) );
AND2x2_ASAP7_75t_L g165 ( .A(n_157), .B(n_158), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_163), .A2(n_190), .B(n_202), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_163), .B(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_164), .A2(n_500), .B(n_507), .Y(n_499) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_166), .B(n_353), .Y(n_365) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_188), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_167), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g303 ( .A(n_167), .B(n_188), .Y(n_303) );
BUFx3_ASAP7_75t_L g311 ( .A(n_167), .Y(n_311) );
OR2x2_ASAP7_75t_L g332 ( .A(n_167), .B(n_207), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_167), .B(n_353), .Y(n_443) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_172), .B(n_185), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_169), .A2(n_246), .B(n_247), .Y(n_245) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_169), .A2(n_561), .B(n_567), .Y(n_560) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_SL g525 ( .A1(n_170), .A2(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_171), .A2(n_491), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_171), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_171), .A2(n_512), .B(n_519), .Y(n_511) );
INVx1_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_184), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g210 ( .A1(n_177), .A2(n_184), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_177), .A2(n_184), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_177), .A2(n_184), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g267 ( .A1(n_177), .A2(n_184), .B(n_268), .C(n_269), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_177), .A2(n_184), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_177), .A2(n_184), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_177), .A2(n_184), .B(n_549), .C(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_182), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_182), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_182), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_183), .A2(n_196), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
INVx1_ASAP7_75t_L g247 ( .A(n_185), .Y(n_247) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_187), .B(n_203), .Y(n_202) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_187), .A2(n_536), .B(n_543), .Y(n_535) );
AND2x2_ASAP7_75t_L g248 ( .A(n_188), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
AND2x2_ASAP7_75t_L g359 ( .A(n_188), .B(n_250), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_188), .A2(n_362), .B1(n_364), .B2(n_366), .C(n_367), .Y(n_361) );
AND2x2_ASAP7_75t_L g375 ( .A(n_188), .B(n_245), .Y(n_375) );
AND2x2_ASAP7_75t_L g401 ( .A(n_188), .B(n_285), .Y(n_401) );
INVx2_ASAP7_75t_SL g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g281 ( .A(n_189), .B(n_250), .Y(n_281) );
BUFx2_ASAP7_75t_L g415 ( .A(n_189), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_197), .C(n_198), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_L g225 ( .A1(n_195), .A2(n_198), .B(n_226), .C(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_198), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_198), .A2(n_565), .B(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_205), .A2(n_342), .A3(n_356), .B1(n_382), .B2(n_383), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_217), .Y(n_205) );
AND2x2_ASAP7_75t_L g322 ( .A(n_206), .B(n_264), .Y(n_322) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g304 ( .A(n_207), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_207), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g376 ( .A(n_207), .B(n_264), .Y(n_376) );
AND2x2_ASAP7_75t_L g387 ( .A(n_207), .B(n_279), .Y(n_387) );
BUFx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g288 ( .A(n_208), .B(n_265), .Y(n_288) );
AND2x2_ASAP7_75t_L g292 ( .A(n_208), .B(n_265), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_208), .B(n_278), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_208), .B(n_230), .Y(n_334) );
OAI211xp5_ASAP7_75t_L g339 ( .A1(n_208), .A2(n_285), .B(n_296), .C(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g393 ( .A(n_208), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_208), .B(n_219), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_217), .B(n_276), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_217), .B(n_292), .Y(n_382) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g287 ( .A(n_218), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
AND2x2_ASAP7_75t_L g279 ( .A(n_219), .B(n_231), .Y(n_279) );
OR2x2_ASAP7_75t_L g294 ( .A(n_219), .B(n_231), .Y(n_294) );
AND2x2_ASAP7_75t_L g317 ( .A(n_219), .B(n_278), .Y(n_317) );
INVx1_ASAP7_75t_L g321 ( .A(n_219), .Y(n_321) );
AND2x2_ASAP7_75t_L g340 ( .A(n_219), .B(n_277), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_219), .A2(n_305), .B1(n_351), .B2(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_219), .B(n_393), .Y(n_417) );
AND2x2_ASAP7_75t_L g432 ( .A(n_219), .B(n_292), .Y(n_432) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx3_ASAP7_75t_L g262 ( .A(n_220), .Y(n_262) );
AND2x2_ASAP7_75t_L g306 ( .A(n_220), .B(n_231), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_220), .B(n_264), .Y(n_308) );
AND3x2_ASAP7_75t_L g370 ( .A(n_220), .B(n_334), .C(n_371), .Y(n_370) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_228), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_221), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_221), .B(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_221), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g405 ( .A(n_230), .B(n_277), .Y(n_405) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g264 ( .A(n_231), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_231), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_231), .B(n_276), .Y(n_338) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_231), .B(n_317), .C(n_393), .Y(n_445) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_240), .Y(n_231) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_251), .B(n_260), .Y(n_250) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_266), .B(n_274), .Y(n_265) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_241), .A2(n_481), .B(n_487), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_261), .B1(n_275), .B2(n_280), .Y(n_242) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_248), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_245), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g357 ( .A(n_245), .Y(n_357) );
OAI31xp33_ASAP7_75t_L g373 ( .A1(n_248), .A2(n_374), .A3(n_375), .B(n_376), .Y(n_373) );
AND2x2_ASAP7_75t_L g398 ( .A(n_248), .B(n_285), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_248), .B(n_311), .Y(n_444) );
AND2x2_ASAP7_75t_L g353 ( .A(n_249), .B(n_285), .Y(n_353) );
AND2x2_ASAP7_75t_L g414 ( .A(n_249), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g284 ( .A(n_250), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g342 ( .A(n_250), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_259), .Y(n_541) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_262), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_263), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AOI221x1_ASAP7_75t_SL g330 ( .A1(n_264), .A2(n_331), .B1(n_333), .B2(n_335), .C(n_337), .Y(n_330) );
INVx2_ASAP7_75t_L g278 ( .A(n_265), .Y(n_278) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_265), .Y(n_372) );
INVx2_ASAP7_75t_L g518 ( .A(n_272), .Y(n_518) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g360 ( .A(n_275), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_276), .B(n_293), .Y(n_385) );
INVx1_ASAP7_75t_SL g448 ( .A(n_276), .Y(n_448) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g366 ( .A(n_279), .B(n_292), .Y(n_366) );
INVx1_ASAP7_75t_L g434 ( .A(n_280), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_280), .B(n_363), .Y(n_447) );
INVx2_ASAP7_75t_SL g286 ( .A(n_281), .Y(n_286) );
AND2x2_ASAP7_75t_L g329 ( .A(n_281), .B(n_285), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_281), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_281), .B(n_356), .Y(n_383) );
AOI21xp33_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_286), .B(n_287), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_284), .B(n_356), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_284), .B(n_311), .Y(n_452) );
OR2x2_ASAP7_75t_L g324 ( .A(n_285), .B(n_303), .Y(n_324) );
AND2x2_ASAP7_75t_L g423 ( .A(n_285), .B(n_414), .Y(n_423) );
OAI22xp5_ASAP7_75t_SL g298 ( .A1(n_286), .A2(n_299), .B1(n_304), .B2(n_307), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_286), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g346 ( .A(n_288), .B(n_294), .Y(n_346) );
INVx1_ASAP7_75t_L g410 ( .A(n_288), .Y(n_410) );
AOI311xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_295), .A3(n_297), .B(n_298), .C(n_309), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_293), .A2(n_425), .B1(n_437), .B2(n_440), .C(n_442), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_293), .B(n_448), .Y(n_450) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g347 ( .A(n_295), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_338), .B(n_339), .C(n_341), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
O2A1O1Ixp33_ASAP7_75t_SL g406 ( .A1(n_300), .A2(n_302), .B(n_407), .C(n_408), .Y(n_406) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_301), .B(n_375), .Y(n_441) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_304), .A2(n_324), .B1(n_325), .B2(n_328), .C(n_330), .Y(n_323) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g409 ( .A(n_306), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_310), .A2(n_368), .B(n_369), .C(n_373), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_311), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_311), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_321), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g435 ( .A(n_324), .Y(n_435) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_327), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g362 ( .A(n_327), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g439 ( .A(n_327), .Y(n_439) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g380 ( .A(n_329), .B(n_356), .Y(n_380) );
INVx1_ASAP7_75t_SL g374 ( .A(n_336), .Y(n_374) );
INVx1_ASAP7_75t_L g351 ( .A(n_342), .Y(n_351) );
NAND3xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_361), .C(n_377), .Y(n_343) );
AOI322xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .A3(n_348), .B1(n_350), .B2(n_354), .C1(n_358), .C2(n_360), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_345), .A2(n_398), .B(n_399), .C(n_406), .Y(n_397) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_348), .A2(n_369), .B1(n_400), .B2(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g358 ( .A(n_356), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g395 ( .A(n_356), .B(n_396), .Y(n_395) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_356), .A2(n_447), .A3(n_448), .B1(n_449), .B2(n_451), .Y(n_446) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g368 ( .A(n_359), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_359), .A2(n_412), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_411) );
AND2x2_ASAP7_75t_L g425 ( .A(n_359), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g428 ( .A(n_363), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g438 ( .A(n_363), .B(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g429 ( .A(n_372), .B(n_393), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_381), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_394), .B(n_397), .C(n_411), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_405), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g420 ( .A(n_417), .Y(n_420) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B(n_427), .Y(n_421) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_433), .B(n_436), .C(n_446), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NOR2x2_ASAP7_75t_L g755 ( .A(n_460), .B(n_469), .Y(n_755) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_463), .A2(n_465), .B(n_756), .Y(n_464) );
XNOR2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_746), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_471), .B2(n_473), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_469), .Y(n_472) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND3x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_668), .C(n_713), .Y(n_475) );
NOR4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_591), .C(n_632), .D(n_649), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_508), .B(n_522), .C(n_554), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_479), .B(n_509), .Y(n_508) );
NOR4xp25_ASAP7_75t_L g615 ( .A(n_479), .B(n_609), .C(n_616), .D(n_622), .Y(n_615) );
AND2x2_ASAP7_75t_L g688 ( .A(n_479), .B(n_577), .Y(n_688) );
AND2x2_ASAP7_75t_L g707 ( .A(n_479), .B(n_653), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_479), .B(n_702), .Y(n_716) );
AND2x2_ASAP7_75t_L g729 ( .A(n_479), .B(n_521), .Y(n_729) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g574 ( .A(n_480), .Y(n_574) );
AND2x2_ASAP7_75t_L g581 ( .A(n_480), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g631 ( .A(n_480), .B(n_489), .Y(n_631) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_480), .B(n_577), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_480), .B(n_489), .Y(n_646) );
AND2x2_ASAP7_75t_L g655 ( .A(n_480), .B(n_580), .Y(n_655) );
BUFx2_ASAP7_75t_L g678 ( .A(n_480), .Y(n_678) );
AND2x2_ASAP7_75t_L g682 ( .A(n_480), .B(n_499), .Y(n_682) );
OR2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_499), .Y(n_488) );
AND2x2_ASAP7_75t_L g521 ( .A(n_489), .B(n_499), .Y(n_521) );
BUFx2_ASAP7_75t_L g584 ( .A(n_489), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_489), .A2(n_617), .B1(n_619), .B2(n_620), .Y(n_616) );
OR2x2_ASAP7_75t_L g638 ( .A(n_489), .B(n_511), .Y(n_638) );
AND2x2_ASAP7_75t_L g702 ( .A(n_489), .B(n_580), .Y(n_702) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g570 ( .A(n_490), .B(n_511), .Y(n_570) );
AND2x2_ASAP7_75t_L g577 ( .A(n_490), .B(n_499), .Y(n_577) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_490), .Y(n_619) );
OR2x2_ASAP7_75t_L g654 ( .A(n_490), .B(n_510), .Y(n_654) );
INVx1_ASAP7_75t_L g573 ( .A(n_499), .Y(n_573) );
INVx3_ASAP7_75t_L g582 ( .A(n_499), .Y(n_582) );
BUFx2_ASAP7_75t_L g606 ( .A(n_499), .Y(n_606) );
AND2x2_ASAP7_75t_L g639 ( .A(n_499), .B(n_574), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_508), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_510), .B(n_582), .Y(n_586) );
INVx1_ASAP7_75t_L g614 ( .A(n_510), .Y(n_614) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g580 ( .A(n_511), .Y(n_580) );
INVx1_ASAP7_75t_L g592 ( .A(n_521), .Y(n_592) );
NAND2x1_ASAP7_75t_SL g522 ( .A(n_523), .B(n_532), .Y(n_522) );
AND2x2_ASAP7_75t_L g590 ( .A(n_523), .B(n_545), .Y(n_590) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_523), .Y(n_664) );
AND2x2_ASAP7_75t_L g691 ( .A(n_523), .B(n_611), .Y(n_691) );
AND2x2_ASAP7_75t_L g699 ( .A(n_523), .B(n_661), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_523), .B(n_557), .Y(n_726) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g558 ( .A(n_524), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g575 ( .A(n_524), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g596 ( .A(n_524), .Y(n_596) );
INVx1_ASAP7_75t_L g602 ( .A(n_524), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_524), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g635 ( .A(n_524), .B(n_560), .Y(n_635) );
OR2x2_ASAP7_75t_L g673 ( .A(n_524), .B(n_628), .Y(n_673) );
AOI32xp33_ASAP7_75t_L g685 ( .A1(n_524), .A2(n_686), .A3(n_689), .B1(n_690), .B2(n_691), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_524), .B(n_661), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_524), .B(n_621), .Y(n_736) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OR2x2_ASAP7_75t_L g647 ( .A(n_533), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_545), .Y(n_533) );
INVx1_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
AND2x2_ASAP7_75t_L g611 ( .A(n_534), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_534), .B(n_559), .Y(n_628) );
AND2x2_ASAP7_75t_L g661 ( .A(n_534), .B(n_637), .Y(n_661) );
AND2x2_ASAP7_75t_L g698 ( .A(n_534), .B(n_560), .Y(n_698) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g557 ( .A(n_535), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_535), .B(n_559), .Y(n_588) );
AND2x2_ASAP7_75t_L g595 ( .A(n_535), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g636 ( .A(n_535), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_542), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_541), .Y(n_538) );
INVx2_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_545), .B(n_559), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_545), .B(n_603), .Y(n_684) );
INVx1_ASAP7_75t_L g706 ( .A(n_545), .Y(n_706) );
INVx1_ASAP7_75t_L g723 ( .A(n_545), .Y(n_723) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g576 ( .A(n_546), .B(n_559), .Y(n_576) );
AND2x2_ASAP7_75t_L g598 ( .A(n_546), .B(n_560), .Y(n_598) );
INVx1_ASAP7_75t_L g637 ( .A(n_546), .Y(n_637) );
AOI221x1_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_569), .B1(n_575), .B2(n_577), .C(n_578), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_555), .A2(n_642), .B1(n_709), .B2(n_710), .Y(n_708) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g695 ( .A(n_556), .B(n_575), .Y(n_695) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g651 ( .A(n_557), .B(n_576), .Y(n_651) );
INVx1_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
AND2x2_ASAP7_75t_L g674 ( .A(n_558), .B(n_661), .Y(n_674) );
AND2x2_ASAP7_75t_L g741 ( .A(n_558), .B(n_636), .Y(n_741) );
INVx2_ASAP7_75t_L g603 ( .A(n_559), .Y(n_603) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_570), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g693 ( .A(n_570), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_571), .B(n_654), .Y(n_657) );
INVx3_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_572), .A2(n_693), .B(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_575), .B(n_601), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_576), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g667 ( .A(n_576), .B(n_595), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_576), .B(n_602), .Y(n_744) );
AND2x2_ASAP7_75t_L g613 ( .A(n_577), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g680 ( .A(n_577), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .B(n_587), .Y(n_578) );
NAND2x1_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g629 ( .A(n_580), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g641 ( .A(n_580), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_580), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g665 ( .A(n_581), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_581), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_581), .B(n_584), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_584), .A2(n_623), .B(n_653), .C(n_655), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_584), .A2(n_671), .B1(n_674), .B2(n_675), .C(n_679), .Y(n_670) );
AND2x2_ASAP7_75t_L g666 ( .A(n_585), .B(n_619), .Y(n_666) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g626 ( .A(n_590), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g697 ( .A(n_590), .B(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_599), .C(n_624), .Y(n_591) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_592), .B(n_711), .C(n_712), .Y(n_710) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
OR2x2_ASAP7_75t_L g683 ( .A(n_594), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_604), .B1(n_607), .B2(n_613), .C(n_615), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_601), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_601), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g623 ( .A(n_606), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_606), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
OR2x2_ASAP7_75t_L g743 ( .A(n_606), .B(n_654), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVxp67_ASAP7_75t_L g717 ( .A(n_609), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_611), .B(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g618 ( .A(n_612), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_614), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_614), .B(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_614), .B(n_681), .Y(n_720) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_618), .Y(n_644) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g734 ( .A(n_623), .B(n_654), .Y(n_734) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g712 ( .A(n_629), .Y(n_712) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI322xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_638), .A3(n_639), .B1(n_640), .B2(n_643), .C1(n_645), .C2(n_647), .Y(n_632) );
OAI322xp33_ASAP7_75t_L g714 ( .A1(n_633), .A2(n_715), .A3(n_716), .B1(n_717), .B2(n_718), .C1(n_719), .C2(n_721), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx4_ASAP7_75t_L g648 ( .A(n_635), .Y(n_648) );
AND2x2_ASAP7_75t_L g709 ( .A(n_635), .B(n_661), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_635), .B(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g733 ( .A(n_638), .Y(n_733) );
INVx1_ASAP7_75t_L g711 ( .A(n_639), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_641), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g728 ( .A(n_641), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_641), .B(n_682), .Y(n_739) );
OR2x2_ASAP7_75t_L g672 ( .A(n_644), .B(n_673), .Y(n_672) );
INVxp33_ASAP7_75t_L g689 ( .A(n_644), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_648), .A2(n_650), .B1(n_652), .B2(n_656), .C(n_658), .Y(n_649) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_648), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g732 ( .A(n_648), .Y(n_732) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx3_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g696 ( .A1(n_655), .A2(n_680), .A3(n_697), .B1(n_699), .B2(n_700), .C1(n_703), .C2(n_707), .Y(n_696) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_666), .B2(n_667), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_692), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_670), .B(n_685), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_673), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
NAND2xp33_ASAP7_75t_SL g690 ( .A(n_676), .B(n_687), .Y(n_690) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g730 ( .A1(n_678), .A2(n_731), .A3(n_733), .B1(n_734), .B2(n_735), .C1(n_737), .C2(n_740), .Y(n_730) );
AOI21xp33_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B(n_683), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_688), .B(n_736), .Y(n_745) );
OAI211xp5_ASAP7_75t_SL g692 ( .A1(n_693), .A2(n_694), .B(n_696), .C(n_708), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_724), .C(n_730), .D(n_742), .Y(n_713) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
CKINVDCx14_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_744), .B(n_745), .Y(n_742) );
CKINVDCx16_ASAP7_75t_R g754 ( .A(n_747), .Y(n_754) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx4f_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
endmodule