module fake_netlist_6_269_n_1464 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_152, n_92, n_105, n_227, n_132, n_102, n_204, n_261, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_231, n_40, n_240, n_139, n_41, n_134, n_273, n_95, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1464);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_152;
input n_92;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_231;
input n_40;
input n_240;
input n_139;
input n_41;
input n_134;
input n_273;
input n_95;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1464;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1372;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_79),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_245),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_32),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_58),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_159),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_9),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_108),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_204),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_72),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_150),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_127),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_186),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_75),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_172),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_123),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_15),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_23),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_252),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_139),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_25),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_236),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_93),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_210),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_87),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_113),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_116),
.Y(n_341)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_66),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_269),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_228),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_85),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_83),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_165),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_271),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_134),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_191),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_188),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_16),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_100),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_254),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_265),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_187),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_132),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_142),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_225),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_171),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_130),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_138),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_200),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_202),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_61),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_160),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_152),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_42),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_154),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_182),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_282),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_125),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_11),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_161),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_25),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_229),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_148),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_305),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_192),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_69),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_50),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_86),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_216),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_19),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_308),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_215),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_4),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_151),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_153),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_164),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_89),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_101),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_207),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_99),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_48),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_298),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_299),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_218),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_149),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_174),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_179),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_30),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_183),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_67),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_169),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_41),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_250),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_175),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_255),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_277),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_214),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_221),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_205),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_5),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_264),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_280),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_208),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_212),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_95),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_96),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_240),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_71),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_78),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_170),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_15),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_56),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_251),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_31),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_62),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_147),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_119),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_211),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_167),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_62),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_122),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_263),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_233),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_181),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_67),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_176),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_80),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_79),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_2),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_0),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_128),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_87),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_75),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_219),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_166),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_10),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_77),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_129),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_302),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_309),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_198),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_55),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_74),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_266),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_19),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_78),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_117),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_136),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_35),
.Y(n_468)
);

BUFx5_ASAP7_75t_L g469 ( 
.A(n_279),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_246),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_68),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_256),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_17),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_290),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_303),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_27),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_293),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_291),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_146),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_10),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_3),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_307),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_45),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_126),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_268),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_227),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_59),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_54),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_177),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_48),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_14),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_111),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_259),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_135),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_285),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_310),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_18),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_292),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_257),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_275),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_222),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_281),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_231),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_163),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_195),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_244),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_261),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_23),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_155),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_203),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_102),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_69),
.Y(n_512)
);

BUFx10_ASAP7_75t_L g513 ( 
.A(n_283),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_92),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_140),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_106),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_104),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_107),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_33),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_209),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_304),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_289),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_86),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_120),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_320),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_365),
.B(n_94),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_342),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_0),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_342),
.B(n_1),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_342),
.B(n_1),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_365),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_2),
.Y(n_532)
);

BUFx12f_ASAP7_75t_L g533 ( 
.A(n_320),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_365),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_365),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_376),
.B(n_3),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_342),
.B(n_4),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_320),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_376),
.B(n_6),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_439),
.B(n_7),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_359),
.B(n_7),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_342),
.Y(n_546)
);

BUFx12f_ASAP7_75t_L g547 ( 
.A(n_419),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_342),
.B(n_8),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_359),
.B(n_8),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_448),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_315),
.Y(n_551)
);

BUFx12f_ASAP7_75t_L g552 ( 
.A(n_315),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_417),
.B(n_9),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_325),
.B(n_11),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_509),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_97),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_418),
.B(n_12),
.Y(n_559)
);

INVx5_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_382),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_382),
.B(n_13),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_405),
.B(n_13),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_448),
.Y(n_564)
);

BUFx12f_ASAP7_75t_L g565 ( 
.A(n_499),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_405),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_355),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_342),
.B(n_341),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_415),
.B(n_14),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_341),
.B(n_16),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_312),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_355),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_354),
.B(n_17),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_311),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_481),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_472),
.B(n_18),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_481),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_313),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_481),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_517),
.B(n_354),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_366),
.B(n_20),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_389),
.B(n_20),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_427),
.B(n_21),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_407),
.B(n_21),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_407),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_411),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_411),
.B(n_412),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_317),
.Y(n_594)
);

BUFx8_ASAP7_75t_L g595 ( 
.A(n_406),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_326),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_412),
.B(n_22),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_329),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_427),
.B(n_22),
.Y(n_599)
);

BUFx8_ASAP7_75t_L g600 ( 
.A(n_406),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_513),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_413),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_437),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_314),
.Y(n_604)
);

BUFx12f_ASAP7_75t_L g605 ( 
.A(n_316),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_497),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_437),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_497),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_402),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_453),
.B(n_24),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_453),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_414),
.B(n_24),
.Y(n_612)
);

INVx5_ASAP7_75t_L g613 ( 
.A(n_474),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_345),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_482),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_372),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_395),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_408),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_324),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_26),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_327),
.B(n_328),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_27),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_334),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_358),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_504),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_318),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_319),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_410),
.B(n_28),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_321),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_339),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_346),
.B(n_28),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_323),
.Y(n_633)
);

BUFx8_ASAP7_75t_L g634 ( 
.A(n_433),
.Y(n_634)
);

INVx5_ASAP7_75t_L g635 ( 
.A(n_358),
.Y(n_635)
);

BUFx12f_ASAP7_75t_L g636 ( 
.A(n_369),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_331),
.B(n_29),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_337),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_340),
.B(n_29),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_434),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_348),
.B(n_30),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_446),
.B(n_31),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_322),
.B(n_32),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_377),
.B(n_33),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_379),
.B(n_34),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_384),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_351),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_352),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_358),
.Y(n_649)
);

INVx6_ASAP7_75t_L g650 ( 
.A(n_358),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_358),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_358),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_332),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_451),
.B(n_35),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_358),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_464),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_469),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_385),
.Y(n_658)
);

BUFx8_ASAP7_75t_L g659 ( 
.A(n_465),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_360),
.B(n_36),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_353),
.B(n_36),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_480),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_469),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_490),
.B(n_37),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_491),
.Y(n_665)
);

BUFx12f_ASAP7_75t_L g666 ( 
.A(n_386),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_391),
.B(n_37),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_330),
.B(n_38),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_361),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_512),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_363),
.B(n_38),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_371),
.B(n_39),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_378),
.B(n_39),
.Y(n_673)
);

BUFx12f_ASAP7_75t_L g674 ( 
.A(n_399),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_383),
.B(n_40),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_362),
.B(n_40),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_400),
.B(n_42),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_556),
.A2(n_430),
.B1(n_431),
.B2(n_428),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_612),
.A2(n_373),
.B1(n_381),
.B2(n_338),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_543),
.A2(n_409),
.B1(n_420),
.B2(n_403),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_574),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_582),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_580),
.Y(n_683)
);

AO22x2_ASAP7_75t_L g684 ( 
.A1(n_543),
.A2(n_422),
.B1(n_435),
.B2(n_429),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_545),
.B(n_440),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_528),
.A2(n_444),
.B1(n_449),
.B2(n_447),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_556),
.A2(n_455),
.B1(n_456),
.B2(n_452),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_621),
.A2(n_394),
.B1(n_396),
.B2(n_392),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_549),
.A2(n_404),
.B1(n_478),
.B2(n_397),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_L g690 ( 
.A1(n_587),
.A2(n_462),
.B1(n_473),
.B2(n_468),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_550),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_550),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_562),
.A2(n_442),
.B1(n_475),
.B2(n_450),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_587),
.A2(n_483),
.B1(n_488),
.B2(n_476),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_668),
.A2(n_523),
.B1(n_508),
.B2(n_471),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_622),
.B(n_416),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_609),
.B(n_459),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_554),
.A2(n_485),
.B1(n_489),
.B2(n_461),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_561),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_531),
.Y(n_701)
);

INVx8_ASAP7_75t_L g702 ( 
.A(n_609),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_531),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_R g704 ( 
.A1(n_536),
.A2(n_501),
.B1(n_505),
.B2(n_494),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_580),
.Y(n_705)
);

AO22x2_ASAP7_75t_L g706 ( 
.A1(n_562),
.A2(n_514),
.B1(n_515),
.B2(n_511),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_534),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_668),
.A2(n_518),
.B1(n_524),
.B2(n_516),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_534),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_532),
.A2(n_335),
.B1(n_336),
.B2(n_333),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_534),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_540),
.A2(n_344),
.B1(n_347),
.B2(n_343),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_613),
.B(n_349),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_SL g714 ( 
.A1(n_643),
.A2(n_356),
.B1(n_357),
.B2(n_350),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_661),
.A2(n_367),
.B1(n_368),
.B2(n_364),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_613),
.B(n_370),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_SL g717 ( 
.A1(n_632),
.A2(n_375),
.B1(n_380),
.B2(n_374),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_583),
.B(n_658),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_676),
.A2(n_390),
.B1(n_393),
.B2(n_387),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_563),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_544),
.A2(n_401),
.B1(n_421),
.B2(n_398),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_594),
.B(n_423),
.Y(n_722)
);

AO22x2_ASAP7_75t_L g723 ( 
.A1(n_563),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_620),
.B(n_424),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_605),
.A2(n_426),
.B1(n_432),
.B2(n_425),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_535),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_671),
.A2(n_522),
.B1(n_521),
.B2(n_520),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_535),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_535),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_570),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_585),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_573),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_597),
.B(n_47),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_585),
.Y(n_734)
);

BUFx6f_ASAP7_75t_SL g735 ( 
.A(n_551),
.Y(n_735)
);

AO22x2_ASAP7_75t_L g736 ( 
.A1(n_570),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_736)
);

AND2x2_ASAP7_75t_SL g737 ( 
.A(n_597),
.B(n_51),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_591),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_646),
.B(n_436),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_541),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_671),
.A2(n_510),
.B1(n_507),
.B2(n_506),
.Y(n_741)
);

AO22x2_ASAP7_75t_L g742 ( 
.A1(n_581),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_629),
.A2(n_503),
.B1(n_502),
.B2(n_500),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_601),
.B(n_438),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_624),
.A2(n_467),
.B1(n_496),
.B2(n_495),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_579),
.Y(n_746)
);

CKINVDCx6p67_ASAP7_75t_R g747 ( 
.A(n_601),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_541),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_653),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_541),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_601),
.B(n_441),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_672),
.A2(n_498),
.B1(n_492),
.B2(n_486),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_631),
.A2(n_484),
.B1(n_479),
.B2(n_477),
.Y(n_753)
);

INVx8_ASAP7_75t_L g754 ( 
.A(n_552),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_568),
.B(n_445),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_636),
.A2(n_470),
.B1(n_454),
.B2(n_466),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_576),
.B(n_457),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_672),
.A2(n_458),
.B1(n_460),
.B2(n_463),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_581),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_553),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_591),
.Y(n_761)
);

INVx1_ASAP7_75t_SL g762 ( 
.A(n_666),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_591),
.Y(n_763)
);

OR2x6_ASAP7_75t_L g764 ( 
.A(n_674),
.B(n_57),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_559),
.A2(n_469),
.B1(n_59),
.B2(n_60),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_645),
.A2(n_469),
.B1(n_60),
.B2(n_61),
.Y(n_766)
);

OAI22xp33_ASAP7_75t_L g767 ( 
.A1(n_675),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_572),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_565),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_553),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_553),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_572),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_644),
.A2(n_469),
.B1(n_71),
.B2(n_72),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_555),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_577),
.A2(n_610),
.B1(n_590),
.B2(n_629),
.Y(n_775)
);

OR2x6_ASAP7_75t_L g776 ( 
.A(n_547),
.B(n_525),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_571),
.B(n_469),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_683),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_700),
.B(n_586),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_705),
.Y(n_780)
);

INVx4_ASAP7_75t_SL g781 ( 
.A(n_777),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_775),
.B(n_594),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_697),
.B(n_606),
.Y(n_783)
);

INVxp33_ASAP7_75t_L g784 ( 
.A(n_755),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_738),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_761),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_702),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_763),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_740),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_740),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_748),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_748),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_685),
.B(n_527),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_701),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_703),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_707),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_709),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_679),
.B(n_662),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_726),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_729),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_750),
.Y(n_803)
);

XOR2xp5_ASAP7_75t_L g804 ( 
.A(n_688),
.B(n_662),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_760),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_770),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_686),
.B(n_571),
.Y(n_807)
);

XOR2xp5_ASAP7_75t_L g808 ( 
.A(n_689),
.B(n_537),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_771),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_774),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_728),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_699),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_691),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_757),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_773),
.B(n_623),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_691),
.Y(n_816)
);

XOR2xp5_ASAP7_75t_L g817 ( 
.A(n_746),
.B(n_537),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_731),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_685),
.A2(n_530),
.B(n_529),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_734),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_728),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_728),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_724),
.B(n_586),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_692),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_681),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_690),
.B(n_596),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_682),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_713),
.B(n_546),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_718),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_680),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_680),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_684),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_684),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_733),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_765),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_693),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

XNOR2xp5_ASAP7_75t_L g838 ( 
.A(n_762),
.B(n_667),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_720),
.B(n_723),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_706),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_739),
.B(n_606),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_752),
.A2(n_569),
.B(n_593),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_706),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_737),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_716),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_744),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_766),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_SL g848 ( 
.A(n_696),
.B(n_526),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_720),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_730),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_730),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_736),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_736),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_742),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_742),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_747),
.B(n_606),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_759),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_759),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_732),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_702),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_698),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_708),
.Y(n_863)
);

INVx4_ASAP7_75t_SL g864 ( 
.A(n_743),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_715),
.B(n_598),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_714),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_710),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_719),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_722),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_735),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_754),
.B(n_764),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_721),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_678),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_793),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_793),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_823),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_869),
.B(n_749),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_819),
.B(n_589),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_828),
.B(n_727),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_778),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_828),
.B(n_741),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_823),
.B(n_758),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_778),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_779),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_819),
.B(n_599),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_780),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_780),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_783),
.B(n_637),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_818),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_845),
.B(n_639),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_847),
.B(n_639),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_846),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_848),
.B(n_826),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_842),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_779),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_820),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_870),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_813),
.Y(n_899)
);

AND2x2_ASAP7_75t_SL g900 ( 
.A(n_848),
.B(n_623),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_782),
.B(n_641),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_816),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_781),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_863),
.Y(n_904)
);

AND2x2_ASAP7_75t_SL g905 ( 
.A(n_826),
.B(n_641),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_811),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_862),
.B(n_660),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_821),
.Y(n_908)
);

AND2x2_ASAP7_75t_SL g909 ( 
.A(n_866),
.B(n_660),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_830),
.B(n_673),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_822),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_829),
.B(n_673),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_841),
.B(n_677),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_868),
.A2(n_548),
.B(n_538),
.Y(n_914)
);

AND2x2_ASAP7_75t_SL g915 ( 
.A(n_834),
.B(n_677),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_784),
.B(n_604),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_784),
.B(n_604),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_781),
.Y(n_918)
);

AND2x2_ASAP7_75t_SL g919 ( 
.A(n_834),
.B(n_538),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_831),
.B(n_548),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_844),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_870),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_825),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_814),
.B(n_617),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_827),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_824),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_835),
.B(n_617),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_781),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_797),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_835),
.B(n_619),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_867),
.B(n_592),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_802),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_844),
.B(n_619),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_785),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_872),
.B(n_786),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_839),
.B(n_640),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_865),
.B(n_717),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_839),
.B(n_640),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_873),
.B(n_656),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_787),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_788),
.B(n_592),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_832),
.B(n_625),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_794),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_859),
.B(n_656),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_795),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_796),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_787),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_798),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_799),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_801),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_833),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_803),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_805),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_836),
.B(n_670),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_837),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_807),
.B(n_712),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_840),
.B(n_843),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_808),
.B(n_695),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_815),
.B(n_603),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_853),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_815),
.B(n_603),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_806),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_809),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_810),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_815),
.B(n_603),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_789),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_790),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_815),
.B(n_791),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_792),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_849),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_850),
.B(n_577),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_886),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_921),
.B(n_804),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_SL g975 ( 
.A(n_898),
.B(n_860),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_876),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_903),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_924),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_880),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_880),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_876),
.B(n_864),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_893),
.B(n_815),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_893),
.B(n_851),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_893),
.B(n_852),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_927),
.B(n_854),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_886),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_887),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_874),
.B(n_875),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_876),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_898),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_877),
.B(n_812),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_887),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_892),
.Y(n_994)
);

BUFx8_ASAP7_75t_SL g995 ( 
.A(n_922),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_874),
.B(n_855),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_883),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_875),
.B(n_856),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_959),
.Y(n_999)
);

BUFx4f_ASAP7_75t_L g1000 ( 
.A(n_972),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_892),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_892),
.B(n_864),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_916),
.B(n_838),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_900),
.B(n_858),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_927),
.B(n_933),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_922),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_897),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_957),
.B(n_812),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_884),
.B(n_895),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_883),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_909),
.B(n_853),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_916),
.B(n_817),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_917),
.B(n_857),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_903),
.B(n_861),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_933),
.B(n_871),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_906),
.Y(n_1016)
);

AND2x2_ASAP7_75t_SL g1017 ( 
.A(n_905),
.B(n_590),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_936),
.B(n_871),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_889),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_889),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_908),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_903),
.B(n_725),
.Y(n_1022)
);

CKINVDCx8_ASAP7_75t_R g1023 ( 
.A(n_920),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_924),
.Y(n_1024)
);

OR2x6_ASAP7_75t_L g1025 ( 
.A(n_936),
.B(n_754),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_895),
.B(n_745),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_938),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_961),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_906),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_900),
.B(n_687),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_908),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_952),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_967),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_938),
.B(n_753),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_918),
.B(n_756),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_918),
.B(n_751),
.Y(n_1036)
);

AND2x6_ASAP7_75t_L g1037 ( 
.A(n_878),
.B(n_610),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_944),
.B(n_764),
.Y(n_1038)
);

AND2x6_ASAP7_75t_L g1039 ( 
.A(n_878),
.B(n_588),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_944),
.B(n_614),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_L g1041 ( 
.A(n_972),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_929),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_930),
.B(n_776),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_939),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_930),
.B(n_776),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_929),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_950),
.B(n_533),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_910),
.B(n_614),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_901),
.B(n_769),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_900),
.B(n_607),
.Y(n_1050)
);

BUFx2_ASAP7_75t_SL g1051 ( 
.A(n_918),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_905),
.B(n_578),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_901),
.B(n_608),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_977),
.B(n_918),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_973),
.Y(n_1056)
);

BUFx5_ASAP7_75t_L g1057 ( 
.A(n_1033),
.Y(n_1057)
);

INVx3_ASAP7_75t_SL g1058 ( 
.A(n_991),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_997),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_977),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1028),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_SL g1062 ( 
.A(n_1006),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_982),
.B(n_905),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_1016),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_981),
.B(n_958),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_994),
.Y(n_1066)
);

CKINVDCx14_ASAP7_75t_R g1067 ( 
.A(n_1012),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_994),
.B(n_928),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_1028),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_1017),
.B(n_909),
.Y(n_1070)
);

INVxp67_ASAP7_75t_SL g1071 ( 
.A(n_1016),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_994),
.B(n_928),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_1001),
.B(n_928),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1005),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_1029),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_1001),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_1025),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1007),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_1029),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_1002),
.B(n_942),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_997),
.Y(n_1081)
);

INVx8_ASAP7_75t_L g1082 ( 
.A(n_1018),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_1027),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_1021),
.B(n_940),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_1025),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_973),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_1027),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_999),
.Y(n_1088)
);

INVx1_ASAP7_75t_SL g1089 ( 
.A(n_1024),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1032),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_993),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_1032),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1007),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1021),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1003),
.B(n_919),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_1015),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_976),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1021),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_975),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_989),
.Y(n_1101)
);

INVx6_ASAP7_75t_L g1102 ( 
.A(n_976),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1010),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_974),
.B(n_904),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_987),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_SL g1106 ( 
.A(n_1045),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_988),
.Y(n_1107)
);

CKINVDCx6p67_ASAP7_75t_R g1108 ( 
.A(n_1045),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_981),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_978),
.B(n_919),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1023),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_1031),
.B(n_976),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1019),
.Y(n_1113)
);

BUFx5_ASAP7_75t_L g1114 ( 
.A(n_1033),
.Y(n_1114)
);

BUFx10_ASAP7_75t_L g1115 ( 
.A(n_1034),
.Y(n_1115)
);

BUFx5_ASAP7_75t_L g1116 ( 
.A(n_1037),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_986),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_990),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1008),
.A2(n_919),
.B1(n_915),
.B2(n_909),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1060),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1070),
.A2(n_1039),
.B1(n_1041),
.B2(n_1000),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1059),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_SL g1123 ( 
.A1(n_1119),
.A2(n_1052),
.B1(n_992),
.B2(n_937),
.Y(n_1123)
);

CKINVDCx14_ASAP7_75t_R g1124 ( 
.A(n_1055),
.Y(n_1124)
);

INVx6_ASAP7_75t_L g1125 ( 
.A(n_1098),
.Y(n_1125)
);

CKINVDCx10_ASAP7_75t_R g1126 ( 
.A(n_1106),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1101),
.B(n_984),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1061),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1061),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1101),
.A2(n_985),
.B1(n_1011),
.B2(n_1030),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1095),
.A2(n_1039),
.B1(n_1037),
.B2(n_1034),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1081),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1110),
.B(n_1037),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1067),
.A2(n_1049),
.B(n_1043),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1074),
.B(n_1004),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1099),
.B(n_1031),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1100),
.A2(n_915),
.B1(n_885),
.B2(n_999),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1069),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1056),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1091),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1097),
.Y(n_1141)
);

BUFx8_ASAP7_75t_SL g1142 ( 
.A(n_1055),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1090),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1067),
.A2(n_1038),
.B(n_1013),
.Y(n_1144)
);

INVx6_ASAP7_75t_L g1145 ( 
.A(n_1098),
.Y(n_1145)
);

CKINVDCx20_ASAP7_75t_R g1146 ( 
.A(n_1062),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_1088),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1062),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1086),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1106),
.A2(n_885),
.B1(n_914),
.B2(n_542),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1103),
.Y(n_1151)
);

BUFx8_ASAP7_75t_L g1152 ( 
.A(n_1077),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1105),
.Y(n_1153)
);

INVx6_ASAP7_75t_L g1154 ( 
.A(n_1066),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1063),
.A2(n_1026),
.B1(n_882),
.B2(n_1044),
.Y(n_1155)
);

BUFx10_ASAP7_75t_L g1156 ( 
.A(n_1065),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1107),
.Y(n_1157)
);

CKINVDCx6p67_ASAP7_75t_R g1158 ( 
.A(n_1058),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1113),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1104),
.A2(n_996),
.B1(n_998),
.B2(n_907),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1096),
.A2(n_1048),
.B1(n_1040),
.B2(n_920),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1064),
.A2(n_1050),
.B1(n_1051),
.B2(n_879),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1065),
.A2(n_1040),
.B1(n_920),
.B2(n_1009),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_1085),
.Y(n_1164)
);

CKINVDCx14_ASAP7_75t_R g1165 ( 
.A(n_1078),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1117),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1111),
.A2(n_920),
.B1(n_1009),
.B2(n_1053),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1117),
.A2(n_1020),
.B1(n_896),
.B2(n_935),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1064),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_1058),
.Y(n_1170)
);

INVx8_ASAP7_75t_L g1171 ( 
.A(n_1082),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1071),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1066),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1071),
.A2(n_881),
.B(n_931),
.Y(n_1174)
);

CKINVDCx14_ASAP7_75t_R g1175 ( 
.A(n_1093),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1075),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1092),
.Y(n_1177)
);

CKINVDCx11_ASAP7_75t_R g1178 ( 
.A(n_1108),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1075),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_1089),
.A2(n_767),
.B(n_1022),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1115),
.A2(n_990),
.B1(n_891),
.B2(n_890),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_SL g1182 ( 
.A(n_1152),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1123),
.A2(n_704),
.B1(n_1115),
.B2(n_1092),
.Y(n_1183)
);

OAI222xp33_ASAP7_75t_L g1184 ( 
.A1(n_1137),
.A2(n_772),
.B1(n_768),
.B2(n_642),
.C1(n_664),
.C2(n_654),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1143),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_SL g1186 ( 
.A1(n_1150),
.A2(n_1035),
.B(n_890),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_L g1187 ( 
.A(n_1158),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1135),
.B(n_1109),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1135),
.B(n_1109),
.Y(n_1189)
);

AOI211xp5_ASAP7_75t_L g1190 ( 
.A1(n_1180),
.A2(n_654),
.B(n_664),
.C(n_912),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1137),
.A2(n_1080),
.B1(n_960),
.B2(n_966),
.Y(n_1191)
);

OAI222xp33_ASAP7_75t_L g1192 ( 
.A1(n_1150),
.A2(n_1080),
.B1(n_962),
.B2(n_593),
.C1(n_896),
.C2(n_969),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1122),
.Y(n_1193)
);

INVxp33_ASAP7_75t_L g1194 ( 
.A(n_1177),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1136),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1177),
.B(n_1083),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1139),
.Y(n_1197)
);

OAI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1155),
.A2(n_912),
.B(n_913),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1136),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1130),
.A2(n_1082),
.B1(n_1116),
.B2(n_659),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1134),
.A2(n_1047),
.B1(n_923),
.B2(n_925),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_1142),
.B(n_1083),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1132),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1127),
.B(n_1087),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1144),
.A2(n_1121),
.B(n_1131),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1167),
.A2(n_942),
.B1(n_1051),
.B2(n_1087),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1170),
.Y(n_1207)
);

OAI21xp33_ASAP7_75t_L g1208 ( 
.A1(n_1161),
.A2(n_888),
.B(n_923),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1181),
.A2(n_1163),
.B1(n_1127),
.B2(n_1160),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1128),
.B(n_956),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1130),
.A2(n_1116),
.B1(n_659),
.B2(n_634),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1160),
.A2(n_1102),
.B1(n_1112),
.B2(n_1084),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1166),
.B(n_891),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1149),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1120),
.B(n_1099),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1168),
.B(n_888),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1126),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1174),
.A2(n_926),
.B(n_945),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1146),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1133),
.A2(n_963),
.B1(n_1116),
.B2(n_934),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1151),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1157),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1138),
.A2(n_1102),
.B1(n_1118),
.B2(n_1014),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1159),
.A2(n_1118),
.B1(n_1036),
.B2(n_1094),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1171),
.A2(n_1116),
.B1(n_600),
.B2(n_595),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1140),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1129),
.A2(n_1094),
.B1(n_899),
.B2(n_1072),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1120),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1162),
.A2(n_1116),
.B1(n_600),
.B2(n_595),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1174),
.A2(n_963),
.B1(n_934),
.B2(n_902),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1153),
.A2(n_963),
.B1(n_934),
.B2(n_902),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1141),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1148),
.B(n_899),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1162),
.A2(n_934),
.B1(n_953),
.B2(n_948),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_SL g1235 ( 
.A1(n_1165),
.A2(n_955),
.B(n_910),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1175),
.A2(n_955),
.B(n_910),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1164),
.A2(n_934),
.B1(n_953),
.B2(n_948),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1169),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1172),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1176),
.A2(n_1068),
.B1(n_1073),
.B2(n_1072),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1179),
.A2(n_949),
.B(n_945),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1204),
.B(n_1171),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1183),
.A2(n_964),
.B1(n_567),
.B2(n_575),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1183),
.A2(n_567),
.B1(n_575),
.B2(n_561),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1188),
.B(n_469),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1200),
.B(n_1057),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1198),
.A2(n_1211),
.B1(n_1209),
.B2(n_1208),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1211),
.A2(n_567),
.B1(n_575),
.B2(n_561),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1216),
.A2(n_1124),
.B1(n_1171),
.B2(n_1152),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1189),
.B(n_1173),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1200),
.A2(n_584),
.B1(n_951),
.B2(n_949),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1238),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1201),
.A2(n_584),
.B1(n_954),
.B2(n_1156),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1233),
.A2(n_1156),
.B1(n_1178),
.B2(n_911),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1229),
.A2(n_911),
.B1(n_908),
.B2(n_968),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1229),
.A2(n_558),
.B1(n_526),
.B2(n_970),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1190),
.A2(n_941),
.B(n_970),
.Y(n_1257)
);

OAI222xp33_ASAP7_75t_L g1258 ( 
.A1(n_1185),
.A2(n_569),
.B1(n_1046),
.B2(n_1042),
.C1(n_665),
.C2(n_618),
.Y(n_1258)
);

OAI21xp33_ASAP7_75t_L g1259 ( 
.A1(n_1186),
.A2(n_665),
.B(n_618),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1239),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1191),
.A2(n_1147),
.B1(n_1057),
.B2(n_1114),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1218),
.B(n_1241),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1192),
.A2(n_980),
.B(n_979),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1235),
.A2(n_1154),
.B1(n_1145),
.B2(n_1125),
.Y(n_1264)
);

OAI222xp33_ASAP7_75t_L g1265 ( 
.A1(n_1213),
.A2(n_983),
.B1(n_1079),
.B2(n_965),
.C1(n_946),
.C2(n_971),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1194),
.B(n_1066),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1205),
.A2(n_965),
.B1(n_967),
.B2(n_943),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1206),
.A2(n_943),
.B1(n_967),
.B2(n_932),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1196),
.B(n_1076),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1236),
.A2(n_1154),
.B1(n_1145),
.B2(n_1125),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1193),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1226),
.B(n_1076),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1225),
.A2(n_943),
.B1(n_906),
.B2(n_1079),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1212),
.A2(n_1114),
.B1(n_1057),
.B2(n_894),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1192),
.A2(n_1073),
.B(n_1068),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1232),
.B(n_1057),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1184),
.A2(n_971),
.B1(n_669),
.B2(n_647),
.C(n_633),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1187),
.A2(n_1224),
.B1(n_1202),
.B2(n_1223),
.Y(n_1278)
);

NAND3xp33_ASAP7_75t_L g1279 ( 
.A(n_1237),
.B(n_628),
.C(n_627),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1210),
.A2(n_894),
.B1(n_1057),
.B2(n_1114),
.Y(n_1280)
);

OAI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1220),
.A2(n_1187),
.B1(n_1234),
.B2(n_1230),
.C(n_1231),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1197),
.B(n_1114),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1203),
.B(n_1214),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1221),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1222),
.B(n_894),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_L g1286 ( 
.A(n_1227),
.B(n_628),
.C(n_627),
.Y(n_1286)
);

AOI222xp33_ASAP7_75t_L g1287 ( 
.A1(n_1207),
.A2(n_650),
.B1(n_669),
.B2(n_648),
.C1(n_638),
.C2(n_630),
.Y(n_1287)
);

OAI22x1_ASAP7_75t_L g1288 ( 
.A1(n_1228),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1182),
.A2(n_1054),
.B1(n_947),
.B2(n_602),
.Y(n_1289)
);

OAI221xp5_ASAP7_75t_L g1290 ( 
.A1(n_1219),
.A2(n_947),
.B1(n_638),
.B2(n_630),
.C(n_657),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1240),
.A2(n_615),
.B1(n_607),
.B2(n_611),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1195),
.A2(n_611),
.B1(n_626),
.B2(n_615),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1195),
.A2(n_616),
.B1(n_626),
.B2(n_655),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1199),
.A2(n_616),
.B1(n_663),
.B2(n_652),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1199),
.A2(n_1215),
.B1(n_1182),
.B2(n_1217),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1278),
.B(n_555),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1250),
.B(n_70),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1245),
.B(n_73),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1283),
.B(n_76),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1283),
.B(n_77),
.Y(n_1300)
);

OAI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1244),
.A2(n_557),
.B(n_80),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1271),
.B(n_81),
.Y(n_1302)
);

OAI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1243),
.A2(n_651),
.B1(n_649),
.B2(n_635),
.C(n_83),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1242),
.B(n_81),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1249),
.B(n_557),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1295),
.B(n_1254),
.Y(n_1306)
);

NOR3xp33_ASAP7_75t_L g1307 ( 
.A(n_1258),
.B(n_82),
.C(n_84),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1247),
.B(n_557),
.Y(n_1308)
);

AOI221xp5_ASAP7_75t_L g1309 ( 
.A1(n_1288),
.A2(n_651),
.B1(n_649),
.B2(n_88),
.C(n_89),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1287),
.B(n_1248),
.C(n_1277),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1284),
.B(n_84),
.Y(n_1311)
);

NOR3xp33_ASAP7_75t_L g1312 ( 
.A(n_1259),
.B(n_85),
.C(n_88),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1284),
.B(n_90),
.Y(n_1313)
);

OAI221xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1251),
.A2(n_91),
.B1(n_98),
.B2(n_103),
.C(n_105),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1262),
.B(n_539),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1252),
.B(n_109),
.Y(n_1316)
);

OA21x2_ASAP7_75t_L g1317 ( 
.A1(n_1246),
.A2(n_110),
.B(n_112),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1257),
.B(n_566),
.C(n_564),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1260),
.B(n_114),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1267),
.B(n_539),
.Y(n_1320)
);

AND2x2_ASAP7_75t_SL g1321 ( 
.A(n_1263),
.B(n_115),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1269),
.B(n_118),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1266),
.B(n_121),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1267),
.A2(n_560),
.B1(n_539),
.B2(n_124),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1260),
.B(n_131),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1261),
.B(n_133),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1253),
.A2(n_560),
.B1(n_141),
.B2(n_143),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1276),
.B(n_137),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1285),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1290),
.A2(n_144),
.B(n_145),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1272),
.B(n_156),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1280),
.B(n_1274),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1255),
.A2(n_157),
.B(n_158),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1282),
.B(n_168),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1307),
.A2(n_1281),
.B1(n_1256),
.B2(n_1263),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_L g1336 ( 
.A(n_1307),
.B(n_1273),
.C(n_1286),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1329),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1302),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1297),
.B(n_1275),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1298),
.B(n_1268),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1304),
.B(n_1264),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1309),
.B(n_1291),
.C(n_1279),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1321),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1299),
.B(n_1270),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1300),
.B(n_1289),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1312),
.A2(n_1301),
.B1(n_1310),
.B2(n_1303),
.Y(n_1346)
);

OAI211xp5_ASAP7_75t_L g1347 ( 
.A1(n_1312),
.A2(n_1292),
.B(n_1293),
.C(n_1294),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1317),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1315),
.B(n_173),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1311),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1351)
);

NOR2x1_ASAP7_75t_L g1352 ( 
.A(n_1318),
.B(n_178),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1313),
.B(n_180),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1332),
.B(n_184),
.Y(n_1354)
);

NAND4xp75_ASAP7_75t_L g1355 ( 
.A(n_1296),
.B(n_185),
.C(n_189),
.D(n_190),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1306),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1316),
.B(n_197),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1337),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1348),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1346),
.B(n_1314),
.C(n_1317),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_1305),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1337),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1350),
.B(n_1319),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1348),
.B(n_1325),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1343),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1343),
.B(n_1326),
.Y(n_1366)
);

AOI211xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1356),
.A2(n_1330),
.B(n_1333),
.C(n_1324),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1339),
.B(n_1344),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1341),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1345),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1335),
.B(n_1328),
.Y(n_1371)
);

XNOR2xp5_ASAP7_75t_L g1372 ( 
.A(n_1346),
.B(n_1323),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1340),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1351),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1351),
.B(n_1322),
.Y(n_1375)
);

OA22x2_ASAP7_75t_L g1376 ( 
.A1(n_1372),
.A2(n_1354),
.B1(n_1308),
.B2(n_1353),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_R g1377 ( 
.A(n_1375),
.B(n_1349),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1358),
.Y(n_1378)
);

NOR2x1_ASAP7_75t_L g1379 ( 
.A(n_1369),
.B(n_1352),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1362),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1364),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1358),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1373),
.B(n_1357),
.Y(n_1383)
);

XNOR2xp5_ASAP7_75t_L g1384 ( 
.A(n_1372),
.B(n_1355),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_1363),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1370),
.B(n_1336),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1364),
.Y(n_1387)
);

AO22x2_ASAP7_75t_L g1388 ( 
.A1(n_1374),
.A2(n_1342),
.B1(n_1320),
.B2(n_1347),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1373),
.B(n_1368),
.Y(n_1389)
);

AO22x2_ASAP7_75t_L g1390 ( 
.A1(n_1374),
.A2(n_1327),
.B1(n_1331),
.B2(n_1334),
.Y(n_1390)
);

AOI22x1_ASAP7_75t_L g1391 ( 
.A1(n_1384),
.A2(n_1375),
.B1(n_1359),
.B2(n_1367),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1385),
.A2(n_1361),
.B1(n_1371),
.B2(n_1360),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1386),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1386),
.Y(n_1394)
);

OAI22x1_ASAP7_75t_L g1395 ( 
.A1(n_1379),
.A2(n_1368),
.B1(n_1365),
.B2(n_1366),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1389),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1380),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1381),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1382),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1381),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1383),
.Y(n_1401)
);

OA22x2_ASAP7_75t_L g1402 ( 
.A1(n_1387),
.A2(n_1388),
.B1(n_1376),
.B2(n_1377),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1398),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1400),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1401),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1397),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1402),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1399),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1396),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1393),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1394),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1407),
.A2(n_1392),
.B1(n_1391),
.B2(n_1376),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1408),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1403),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1404),
.Y(n_1415)
);

OA22x2_ASAP7_75t_L g1416 ( 
.A1(n_1405),
.A2(n_1395),
.B1(n_1378),
.B2(n_1390),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1406),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1414),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1415),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1413),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1412),
.A2(n_1409),
.B1(n_1410),
.B2(n_1411),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1416),
.Y(n_1422)
);

AOI31xp33_ASAP7_75t_L g1423 ( 
.A1(n_1417),
.A2(n_199),
.A3(n_201),
.B(n_206),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1418),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_L g1425 ( 
.A(n_1422),
.B(n_213),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1419),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1420),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1421),
.B(n_217),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1426),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1424),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1427),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1425),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1429),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1432),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1430),
.B(n_1428),
.Y(n_1435)
);

INVxp33_ASAP7_75t_SL g1436 ( 
.A(n_1431),
.Y(n_1436)
);

NOR3xp33_ASAP7_75t_L g1437 ( 
.A(n_1432),
.B(n_1423),
.C(n_223),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1436),
.A2(n_220),
.B1(n_224),
.B2(n_226),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1433),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1435),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1437),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1434),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1434),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1439),
.Y(n_1444)
);

OAI22x1_ASAP7_75t_L g1445 ( 
.A1(n_1440),
.A2(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1441),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_1446)
);

AOI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1442),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_1447)
);

OAI22x1_ASAP7_75t_L g1448 ( 
.A1(n_1443),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_1448)
);

AO22x2_ASAP7_75t_L g1449 ( 
.A1(n_1438),
.A2(n_253),
.B1(n_258),
.B2(n_260),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1439),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1444),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1450),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1449),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1449),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1445),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1452),
.A2(n_1446),
.B1(n_1448),
.B2(n_1447),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1455),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1456),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1457),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1458),
.A2(n_1454),
.B1(n_1453),
.B2(n_1451),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1459),
.A2(n_274),
.B1(n_276),
.B2(n_278),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1460),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1462),
.A2(n_1461),
.B1(n_284),
.B2(n_287),
.C(n_288),
.Y(n_1463)
);

AOI211xp5_ASAP7_75t_L g1464 ( 
.A1(n_1463),
.A2(n_294),
.B(n_295),
.C(n_297),
.Y(n_1464)
);


endmodule