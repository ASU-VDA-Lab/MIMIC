module fake_jpeg_32180_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_1),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_1),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_59),
.B1(n_74),
.B2(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_98),
.B1(n_58),
.B2(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_68),
.B1(n_75),
.B2(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_106),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_81),
.B(n_80),
.C(n_79),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_109),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_72),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_66),
.B1(n_74),
.B2(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_64),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_115),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_117),
.B1(n_21),
.B2(n_48),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_61),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_63),
.B1(n_75),
.B2(n_57),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_52),
.B1(n_71),
.B2(n_26),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_68),
.B1(n_65),
.B2(n_62),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_132),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_71),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_3),
.Y(n_125)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_22),
.B(n_50),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_19),
.B(n_30),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_3),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_40),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_32),
.B1(n_47),
.B2(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_139),
.B1(n_121),
.B2(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_145),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_15),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_152),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_16),
.B(n_18),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_151),
.B(n_157),
.Y(n_171)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g164 ( 
.A(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_160),
.B1(n_120),
.B2(n_43),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_37),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_38),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_141),
.B(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_51),
.B1(n_41),
.B2(n_42),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_144),
.B1(n_149),
.B2(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_162),
.B(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_169),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_179),
.B1(n_166),
.B2(n_167),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_177),
.Y(n_181)
);

OAI221xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_175),
.B1(n_165),
.B2(n_171),
.C(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_147),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_148),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_142),
.Y(n_188)
);


endmodule