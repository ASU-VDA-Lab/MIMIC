module fake_jpeg_10783_n_477 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_477);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_477;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_68),
.B1(n_50),
.B2(n_41),
.Y(n_120)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_58),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_61),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_62),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_63),
.B(n_64),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_20),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_75),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_77),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_25),
.B(n_15),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_79),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_28),
.B(n_48),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_80),
.B(n_14),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_86),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_46),
.B(n_1),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_11),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_96),
.Y(n_125)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_33),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_12),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_37),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_38),
.B(n_12),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_38),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_117),
.Y(n_184)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_12),
.Y(n_117)
);

BUFx16f_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_120),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_45),
.B1(n_48),
.B2(n_47),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_122),
.A2(n_123),
.B1(n_131),
.B2(n_138),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_51),
.B1(n_49),
.B2(n_43),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_35),
.B1(n_50),
.B2(n_41),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_96),
.A2(n_34),
.B1(n_49),
.B2(n_43),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_57),
.A2(n_35),
.B1(n_21),
.B2(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_68),
.A2(n_21),
.B1(n_40),
.B2(n_30),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_39),
.B1(n_34),
.B2(n_30),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_39),
.B1(n_40),
.B2(n_6),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_143),
.A2(n_145),
.B1(n_150),
.B2(n_152),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_89),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_182),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_70),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_94),
.A2(n_7),
.B1(n_14),
.B2(n_83),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_82),
.A2(n_7),
.B1(n_73),
.B2(n_66),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_155),
.A2(n_158),
.B1(n_160),
.B2(n_169),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_7),
.B1(n_114),
.B2(n_116),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_69),
.A2(n_58),
.B1(n_105),
.B2(n_60),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_56),
.A2(n_62),
.B1(n_99),
.B2(n_97),
.Y(n_169)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_99),
.A2(n_93),
.B1(n_103),
.B2(n_90),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_95),
.A2(n_102),
.B1(n_88),
.B2(n_87),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_176),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_85),
.A2(n_109),
.B1(n_101),
.B2(n_67),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_196),
.B1(n_123),
.B2(n_183),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_84),
.B1(n_71),
.B2(n_98),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_185),
.Y(n_255)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_112),
.A2(n_118),
.B1(n_81),
.B2(n_104),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_118),
.A2(n_104),
.B1(n_32),
.B2(n_96),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_96),
.A2(n_32),
.B1(n_54),
.B2(n_119),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_198),
.A2(n_215),
.B1(n_260),
.B2(n_263),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_199),
.B(n_210),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

AO22x1_ASAP7_75t_SL g201 ( 
.A1(n_126),
.A2(n_127),
.B1(n_124),
.B2(n_132),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_201),
.B(n_253),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_171),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_230),
.B(n_240),
.Y(n_271)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_203),
.Y(n_299)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_204),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_209),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_180),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_129),
.B(n_181),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_208),
.B(n_220),
.C(n_223),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_184),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_137),
.B(n_184),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_212),
.B(n_227),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_213),
.B(n_219),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_148),
.B(n_153),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_136),
.B(n_171),
.C(n_144),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_125),
.B(n_159),
.C(n_130),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_135),
.B(n_165),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_226),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_187),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_138),
.B(n_150),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_143),
.A2(n_196),
.B(n_195),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_162),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_231),
.B(n_237),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_232),
.Y(n_305)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_141),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_236),
.Y(n_297)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_157),
.Y(n_235)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_142),
.B(n_154),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_162),
.B(n_156),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_166),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_156),
.B(n_168),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_243),
.A2(n_249),
.B(n_256),
.Y(n_300)
);

BUFx4f_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx11_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_192),
.A2(n_169),
.B(n_174),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_247),
.A2(n_217),
.B(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_170),
.B(n_178),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_167),
.B(n_179),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_151),
.B(n_133),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_163),
.B(n_186),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_258),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_146),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_263),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx6_ASAP7_75t_SL g261 ( 
.A(n_146),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_238),
.Y(n_307)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_160),
.B1(n_217),
.B2(n_262),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_277),
.B1(n_279),
.B2(n_285),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_202),
.A2(n_201),
.B(n_220),
.C(n_208),
.Y(n_273)
);

A2O1A1Ixp33_ASAP7_75t_L g340 ( 
.A1(n_273),
.A2(n_300),
.B(n_307),
.C(n_296),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_250),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_255),
.B1(n_216),
.B2(n_229),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_246),
.A2(n_229),
.B1(n_198),
.B2(n_257),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_306),
.B1(n_286),
.B2(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_201),
.B1(n_198),
.B2(n_230),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_208),
.A2(n_202),
.B(n_253),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_296),
.B(n_270),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_198),
.A2(n_247),
.B1(n_223),
.B2(n_261),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_224),
.B(n_252),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_286),
.A2(n_244),
.B(n_211),
.Y(n_316)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_221),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_274),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_206),
.A2(n_248),
.B(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_301),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_214),
.B(n_222),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_235),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_203),
.A2(n_233),
.B1(n_241),
.B2(n_260),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_317),
.Y(n_350)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_211),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_313),
.B(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_316),
.A2(n_326),
.B(n_291),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_275),
.B(n_200),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_325),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_232),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_320),
.B(n_335),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_267),
.A2(n_270),
.B1(n_279),
.B2(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_328),
.B1(n_332),
.B2(n_305),
.Y(n_361)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_269),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_324),
.B(n_341),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_250),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_297),
.A2(n_244),
.B1(n_285),
.B2(n_273),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_272),
.A2(n_271),
.B1(n_282),
.B2(n_264),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_329),
.A2(n_346),
.B1(n_306),
.B2(n_299),
.Y(n_359)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_330),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_331),
.B(n_336),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_347),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_308),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_268),
.C(n_287),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_297),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_298),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_276),
.A2(n_281),
.B1(n_280),
.B2(n_292),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_337),
.A2(n_305),
.B1(n_265),
.B2(n_283),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_269),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_338),
.Y(n_349)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_340),
.B(n_329),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_303),
.A2(n_289),
.B(n_290),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_303),
.Y(n_342)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_268),
.B(n_290),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_343),
.Y(n_352)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_345),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_276),
.A2(n_292),
.B1(n_266),
.B2(n_287),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_360),
.C(n_366),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_313),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_371),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_314),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_359),
.A2(n_322),
.B1(n_315),
.B2(n_317),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_288),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_361),
.A2(n_376),
.B1(n_319),
.B2(n_325),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_299),
.C(n_288),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_343),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_373),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_288),
.B(n_291),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_312),
.B(n_299),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_322),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_349),
.A2(n_321),
.B1(n_326),
.B2(n_328),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_389),
.B(n_398),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_361),
.A2(n_314),
.B1(n_353),
.B2(n_354),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_380),
.A2(n_393),
.B1(n_352),
.B2(n_357),
.Y(n_417)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_381),
.Y(n_404)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_383),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_374),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_351),
.B(n_331),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_386),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_375),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_388),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_375),
.B(n_338),
.Y(n_386)
);

XOR2x2_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_350),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_349),
.A2(n_318),
.B1(n_332),
.B2(n_335),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_336),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_348),
.C(n_364),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_365),
.B(n_327),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_395),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_364),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_355),
.A2(n_340),
.B1(n_320),
.B2(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_401),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_359),
.A2(n_311),
.B1(n_316),
.B2(n_339),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_391),
.B(n_358),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_408),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_414),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_366),
.C(n_356),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_407),
.B(n_409),
.C(n_410),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_356),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_354),
.C(n_353),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_389),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_394),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_388),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_369),
.C(n_371),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_412),
.B(n_378),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_369),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_365),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_417),
.A2(n_418),
.B1(n_401),
.B2(n_395),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_380),
.A2(n_352),
.B1(n_362),
.B2(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_423),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_385),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_381),
.B(n_382),
.C(n_378),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_428),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_413),
.B1(n_421),
.B2(n_419),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_427),
.B(n_403),
.Y(n_447)
);

BUFx12_ASAP7_75t_L g428 ( 
.A(n_421),
.Y(n_428)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_402),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_429),
.B(n_430),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_383),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_330),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_431),
.A2(n_434),
.B1(n_435),
.B2(n_418),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_409),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_406),
.B(n_342),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_437),
.B(n_441),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_408),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_445),
.Y(n_453)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_440),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_425),
.A2(n_417),
.B1(n_413),
.B2(n_412),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_447),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_407),
.C(n_416),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_433),
.C(n_424),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_426),
.A2(n_419),
.B1(n_410),
.B2(n_400),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_428),
.A2(n_372),
.B(n_316),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_448),
.A2(n_373),
.B(n_428),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_427),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_452),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_437),
.B(n_424),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_443),
.A2(n_441),
.B(n_448),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_454),
.B(n_440),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_455),
.B(n_444),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_457),
.B(n_445),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_459),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_446),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_460),
.Y(n_465)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_464),
.B(n_457),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_438),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_462),
.A2(n_463),
.B(n_450),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_469),
.Y(n_471)
);

AOI322xp5_ASAP7_75t_L g470 ( 
.A1(n_467),
.A2(n_453),
.A3(n_390),
.B1(n_436),
.B2(n_377),
.C1(n_370),
.C2(n_368),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_461),
.A2(n_453),
.B(n_447),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_472),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_468),
.B(n_362),
.Y(n_472)
);

AOI322xp5_ASAP7_75t_L g473 ( 
.A1(n_471),
.A2(n_465),
.A3(n_390),
.B1(n_377),
.B2(n_370),
.C1(n_265),
.C2(n_367),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_473),
.B(n_346),
.C(n_347),
.Y(n_475)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_475),
.A2(n_345),
.B1(n_474),
.B2(n_291),
.C(n_305),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_283),
.B(n_265),
.Y(n_477)
);


endmodule