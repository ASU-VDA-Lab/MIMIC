module real_jpeg_29583_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_0),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_56),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_1),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_81),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_81),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_26),
.B1(n_33),
.B2(n_81),
.Y(n_197)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_32),
.B1(n_40),
.B2(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_42),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_58),
.B(n_62),
.C(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_5),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_5),
.B(n_60),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_5),
.B(n_40),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_40),
.B(n_44),
.C(n_182),
.D(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_72),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_25),
.B(n_195),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_5),
.A2(n_64),
.B(n_76),
.C(n_112),
.D(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_64),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_26),
.B1(n_33),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_7),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_50),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_10),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_11),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_119)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_12),
.B(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_12),
.B(n_26),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_13),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_67),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_227)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_21),
.B(n_113),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_82),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_22),
.B(n_82),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_54),
.C(n_68),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_38),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_25),
.A2(n_36),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_25),
.A2(n_34),
.B(n_85),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_25),
.A2(n_84),
.B1(n_105),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_25),
.A2(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_25),
.B(n_197),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_29),
.A2(n_203),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_29),
.B(n_100),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_31),
.A2(n_35),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_33),
.A2(n_41),
.A3(n_46),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_33),
.B(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g84 ( 
.A(n_35),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_39),
.A2(n_51),
.B(n_146),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_40),
.A2(n_63),
.A3(n_224),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_41),
.B(n_74),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_43),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_44),
.A2(n_48),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_44),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_44),
.A2(n_48),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_51),
.B(n_148),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_51),
.A2(n_146),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_51),
.B(n_100),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_59),
.A2(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_60),
.B(n_96),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_64),
.B(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_66),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_70),
.A2(n_71),
.B1(n_108),
.B2(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_80),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_71),
.A2(n_75),
.B(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_72),
.A2(n_76),
.B1(n_110),
.B2(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_89),
.A2(n_90),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_106),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_92),
.B1(n_106),
.B2(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B(n_95),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_103),
.A2(n_198),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_111),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_133),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_132),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_174),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_158),
.B(n_173),
.Y(n_137)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_155),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_143),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.C(n_152),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_159),
.B(n_161),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_162),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_167),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_168),
.B(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_170),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_252),
.C(n_253),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_247),
.B(n_251),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_235),
.B(n_246),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_219),
.B(n_234),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_199),
.B(n_218),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_184),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_211),
.B(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_217),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_216),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_221),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_237),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);


endmodule