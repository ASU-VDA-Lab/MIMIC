module real_jpeg_29978_n_18 (n_17, n_8, n_0, n_2, n_10, n_338, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_338;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_0),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_0),
.A2(n_56),
.B1(n_58),
.B2(n_96),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_0),
.A2(n_61),
.B1(n_62),
.B2(n_96),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_28),
.B1(n_56),
.B2(n_58),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_1),
.A2(n_28),
.B1(n_61),
.B2(n_62),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_2),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_111),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_111),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_2),
.A2(n_56),
.B1(n_58),
.B2(n_111),
.Y(n_204)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_4),
.B(n_56),
.Y(n_116)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_51),
.B1(n_56),
.B2(n_58),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_277)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_94),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_7),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_94),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_7),
.A2(n_56),
.B1(n_58),
.B2(n_94),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_8),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_56),
.B1(n_58),
.B2(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_285)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_37),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_37),
.B1(n_56),
.B2(n_58),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_11),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_101),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_56),
.B1(n_58),
.B2(n_101),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_101),
.Y(n_258)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_13),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_30),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_13),
.B(n_32),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_61),
.B(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_61),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_13),
.B(n_74),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_13),
.A2(n_119),
.B1(n_138),
.B2(n_204),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_13),
.A2(n_33),
.B(n_219),
.Y(n_218)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_16),
.A2(n_61),
.B1(n_62),
.B2(n_72),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_17),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_17),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_17),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_22),
.B(n_43),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_24),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_26),
.A2(n_35),
.B(n_108),
.C(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_32),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_32),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_29),
.A2(n_32),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_29),
.A2(n_32),
.B1(n_146),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_29),
.A2(n_32),
.B1(n_165),
.B2(n_258),
.Y(n_257)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_68),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_33),
.A2(n_62),
.A3(n_68),
.B1(n_220),
.B2(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_34),
.B(n_108),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_82),
.B(n_333),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_75),
.C(n_77),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_44),
.A2(n_45),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_64),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_46),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_48),
.A2(n_79),
.B1(n_81),
.B2(n_285),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_52),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_52),
.A2(n_64),
.B1(n_311),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_53),
.A2(n_59),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_53),
.A2(n_59),
.B1(n_136),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_53),
.A2(n_59),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_53),
.A2(n_59),
.B1(n_179),
.B2(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_53),
.B(n_108),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_53),
.A2(n_59),
.B1(n_100),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_53),
.A2(n_59),
.B1(n_63),
.B2(n_267),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_54),
.A2(n_58),
.A3(n_61),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_55),
.B(n_56),
.Y(n_183)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_56),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_61),
.B(n_72),
.Y(n_228)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_73),
.B2(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_65),
.A2(n_66),
.B1(n_74),
.B2(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_74),
.B1(n_93),
.B2(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_66),
.A2(n_74),
.B1(n_149),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_66),
.A2(n_74),
.B1(n_167),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_71),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_71),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_67),
.A2(n_71),
.B1(n_95),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_67),
.A2(n_71),
.B1(n_127),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_67),
.A2(n_71),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_75),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_79),
.A2(n_81),
.B1(n_110),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_79),
.A2(n_81),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_326),
.B(n_332),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_302),
.A3(n_321),
.B1(n_324),
.B2(n_325),
.C(n_337),
.Y(n_83)
);

AOI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_254),
.A3(n_291),
.B1(n_296),
.B2(n_301),
.C(n_338),
.Y(n_84)
);

NOR3xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_151),
.C(n_169),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_131),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_87),
.B(n_131),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_112),
.C(n_123),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_88),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_106),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_98),
.C(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_102),
.A2(n_105),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_102),
.A2(n_105),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_108),
.B(n_119),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_112),
.A2(n_123),
.B1(n_124),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_112),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_116),
.A2(n_118),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_138),
.B1(n_140),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_119),
.A2(n_138),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_119),
.A2(n_138),
.B1(n_198),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_119),
.A2(n_138),
.B1(n_193),
.B2(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_119),
.A2(n_138),
.B(n_158),
.Y(n_269)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_130),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_125),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_128),
.B(n_130),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_129),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_141),
.C(n_142),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_137),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.C(n_150),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g297 ( 
.A1(n_152),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_153),
.B(n_154),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_168),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_156),
.B(n_161),
.C(n_168),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_157),
.B(n_159),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_160),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_248),
.B(n_253),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_234),
.B(n_247),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_213),
.B(n_233),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_194),
.B(n_212),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_174),
.B(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_211),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_200),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_210),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_215),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_217),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_225),
.C(n_232),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_250),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_271),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_255),
.B(n_271),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.C(n_270),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_262),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_256),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.CI(n_261),
.CON(n_256),
.SN(n_256)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_258),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_260),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_268),
.B2(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_263),
.B(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_269),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_268),
.A2(n_283),
.B(n_286),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_289),
.B2(n_290),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_280),
.C(n_290),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_278),
.B(n_279),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_277),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_304),
.C(n_313),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_279),
.B(n_304),
.CI(n_313),
.CON(n_323),
.SN(n_323)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_292),
.A2(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_314),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_305),
.A2(n_306),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.C(n_311),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_319),
.C(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_323),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule