module real_aes_382_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_0), .A2(n_13), .B1(n_156), .B2(n_158), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_1), .A2(n_69), .B1(n_134), .B2(n_138), .Y(n_133) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_2), .A2(n_55), .B1(n_95), .B2(n_99), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_3), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_3), .Y(n_184) );
INVx1_ASAP7_75t_L g201 ( .A(n_4), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_5), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g174 ( .A(n_6), .Y(n_174) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_7), .A2(n_20), .B1(n_95), .B2(n_96), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_8), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_9), .A2(n_71), .B1(n_88), .B2(n_109), .Y(n_87) );
INVx2_ASAP7_75t_L g221 ( .A(n_10), .Y(n_221) );
INVx1_ASAP7_75t_L g291 ( .A(n_11), .Y(n_291) );
INVx1_ASAP7_75t_L g183 ( .A(n_12), .Y(n_183) );
INVx1_ASAP7_75t_L g288 ( .A(n_14), .Y(n_288) );
INVx1_ASAP7_75t_SL g342 ( .A(n_15), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_15), .A2(n_83), .B1(n_84), .B2(n_342), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_16), .B(n_241), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_17), .A2(n_179), .B1(n_186), .B2(n_187), .Y(n_178) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_17), .Y(n_186) );
AOI33xp33_ASAP7_75t_L g328 ( .A1(n_18), .A2(n_41), .A3(n_226), .B1(n_234), .B2(n_329), .B3(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g265 ( .A(n_19), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g193 ( .A1(n_20), .A2(n_55), .B1(n_58), .B2(n_194), .C(n_196), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_21), .A2(n_43), .B1(n_143), .B2(n_145), .Y(n_142) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_22), .A2(n_70), .B(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g251 ( .A(n_22), .B(n_70), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_23), .B(n_224), .Y(n_339) );
INVx3_ASAP7_75t_L g95 ( .A(n_24), .Y(n_95) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_25), .A2(n_39), .B1(n_114), .B2(n_118), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_26), .A2(n_52), .B1(n_163), .B2(n_167), .Y(n_162) );
INVx1_ASAP7_75t_SL g104 ( .A(n_27), .Y(n_104) );
INVx1_ASAP7_75t_L g203 ( .A(n_28), .Y(n_203) );
AND2x2_ASAP7_75t_L g229 ( .A(n_28), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g247 ( .A(n_28), .B(n_201), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_29), .A2(n_40), .B1(n_124), .B2(n_128), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_30), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_31), .B(n_224), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_32), .A2(n_219), .B1(n_282), .B2(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g177 ( .A(n_33), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_33), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_34), .B(n_241), .Y(n_343) );
INVx1_ASAP7_75t_L g595 ( .A(n_34), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_35), .B(n_255), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_36), .B(n_241), .Y(n_258) );
AO22x2_ASAP7_75t_L g107 ( .A1(n_37), .A2(n_58), .B1(n_95), .B2(n_108), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_38), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_42), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g227 ( .A(n_44), .Y(n_227) );
INVx1_ASAP7_75t_L g243 ( .A(n_44), .Y(n_243) );
AND2x2_ASAP7_75t_L g248 ( .A(n_45), .B(n_249), .Y(n_248) );
AOI221xp5_ASAP7_75t_L g256 ( .A1(n_46), .A2(n_60), .B1(n_224), .B2(n_232), .C(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_47), .B(n_224), .Y(n_316) );
INVx1_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_49), .B(n_219), .Y(n_274) );
AOI21xp5_ASAP7_75t_SL g312 ( .A1(n_50), .A2(n_232), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g285 ( .A(n_51), .Y(n_285) );
INVx1_ASAP7_75t_L g238 ( .A(n_53), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_54), .A2(n_232), .B(n_237), .Y(n_231) );
INVxp33_ASAP7_75t_L g198 ( .A(n_55), .Y(n_198) );
INVx1_ASAP7_75t_L g230 ( .A(n_56), .Y(n_230) );
INVx1_ASAP7_75t_L g245 ( .A(n_56), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_57), .B(n_224), .Y(n_331) );
INVxp67_ASAP7_75t_L g197 ( .A(n_58), .Y(n_197) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_59), .A2(n_83), .B1(n_84), .B2(n_588), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_59), .Y(n_588) );
AND2x2_ASAP7_75t_L g344 ( .A(n_61), .B(n_218), .Y(n_344) );
INVx1_ASAP7_75t_L g286 ( .A(n_62), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_63), .A2(n_232), .B(n_341), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_64), .A2(n_232), .B(n_303), .C(n_307), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_65), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_66), .B(n_218), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_67), .A2(n_180), .B1(n_181), .B2(n_185), .Y(n_179) );
INVx1_ASAP7_75t_L g185 ( .A(n_67), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_68), .A2(n_232), .B1(n_326), .B2(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g314 ( .A(n_72), .Y(n_314) );
INVx1_ASAP7_75t_L g82 ( .A(n_73), .Y(n_82) );
AND2x2_ASAP7_75t_L g332 ( .A(n_74), .B(n_218), .Y(n_332) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_75), .A2(n_263), .B(n_264), .C(n_267), .Y(n_262) );
BUFx2_ASAP7_75t_SL g195 ( .A(n_76), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_77), .B(n_241), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_190), .B1(n_204), .B2(n_574), .C(n_579), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_172), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_84), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_141), .Y(n_85) );
NAND4xp25_ASAP7_75t_L g86 ( .A(n_87), .B(n_113), .C(n_123), .D(n_133), .Y(n_86) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx4_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx8_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x4_ASAP7_75t_L g91 ( .A(n_92), .B(n_100), .Y(n_91) );
AND2x2_ASAP7_75t_L g116 ( .A(n_92), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g136 ( .A(n_92), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g154 ( .A(n_92), .B(n_149), .Y(n_154) );
AND2x4_ASAP7_75t_L g92 ( .A(n_93), .B(n_97), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x4_ASAP7_75t_L g112 ( .A(n_94), .B(n_97), .Y(n_112) );
INVx1_ASAP7_75t_L g122 ( .A(n_94), .Y(n_122) );
AND2x2_ASAP7_75t_L g132 ( .A(n_94), .B(n_98), .Y(n_132) );
INVx2_ASAP7_75t_L g96 ( .A(n_95), .Y(n_96) );
INVx1_ASAP7_75t_L g99 ( .A(n_95), .Y(n_99) );
OAI22x1_ASAP7_75t_L g102 ( .A1(n_95), .A2(n_103), .B1(n_104), .B2(n_105), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_95), .Y(n_103) );
INVx1_ASAP7_75t_L g108 ( .A(n_95), .Y(n_108) );
INVxp67_ASAP7_75t_L g148 ( .A(n_97), .Y(n_148) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g121 ( .A(n_98), .B(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g120 ( .A(n_100), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g140 ( .A(n_100), .B(n_132), .Y(n_140) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_106), .Y(n_100) );
AND2x2_ASAP7_75t_L g117 ( .A(n_101), .B(n_107), .Y(n_117) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g137 ( .A(n_102), .B(n_106), .Y(n_137) );
AND2x2_ASAP7_75t_L g149 ( .A(n_102), .B(n_107), .Y(n_149) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_102), .Y(n_171) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g131 ( .A(n_107), .Y(n_131) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g144 ( .A(n_112), .B(n_117), .Y(n_144) );
AND2x2_ASAP7_75t_L g166 ( .A(n_112), .B(n_137), .Y(n_166) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx3_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g127 ( .A(n_117), .B(n_121), .Y(n_127) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx8_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g157 ( .A(n_121), .B(n_137), .Y(n_157) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx5_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_L g170 ( .A(n_132), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx6_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND4xp25_ASAP7_75t_L g141 ( .A(n_142), .B(n_150), .C(n_155), .D(n_162), .Y(n_141) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x4_ASAP7_75t_L g159 ( .A(n_149), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B1(n_175), .B2(n_189), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_174), .A2(n_239), .B(n_246), .C(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B1(n_178), .B2(n_188), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_178), .Y(n_188) );
INVx1_ASAP7_75t_L g187 ( .A(n_179), .Y(n_187) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
AND3x1_ASAP7_75t_SL g192 ( .A(n_193), .B(n_199), .C(n_202), .Y(n_192) );
INVxp67_ASAP7_75t_L g586 ( .A(n_193), .Y(n_586) );
CKINVDCx8_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g584 ( .A(n_199), .Y(n_584) );
AO21x1_ASAP7_75t_SL g592 ( .A1(n_199), .A2(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g225 ( .A(n_200), .B(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_SL g591 ( .A(n_200), .B(n_202), .Y(n_591) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g236 ( .A(n_201), .B(n_227), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_202), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2x1p5_ASAP7_75t_L g233 ( .A(n_203), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND4xp75_ASAP7_75t_L g207 ( .A(n_208), .B(n_446), .C(n_491), .D(n_560), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2x1_ASAP7_75t_L g209 ( .A(n_210), .B(n_406), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_362), .C(n_387), .Y(n_210) );
OAI222xp33_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_276), .B1(n_317), .B2(n_333), .C1(n_349), .C2(n_356), .Y(n_211) );
INVxp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_252), .Y(n_213) );
AND2x2_ASAP7_75t_L g571 ( .A(n_214), .B(n_385), .Y(n_571) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_216), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_216), .B(n_260), .Y(n_361) );
INVx3_ASAP7_75t_L g376 ( .A(n_216), .Y(n_376) );
AND2x2_ASAP7_75t_L g509 ( .A(n_216), .B(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_222), .B(n_248), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_217), .A2(n_218), .B1(n_262), .B2(n_268), .Y(n_261) );
AO21x2_ASAP7_75t_L g394 ( .A1(n_217), .A2(n_222), .B(n_248), .Y(n_394) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_219), .B(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_220), .Y(n_255) );
AND2x2_ASAP7_75t_SL g250 ( .A(n_221), .B(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g282 ( .A(n_221), .B(n_251), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_231), .Y(n_222) );
INVx1_ASAP7_75t_L g275 ( .A(n_224), .Y(n_275) );
AND2x4_ASAP7_75t_L g224 ( .A(n_225), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g299 ( .A(n_225), .Y(n_299) );
OR2x6_ASAP7_75t_L g239 ( .A(n_226), .B(n_235), .Y(n_239) );
INVxp33_ASAP7_75t_L g329 ( .A(n_226), .Y(n_329) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_226), .Y(n_594) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g293 ( .A(n_227), .B(n_244), .Y(n_293) );
INVx1_ASAP7_75t_L g300 ( .A(n_228), .Y(n_300) );
BUFx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g235 ( .A(n_230), .Y(n_235) );
AND2x6_ASAP7_75t_L g290 ( .A(n_230), .B(n_242), .Y(n_290) );
INVxp67_ASAP7_75t_L g273 ( .A(n_232), .Y(n_273) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_236), .Y(n_232) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_233), .Y(n_593) );
INVx1_ASAP7_75t_L g330 ( .A(n_234), .Y(n_330) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .C(n_246), .Y(n_237) );
INVxp67_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_239), .A2(n_266), .B1(n_285), .B2(n_286), .Y(n_284) );
INVx2_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_239), .A2(n_246), .B(n_314), .C(n_315), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g341 ( .A1(n_239), .A2(n_246), .B(n_342), .C(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g266 ( .A(n_241), .Y(n_266) );
AND2x4_ASAP7_75t_L g578 ( .A(n_241), .B(n_247), .Y(n_578) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_246), .B(n_282), .Y(n_294) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_246), .A2(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
INVx5_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_247), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_249), .Y(n_337) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g439 ( .A(n_252), .B(n_392), .Y(n_439) );
AND2x2_ASAP7_75t_L g441 ( .A(n_252), .B(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g476 ( .A(n_252), .Y(n_476) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_260), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_L g359 ( .A(n_254), .Y(n_359) );
INVx1_ASAP7_75t_L g378 ( .A(n_254), .Y(n_378) );
AND2x4_ASAP7_75t_L g385 ( .A(n_254), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_254), .B(n_323), .Y(n_401) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_254), .Y(n_510) );
INVx1_ASAP7_75t_L g520 ( .A(n_254), .Y(n_520) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_259), .Y(n_254) );
INVx2_ASAP7_75t_SL g307 ( .A(n_255), .Y(n_307) );
INVx1_ASAP7_75t_L g320 ( .A(n_260), .Y(n_320) );
INVx2_ASAP7_75t_L g373 ( .A(n_260), .Y(n_373) );
INVx1_ASAP7_75t_L g454 ( .A(n_260), .Y(n_454) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_273), .B1(n_274), .B2(n_275), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_SL g277 ( .A(n_278), .B(n_308), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_278), .B(n_335), .Y(n_429) );
INVx2_ASAP7_75t_L g450 ( .A(n_278), .Y(n_450) );
AND2x2_ASAP7_75t_L g458 ( .A(n_278), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_295), .Y(n_278) );
AND2x4_ASAP7_75t_L g348 ( .A(n_279), .B(n_296), .Y(n_348) );
INVx1_ASAP7_75t_L g355 ( .A(n_279), .Y(n_355) );
AND2x2_ASAP7_75t_L g531 ( .A(n_279), .B(n_336), .Y(n_531) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g369 ( .A(n_280), .B(n_296), .Y(n_369) );
INVx2_ASAP7_75t_L g405 ( .A(n_280), .Y(n_405) );
AND2x2_ASAP7_75t_L g484 ( .A(n_280), .B(n_336), .Y(n_484) );
NOR2x1_ASAP7_75t_SL g527 ( .A(n_280), .B(n_309), .Y(n_527) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_282), .A2(n_312), .B(n_316), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_294), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_291), .B2(n_292), .Y(n_287) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g367 ( .A(n_295), .Y(n_367) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g381 ( .A(n_296), .B(n_309), .Y(n_381) );
INVx1_ASAP7_75t_L g397 ( .A(n_296), .Y(n_397) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_296), .Y(n_505) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_302), .Y(n_296) );
NOR3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .C(n_301), .Y(n_298) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_307), .A2(n_324), .B(n_332), .Y(n_323) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_307), .A2(n_324), .B(n_332), .Y(n_374) );
AND2x2_ASAP7_75t_L g368 ( .A(n_308), .B(n_369), .Y(n_368) );
OR2x6_ASAP7_75t_L g449 ( .A(n_308), .B(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g487 ( .A(n_308), .B(n_484), .Y(n_487) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx4_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_309), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g416 ( .A(n_309), .Y(n_416) );
OR2x2_ASAP7_75t_L g422 ( .A(n_309), .B(n_336), .Y(n_422) );
AND2x4_ASAP7_75t_L g436 ( .A(n_309), .B(n_397), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_309), .B(n_405), .Y(n_437) );
OR2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g481 ( .A(n_320), .B(n_400), .Y(n_481) );
BUFx2_ASAP7_75t_L g533 ( .A(n_320), .Y(n_533) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g564 ( .A(n_322), .B(n_476), .Y(n_564) );
INVx2_ASAP7_75t_L g358 ( .A(n_323), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_325), .B(n_331), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_345), .Y(n_333) );
AND2x2_ASAP7_75t_L g380 ( .A(n_334), .B(n_381), .Y(n_380) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_335), .B(n_355), .Y(n_365) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g353 ( .A(n_336), .Y(n_353) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_336), .Y(n_459) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_336), .Y(n_526) );
INVx1_ASAP7_75t_L g566 ( .A(n_336), .Y(n_566) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_344), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
BUFx2_ASAP7_75t_L g480 ( .A(n_345), .Y(n_480) );
NOR2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AND2x4_ASAP7_75t_L g396 ( .A(n_346), .B(n_397), .Y(n_396) );
NOR2xp67_ASAP7_75t_SL g428 ( .A(n_346), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g501 ( .A(n_346), .B(n_484), .Y(n_501) );
AND2x4_ASAP7_75t_SL g504 ( .A(n_346), .B(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g553 ( .A(n_346), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g420 ( .A(n_347), .Y(n_420) );
INVx4_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g415 ( .A(n_348), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_348), .B(n_413), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_348), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_348), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g498 ( .A(n_352), .B(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g414 ( .A(n_353), .Y(n_414) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_357), .B(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g532 ( .A(n_357), .B(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g540 ( .A(n_357), .B(n_469), .Y(n_540) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g409 ( .A(n_358), .B(n_394), .Y(n_409) );
AND2x4_ASAP7_75t_L g442 ( .A(n_358), .B(n_376), .Y(n_442) );
INVx1_ASAP7_75t_L g559 ( .A(n_358), .Y(n_559) );
AND2x2_ASAP7_75t_L g445 ( .A(n_360), .B(n_385), .Y(n_445) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g466 ( .A(n_361), .B(n_401), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_370), .B1(n_379), .B2(n_382), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B(n_368), .Y(n_363) );
OAI22xp5_ASAP7_75t_SL g545 ( .A1(n_364), .A2(n_433), .B1(n_541), .B2(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_365), .B(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g434 ( .A(n_365), .B(n_366), .Y(n_434) );
AND2x2_ASAP7_75t_SL g464 ( .A(n_365), .B(n_436), .Y(n_464) );
AOI211xp5_ASAP7_75t_SL g552 ( .A1(n_365), .A2(n_553), .B(n_555), .C(n_556), .Y(n_552) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_366), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_366), .B(n_412), .Y(n_538) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g443 ( .A(n_368), .Y(n_443) );
INVx2_ASAP7_75t_L g499 ( .A(n_369), .Y(n_499) );
AND2x2_ASAP7_75t_L g573 ( .A(n_369), .B(n_566), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_370), .A2(n_522), .B(n_528), .Y(n_521) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g508 ( .A(n_372), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g518 ( .A(n_372), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x2_ASAP7_75t_L g425 ( .A(n_373), .B(n_378), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g427 ( .A(n_373), .B(n_394), .Y(n_427) );
AND2x2_ASAP7_75t_L g469 ( .A(n_373), .B(n_394), .Y(n_469) );
INVx2_ASAP7_75t_L g386 ( .A(n_374), .Y(n_386) );
AND2x4_ASAP7_75t_L g392 ( .A(n_374), .B(n_393), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx3_ASAP7_75t_L g384 ( .A(n_376), .Y(n_384) );
INVx3_ASAP7_75t_L g390 ( .A(n_377), .Y(n_390) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_381), .A2(n_487), .B(n_563), .Y(n_567) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_384), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_384), .B(n_459), .Y(n_474) );
OR2x2_ASAP7_75t_L g489 ( .A(n_384), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g496 ( .A(n_384), .B(n_400), .Y(n_496) );
AND2x2_ASAP7_75t_L g452 ( .A(n_385), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g468 ( .A(n_385), .B(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g485 ( .A(n_385), .B(n_454), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_395), .B1(n_398), .B2(n_402), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g462 ( .A(n_390), .B(n_391), .Y(n_462) );
NOR2xp67_ASAP7_75t_SL g500 ( .A(n_390), .B(n_408), .Y(n_500) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_394), .B(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g403 ( .A(n_396), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g467 ( .A(n_396), .B(n_413), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_396), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g570 ( .A(n_404), .B(n_436), .Y(n_570) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_405), .B(n_516), .Y(n_515) );
NOR2xp67_ASAP7_75t_SL g406 ( .A(n_407), .B(n_430), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_417), .C(n_426), .Y(n_407) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_408), .A2(n_461), .B(n_471), .C(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g550 ( .A(n_409), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g461 ( .A(n_413), .B(n_437), .Y(n_461) );
AND2x2_ASAP7_75t_L g548 ( .A(n_413), .B(n_527), .Y(n_548) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g516 ( .A(n_416), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_423), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_420), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
NAND2xp33_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_438), .B1(n_440), .B2(n_443), .C(n_444), .Y(n_430) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .C(n_435), .D(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g549 ( .A(n_436), .B(n_512), .Y(n_549) );
INVx2_ASAP7_75t_L g555 ( .A(n_436), .Y(n_555) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_439), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g542 ( .A(n_442), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NAND4xp75_ASAP7_75t_L g447 ( .A(n_448), .B(n_470), .C(n_477), .D(n_486), .Y(n_447) );
OA211x2_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_451), .B(n_455), .C(n_463), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_449), .B(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g543 ( .A(n_453), .Y(n_543) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g551 ( .A(n_454), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_456), .B(n_462), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g512 ( .A(n_459), .Y(n_512) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_468), .Y(n_463) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_467), .A2(n_518), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g546 ( .A(n_468), .Y(n_546) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_469), .B(n_559), .Y(n_558) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVxp67_ASAP7_75t_L g544 ( .A(n_480), .Y(n_544) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
AND2x2_ASAP7_75t_SL g503 ( .A(n_484), .B(n_504), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_485), .A2(n_548), .B1(n_570), .B2(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND3x1_ASAP7_75t_L g492 ( .A(n_493), .B(n_534), .C(n_547), .Y(n_492) );
NOR3x1_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .C(n_521), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_502), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_500), .B2(n_501), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_511), .B1(n_513), .B2(n_517), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g565 ( .A(n_515), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_532), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g554 ( .A(n_531), .Y(n_554) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_532), .A2(n_563), .B(n_565), .Y(n_562) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_545), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_539), .B1(n_541), .B2(n_544), .Y(n_535) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B(n_550), .C(n_552), .Y(n_547) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2x1_ASAP7_75t_SL g560 ( .A(n_561), .B(n_568), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_572), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_575), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI222xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_587), .B2(n_589), .C1(n_592), .C2(n_595), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
endmodule