module fake_netlist_1_3165_n_516 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_516);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_516;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_44), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_9), .Y(n_76) );
BUFx6f_ASAP7_75t_L g77 ( .A(n_48), .Y(n_77) );
BUFx2_ASAP7_75t_SL g78 ( .A(n_24), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_50), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_31), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_69), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_21), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_22), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_2), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_9), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_62), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_32), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
AND2x2_ASAP7_75t_L g95 ( .A(n_46), .B(n_73), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_35), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_16), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_23), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_5), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_55), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_13), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_4), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_47), .B(n_66), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_61), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_11), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_81), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_97), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_97), .Y(n_112) );
BUFx8_ASAP7_75t_L g113 ( .A(n_95), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_89), .Y(n_114) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_75), .A2(n_34), .B(n_72), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_89), .B(n_83), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_77), .B(n_0), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_101), .B(n_1), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_79), .B(n_2), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_76), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_84), .B(n_3), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_77), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_90), .B(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_87), .Y(n_132) );
OR2x2_ASAP7_75t_L g133 ( .A(n_116), .B(n_91), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_115), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_110), .Y(n_135) );
AOI22xp33_ASAP7_75t_L g136 ( .A1(n_124), .A2(n_88), .B1(n_108), .B2(n_79), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_110), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_115), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_125), .Y(n_140) );
AO22x2_ASAP7_75t_L g141 ( .A1(n_116), .A2(n_85), .B1(n_93), .B2(n_96), .Y(n_141) );
NAND2xp33_ASAP7_75t_L g142 ( .A(n_119), .B(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_118), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_118), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_119), .B(n_99), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_118), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_124), .B(n_95), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_112), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_120), .B(n_88), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_120), .B(n_90), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_123), .B(n_86), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_127), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_122), .B(n_94), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_111), .Y(n_158) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_147), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_134), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_135), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_145), .B(n_113), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_155), .B(n_113), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_153), .B(n_113), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_153), .B(n_131), .Y(n_167) );
INVx3_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_135), .Y(n_169) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_153), .B(n_105), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_133), .B(n_114), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_149), .B(n_123), .Y(n_174) );
INVx5_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
BUFx12f_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
NOR2xp67_ASAP7_75t_L g177 ( .A(n_151), .B(n_128), .Y(n_177) );
BUFx8_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
AND2x2_ASAP7_75t_SL g183 ( .A(n_153), .B(n_105), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_149), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_154), .B(n_142), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_157), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_138), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_141), .A2(n_122), .B1(n_126), .B2(n_129), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_146), .Y(n_191) );
INVxp67_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_170), .A2(n_141), .B1(n_149), .B2(n_157), .Y(n_193) );
BUFx3_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
AND3x2_ASAP7_75t_L g195 ( .A(n_192), .B(n_85), .C(n_93), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_175), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_170), .A2(n_149), .B1(n_141), .B2(n_157), .Y(n_201) );
AOI21xp33_ASAP7_75t_L g202 ( .A1(n_163), .A2(n_141), .B(n_136), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_184), .B(n_157), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_160), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_170), .B(n_151), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_183), .B(n_157), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_176), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_176), .B(n_104), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_171), .Y(n_211) );
OAI221xp5_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_129), .B1(n_132), .B2(n_128), .C(n_158), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_183), .A2(n_132), .B1(n_158), .B2(n_144), .Y(n_213) );
INVx2_ASAP7_75t_SL g214 ( .A(n_175), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_171), .Y(n_215) );
INVx2_ASAP7_75t_SL g216 ( .A(n_175), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_161), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_185), .A2(n_143), .B(n_144), .C(n_156), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_175), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_173), .B(n_148), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_183), .B(n_152), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_184), .B(n_175), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_184), .B(n_152), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
OAI221xp5_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_189), .B1(n_166), .B2(n_165), .C(n_167), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_217), .Y(n_227) );
OAI211xp5_ASAP7_75t_L g228 ( .A1(n_201), .A2(n_177), .B(n_174), .C(n_117), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_197), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_198), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_201), .A2(n_178), .B1(n_181), .B2(n_175), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_209), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_207), .A2(n_181), .B1(n_188), .B2(n_179), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_207), .A2(n_179), .B1(n_188), .B2(n_186), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_186), .B1(n_168), .B2(n_187), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_213), .A2(n_169), .B1(n_190), .B2(n_187), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_217), .Y(n_240) );
OAI221xp5_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_177), .B1(n_190), .B2(n_182), .C(n_161), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_211), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g243 ( .A1(n_212), .A2(n_159), .B1(n_164), .B2(n_182), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_215), .Y(n_245) );
AO31x2_ASAP7_75t_L g246 ( .A1(n_218), .A2(n_148), .A3(n_111), .B(n_117), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_215), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_225), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_225), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
NOR2x1p5_ASAP7_75t_L g252 ( .A(n_203), .B(n_159), .Y(n_252) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_226), .A2(n_202), .B1(n_210), .B2(n_222), .C(n_103), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_206), .B(n_196), .Y(n_254) );
AOI322xp5_ASAP7_75t_L g255 ( .A1(n_251), .A2(n_108), .A3(n_103), .B1(n_121), .B2(n_98), .C1(n_100), .C2(n_102), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_252), .B(n_203), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g257 ( .A1(n_241), .A2(n_203), .B1(n_219), .B2(n_194), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_243), .A2(n_208), .B1(n_219), .B2(n_194), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_204), .B1(n_198), .B2(n_169), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_204), .B1(n_168), .B2(n_224), .C(n_156), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_227), .Y(n_261) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_250), .A2(n_130), .B(n_92), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_240), .A2(n_112), .B1(n_224), .B2(n_78), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_228), .A2(n_112), .B1(n_146), .B2(n_168), .C(n_98), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_233), .B(n_191), .Y(n_267) );
OAI21xp5_ASAP7_75t_SL g268 ( .A1(n_234), .A2(n_195), .B(n_223), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_235), .Y(n_269) );
INVx11_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
OAI211xp5_ASAP7_75t_L g271 ( .A1(n_237), .A2(n_112), .B(n_109), .C(n_92), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_245), .B(n_223), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_245), .A2(n_78), .B1(n_148), .B2(n_150), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_247), .A2(n_148), .B1(n_150), .B2(n_134), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_269), .B(n_247), .Y(n_275) );
OAI31xp33_ASAP7_75t_SL g276 ( .A1(n_259), .A2(n_248), .A3(n_249), .B(n_244), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_253), .B(n_248), .C(n_249), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_261), .B(n_235), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_265), .B(n_246), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_264), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_258), .A2(n_231), .B1(n_236), .B2(n_244), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_267), .B(n_270), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_257), .A2(n_231), .B1(n_235), .B2(n_244), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_256), .A2(n_223), .B1(n_242), .B2(n_239), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_262), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_268), .B(n_107), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_272), .B(n_229), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_256), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_263), .B(n_246), .Y(n_292) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_254), .A2(n_250), .B(n_229), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_263), .A2(n_223), .B1(n_242), .B2(n_239), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_262), .B(n_230), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_271), .B(n_246), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_275), .B(n_246), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_275), .B(n_246), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_278), .B(n_246), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_287), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_230), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_289), .B(n_262), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_285), .A2(n_273), .B1(n_266), .B2(n_260), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_289), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_295), .B(n_77), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_284), .B(n_288), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_277), .A2(n_273), .B1(n_94), .B2(n_106), .C(n_77), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_292), .A2(n_94), .B1(n_106), .B2(n_274), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_295), .B(n_77), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_291), .B(n_255), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_292), .B(n_77), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_280), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_276), .B(n_106), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_280), .B(n_4), .Y(n_320) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_286), .A2(n_274), .B1(n_199), .B2(n_220), .C(n_216), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_282), .Y(n_323) );
INVx5_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_282), .B(n_250), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_308), .B(n_296), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_314), .A2(n_296), .B1(n_281), .B2(n_294), .C(n_130), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_304), .B(n_283), .Y(n_330) );
AOI211xp5_ASAP7_75t_L g331 ( .A1(n_310), .A2(n_276), .B(n_283), .C(n_130), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_290), .Y(n_333) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_317), .B(n_5), .C(n_6), .D(n_7), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_298), .B(n_6), .C(n_7), .D(n_8), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_304), .B(n_290), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_290), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_8), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_300), .B(n_10), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_309), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_10), .Y(n_342) );
AND2x4_ASAP7_75t_SL g343 ( .A(n_305), .B(n_313), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_298), .B(n_11), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_302), .B(n_12), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_324), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_302), .B(n_12), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_13), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_305), .B(n_14), .Y(n_350) );
XOR2xp5_ASAP7_75t_L g351 ( .A(n_320), .B(n_16), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_320), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_297), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_318), .B(n_150), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_318), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_326), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_323), .B(n_150), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_326), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_322), .B(n_150), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_325), .B(n_139), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_297), .B(n_139), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_301), .B(n_139), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_301), .B(n_139), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_312), .B(n_134), .Y(n_367) );
NOR3xp33_ASAP7_75t_SL g368 ( .A(n_319), .B(n_17), .C(n_18), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_343), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_343), .B(n_316), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_339), .B(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_341), .B(n_316), .Y(n_373) );
XOR2x2_ASAP7_75t_L g374 ( .A(n_351), .B(n_307), .Y(n_374) );
AOI31xp33_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_307), .A3(n_311), .B(n_321), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_336), .B(n_316), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_331), .B(n_324), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_346), .B(n_315), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_356), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_315), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_332), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_327), .B(n_315), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_338), .B(n_315), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_339), .B(n_324), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_334), .B(n_324), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_352), .B(n_324), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_338), .B(n_324), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
XOR2xp5_ASAP7_75t_L g390 ( .A(n_340), .B(n_19), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_359), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_330), .B(n_25), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_346), .B(n_198), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_328), .A2(n_160), .B1(n_172), .B2(n_180), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_340), .B(n_26), .Y(n_396) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_345), .B(n_164), .C(n_30), .D(n_33), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_342), .A2(n_160), .B1(n_172), .B2(n_180), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_342), .B(n_29), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_333), .B(n_37), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_353), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_363), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_345), .B(n_38), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_347), .B(n_39), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_333), .B(n_40), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_348), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_337), .B(n_41), .Y(n_408) );
INVx3_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
O2A1O1Ixp33_ASAP7_75t_L g410 ( .A1(n_347), .A2(n_220), .B(n_214), .C(n_199), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_344), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_348), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_355), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_374), .A2(n_344), .B(n_368), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_369), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_387), .B(n_350), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_402), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_371), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_387), .B(n_361), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_412), .B(n_362), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_381), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_407), .B(n_358), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_391), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_390), .B(n_367), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_377), .B(n_366), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_375), .B(n_365), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
XOR2x2_ASAP7_75t_L g431 ( .A(n_377), .B(n_364), .Y(n_431) );
XNOR2xp5_ASAP7_75t_L g432 ( .A(n_370), .B(n_364), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_388), .B(n_42), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_411), .B(n_43), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_385), .B(n_378), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_393), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_393), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_406), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_384), .Y(n_440) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_376), .A2(n_214), .B1(n_180), .B2(n_172), .C1(n_198), .C2(n_196), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_386), .B(n_45), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_379), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_409), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_372), .B(n_382), .Y(n_445) );
XOR2x2_ASAP7_75t_L g446 ( .A(n_385), .B(n_49), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_386), .B(n_51), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_397), .B(n_206), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_378), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_380), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_383), .B(n_54), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_410), .A2(n_56), .B(n_57), .C(n_58), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_60), .A3(n_63), .B(n_64), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_410), .A2(n_206), .B(n_205), .Y(n_455) );
XOR2x2_ASAP7_75t_L g456 ( .A(n_404), .B(n_65), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_413), .B(n_67), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_408), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_400), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_405), .B(n_68), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_398), .B(n_70), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_396), .B(n_399), .C(n_403), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_398), .B(n_196), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_395), .A2(n_196), .B(n_205), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_392), .A2(n_198), .B1(n_205), .B2(n_206), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_395), .B(n_205), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_377), .A2(n_205), .B(n_206), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_394), .Y(n_471) );
XNOR2xp5_ASAP7_75t_L g472 ( .A(n_374), .B(n_71), .Y(n_472) );
AOI222xp33_ASAP7_75t_L g473 ( .A1(n_374), .A2(n_74), .B1(n_172), .B2(n_180), .C1(n_340), .C2(n_339), .Y(n_473) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_390), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_387), .B(n_412), .Y(n_475) );
XOR2x2_ASAP7_75t_L g476 ( .A(n_374), .B(n_390), .Y(n_476) );
OAI21xp33_ASAP7_75t_SL g477 ( .A1(n_427), .A2(n_415), .B(n_436), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_429), .A2(n_414), .B1(n_473), .B2(n_415), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_448), .B(n_453), .Y(n_480) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_472), .A2(n_414), .B(n_453), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_474), .B(n_475), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g483 ( .A1(n_416), .A2(n_425), .B1(n_419), .B2(n_471), .C(n_422), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_470), .A2(n_431), .B(n_446), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_457), .B(n_439), .Y(n_485) );
XNOR2x2_ASAP7_75t_L g486 ( .A(n_476), .B(n_456), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_435), .B(n_430), .Y(n_487) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_470), .B(n_469), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_428), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_418), .A2(n_423), .B1(n_444), .B2(n_440), .C(n_459), .Y(n_490) );
XNOR2xp5_ASAP7_75t_L g491 ( .A(n_432), .B(n_462), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_450), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_442), .B(n_434), .C(n_458), .Y(n_493) );
AO22x2_ASAP7_75t_L g494 ( .A1(n_486), .A2(n_449), .B1(n_438), .B2(n_437), .Y(n_494) );
OA22x2_ASAP7_75t_L g495 ( .A1(n_478), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_495) );
OA22x2_ASAP7_75t_L g496 ( .A1(n_491), .A2(n_451), .B1(n_461), .B2(n_460), .Y(n_496) );
NOR4xp25_ASAP7_75t_L g497 ( .A(n_477), .B(n_452), .C(n_443), .D(n_447), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_479), .Y(n_498) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_481), .A2(n_454), .B(n_465), .C(n_426), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g500 ( .A1(n_481), .A2(n_441), .B(n_455), .C(n_466), .Y(n_500) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_484), .A2(n_424), .A3(n_455), .B(n_468), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_487), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_494), .A2(n_482), .B1(n_480), .B2(n_483), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_499), .B(n_492), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_502), .B(n_490), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_494), .A2(n_488), .B1(n_485), .B2(n_489), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_500), .B(n_493), .C(n_463), .Y(n_507) );
NAND5xp2_ASAP7_75t_L g508 ( .A(n_503), .B(n_501), .C(n_495), .D(n_497), .E(n_464), .Y(n_508) );
AOI22xp5_ASAP7_75t_SL g509 ( .A1(n_506), .A2(n_496), .B1(n_498), .B2(n_467), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_504), .A2(n_445), .B1(n_421), .B2(n_420), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_510), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_509), .Y(n_512) );
NOR3x2_ASAP7_75t_L g513 ( .A(n_512), .B(n_508), .C(n_507), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_513), .Y(n_514) );
XNOR2xp5_ASAP7_75t_L g515 ( .A(n_514), .B(n_511), .Y(n_515) );
NAND3x2_ASAP7_75t_L g516 ( .A(n_515), .B(n_505), .C(n_433), .Y(n_516) );
endmodule