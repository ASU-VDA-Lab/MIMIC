module fake_jpeg_10687_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_79),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_2),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_26),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_70),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_63),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_63),
.B1(n_52),
.B2(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_56),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_69),
.B(n_61),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_67),
.B1(n_65),
.B2(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_50),
.B1(n_53),
.B2(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_78),
.B1(n_60),
.B2(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_12),
.B(n_13),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_104),
.Y(n_121)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_108),
.Y(n_134)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_75),
.B1(n_56),
.B2(n_55),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_107),
.B1(n_37),
.B2(n_38),
.Y(n_135)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_113),
.B(n_31),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_115),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_48),
.B1(n_43),
.B2(n_44),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_28),
.A3(n_47),
.B1(n_46),
.B2(n_45),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_5),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_6),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_114),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_136),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_126),
.B1(n_129),
.B2(n_133),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_131),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_124),
.B(n_122),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_15),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_138),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_22),
.B(n_24),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_25),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_135),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_144),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_132),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_137),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_155),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_128),
.C(n_131),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_159),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_148),
.C(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_141),
.B1(n_158),
.B2(n_160),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_153),
.B1(n_151),
.B2(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_148),
.B1(n_155),
.B2(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_156),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_165),
.B(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_167),
.B(n_166),
.Y(n_174)
);


endmodule