module fake_jpeg_21995_n_282 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_282);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_282;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_20),
.B1(n_25),
.B2(n_21),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_31),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_18),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_40),
.B(n_18),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_24),
.C(n_32),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_38),
.C(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_62),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_58),
.B1(n_85),
.B2(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_64),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_70),
.B1(n_75),
.B2(n_47),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_67),
.B(n_73),
.Y(n_110)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_20),
.B1(n_32),
.B2(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_80),
.B(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_20),
.B1(n_27),
.B2(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_27),
.B1(n_37),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_84),
.B1(n_19),
.B2(n_30),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_50),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_48),
.Y(n_104)
);

AO22x2_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_35),
.B1(n_27),
.B2(n_30),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_30),
.B1(n_48),
.B2(n_23),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_30),
.B1(n_31),
.B2(n_22),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_19),
.B1(n_29),
.B2(n_26),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_91),
.B1(n_99),
.B2(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_47),
.B1(n_42),
.B2(n_29),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_96),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_42),
.B1(n_26),
.B2(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_97),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_107),
.B(n_71),
.Y(n_125)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_29),
.B1(n_31),
.B2(n_16),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_109),
.B1(n_112),
.B2(n_77),
.Y(n_133)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_68),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_22),
.B1(n_23),
.B2(n_7),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_61),
.B1(n_70),
.B2(n_59),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_66),
.B(n_78),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_120),
.B(n_127),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_112),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_124),
.C(n_138),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_121),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_65),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g121 ( 
.A(n_111),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_128),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_134),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_131),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_72),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_9),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_102),
.B1(n_110),
.B2(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_106),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_0),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_72),
.C(n_60),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_96),
.B1(n_103),
.B2(n_97),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_143),
.B1(n_151),
.B2(n_159),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_157),
.C(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_102),
.B1(n_88),
.B2(n_100),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_122),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_109),
.B1(n_56),
.B2(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_109),
.B1(n_86),
.B2(n_81),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_81),
.B1(n_28),
.B2(n_2),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_161),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_9),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_155),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_0),
.Y(n_155)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_28),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_127),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_28),
.C(n_1),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_28),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_159)
);

INVx13_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_0),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_137),
.B(n_128),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_9),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_177),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_195),
.B1(n_185),
.B2(n_148),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_114),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_146),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_120),
.B(n_127),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_182),
.B(n_162),
.C(n_155),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_117),
.B1(n_135),
.B2(n_121),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_185),
.A2(n_192),
.B1(n_143),
.B2(n_159),
.Y(n_196)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_129),
.B1(n_136),
.B2(n_123),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_148),
.B(n_158),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_196),
.A2(n_205),
.B1(n_207),
.B2(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_169),
.B1(n_149),
.B2(n_160),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_204),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_144),
.B1(n_141),
.B2(n_142),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_157),
.C(n_164),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_180),
.C(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_152),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_212),
.B(n_170),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_150),
.A3(n_162),
.B1(n_163),
.B2(n_155),
.C1(n_154),
.C2(n_10),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_203),
.B1(n_209),
.B2(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_226),
.Y(n_239)
);

NAND2x1p5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_225),
.C(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_175),
.B(n_183),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_173),
.C(n_179),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_178),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_230),
.B1(n_231),
.B2(n_190),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_177),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_202),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.C(n_176),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_192),
.C(n_196),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_243),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_210),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_223),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_220),
.B(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.C(n_251),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_224),
.B(n_220),
.Y(n_247)
);

AOI221xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_219),
.B1(n_216),
.B2(n_215),
.C(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_254),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_215),
.B1(n_218),
.B2(n_186),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_253),
.B1(n_244),
.B2(n_170),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_201),
.B(n_218),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_201),
.B1(n_176),
.B2(n_187),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_260),
.Y(n_269)
);

BUFx4f_ASAP7_75t_SL g258 ( 
.A(n_246),
.Y(n_258)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_242),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_10),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_255),
.A3(n_10),
.B1(n_4),
.B2(n_6),
.C1(n_8),
.C2(n_14),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_3),
.C(n_6),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_254),
.B(n_245),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_259),
.B(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_267),
.B(n_265),
.C(n_270),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_3),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

O2A1O1Ixp33_ASAP7_75t_SL g279 ( 
.A1(n_277),
.A2(n_267),
.B(n_271),
.C(n_269),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_279),
.A2(n_264),
.B1(n_12),
.B2(n_14),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_280),
.A2(n_278),
.B1(n_11),
.B2(n_12),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_11),
.B(n_12),
.Y(n_282)
);


endmodule