module real_jpeg_27970_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_326, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_326;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_0),
.A2(n_42),
.B1(n_62),
.B2(n_63),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_0),
.A2(n_42),
.B1(n_53),
.B2(n_55),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_1),
.A2(n_53),
.B1(n_55),
.B2(n_73),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_53),
.B1(n_55),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_107),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_107),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_107),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_53),
.Y(n_78)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_53),
.B1(n_55),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_4),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_86),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_86),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_86),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_5),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_40),
.B1(n_53),
.B2(n_55),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_47),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_9),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_53),
.B1(n_55),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_128),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_128),
.Y(n_296)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_32),
.B(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_12),
.B(n_67),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_12),
.A2(n_35),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_12),
.B(n_93),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_12),
.A2(n_82),
.B1(n_104),
.B2(n_174),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_12),
.A2(n_31),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_53),
.B1(n_55),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_13),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_80),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_80),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_278)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_305),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_273),
.A3(n_300),
.B1(n_303),
.B2(n_304),
.C(n_325),
.Y(n_19)
);

AOI321xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_224),
.A3(n_262),
.B1(n_267),
.B2(n_272),
.C(n_326),
.Y(n_20)
);

NOR3xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_120),
.C(n_139),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_97),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_23),
.B(n_97),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_74),
.C(n_87),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_24),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_60),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_26),
.B(n_44),
.C(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_27)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_28),
.A2(n_34),
.B1(n_41),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_28),
.A2(n_34),
.B1(n_91),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_28),
.A2(n_34),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_28),
.A2(n_34),
.B(n_313),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_29),
.A2(n_31),
.A3(n_36),
.B1(n_190),
.B2(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_31),
.A2(n_32),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_32),
.B(n_70),
.Y(n_190)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g151 ( 
.A1(n_35),
.A2(n_51),
.A3(n_55),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_35),
.B(n_37),
.Y(n_198)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_39),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_57),
.B2(n_59),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_48),
.A2(n_59),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_48),
.A2(n_59),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_50),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_49),
.A2(n_50),
.B1(n_102),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_50),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_49),
.A2(n_50),
.B1(n_149),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_49),
.A2(n_50),
.B1(n_237),
.B2(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_49),
.A2(n_50),
.B(n_249),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_50),
.B(n_70),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_52),
.B(n_53),
.Y(n_153)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_53),
.B(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_60)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_67),
.B1(n_115),
.B2(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_61),
.A2(n_67),
.B1(n_135),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_61),
.A2(n_67),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B(n_66),
.C(n_67),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_65),
.Y(n_66)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_68),
.B(n_70),
.C(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_70),
.B(n_82),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_72),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_74),
.A2(n_87),
.B1(n_88),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_85),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_78),
.A2(n_81),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_104),
.B1(n_106),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_82),
.A2(n_104),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_82),
.A2(n_104),
.B1(n_168),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_82),
.A2(n_104),
.B1(n_163),
.B2(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_82),
.A2(n_104),
.B(n_127),
.Y(n_239)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_96),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_89),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_93),
.B1(n_118),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_92),
.A2(n_93),
.B1(n_137),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_92),
.A2(n_93),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_92),
.A2(n_93),
.B1(n_282),
.B2(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_94),
.B(n_96),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_95),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_108),
.C(n_109),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_103),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_116),
.C(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_112),
.A2(n_113),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_112),
.A2(n_113),
.B1(n_256),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_112),
.A2(n_113),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_121),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_122),
.B(n_123),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_138),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_125),
.B(n_131),
.C(n_138),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_126),
.B(n_129),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_130),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_132),
.B(n_134),
.C(n_136),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_218),
.B(n_223),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_204),
.B(n_217),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_183),
.B(n_203),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_164),
.B(n_182),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_146),
.B1(n_150),
.B2(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_160),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_181),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_170),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_176),
.B(n_180),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_185),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_196),
.B1(n_201),
.B2(n_202),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_195),
.C(n_202),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_199),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_241),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_241),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.C(n_240),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_232),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_226),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.CI(n_231),
.CON(n_226),
.SN(n_226)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_229),
.C(n_231),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_230),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_239),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_238),
.A2(n_254),
.B(n_257),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_260),
.B2(n_261),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_251),
.C(n_261),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_248),
.B(n_250),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_248),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_275),
.C(n_287),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_250),
.B(n_275),
.CI(n_287),
.CON(n_302),
.SN(n_302)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_268),
.B(n_271),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_288),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_288),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_286),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_277),
.B1(n_290),
.B2(n_298),
.Y(n_289)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_280),
.C(n_285),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_298),
.C(n_299),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_285),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_291),
.C(n_295),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_299),
.Y(n_288)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_302),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_302),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_320),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_318),
.B2(n_319),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_314),
.B2(n_315),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);


endmodule