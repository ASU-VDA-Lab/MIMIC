module fake_jpeg_4512_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_20),
.B1(n_33),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_51),
.B1(n_55),
.B2(n_18),
.Y(n_86)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_33),
.B1(n_20),
.B2(n_32),
.Y(n_51)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_18),
.B1(n_27),
.B2(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_23),
.Y(n_77)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_16),
.B1(n_31),
.B2(n_24),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_10),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_20),
.B1(n_43),
.B2(n_23),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_83),
.B1(n_69),
.B2(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_69),
.B1(n_53),
.B2(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_97),
.Y(n_125)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_79),
.B1(n_90),
.B2(n_92),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_34),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_101),
.B(n_108),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_61),
.B(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_34),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_115),
.B1(n_117),
.B2(n_90),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_54),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_119),
.B(n_105),
.C(n_107),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_85),
.B1(n_93),
.B2(n_76),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_34),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_58),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_34),
.C(n_39),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_53),
.B1(n_56),
.B2(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_28),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_111),
.B1(n_117),
.B2(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_82),
.B1(n_70),
.B2(n_78),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_129),
.B1(n_130),
.B2(n_135),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_39),
.CI(n_36),
.CON(n_128),
.SN(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_145),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_85),
.B1(n_76),
.B2(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_85),
.B1(n_73),
.B2(n_26),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_136),
.B1(n_143),
.B2(n_111),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_115),
.C(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_52),
.B1(n_27),
.B2(n_26),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_28),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_114),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_27),
.B1(n_25),
.B2(n_21),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_79),
.B1(n_39),
.B2(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_96),
.A2(n_39),
.B1(n_92),
.B2(n_90),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_155),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_100),
.B1(n_102),
.B2(n_112),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_163),
.B1(n_173),
.B2(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_100),
.C(n_134),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_132),
.B1(n_126),
.B2(n_138),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_161),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_101),
.B(n_118),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_160),
.B(n_136),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_102),
.B(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_167),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_131),
.B(n_116),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_133),
.C(n_143),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_111),
.B1(n_106),
.B2(n_112),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_178),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_150),
.C(n_152),
.Y(n_178)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_183),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_192),
.B(n_169),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_151),
.B(n_164),
.Y(n_207)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_191),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_129),
.B1(n_144),
.B2(n_132),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_197),
.B1(n_200),
.B2(n_164),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_29),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_125),
.C(n_126),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_138),
.B(n_97),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_137),
.B1(n_139),
.B2(n_39),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_174),
.B1(n_25),
.B2(n_29),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_155),
.B(n_37),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_208),
.B1(n_216),
.B2(n_221),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_206),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_225),
.C(n_176),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_159),
.B1(n_156),
.B2(n_161),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_205),
.A2(n_209),
.B1(n_213),
.B2(n_187),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_177),
.B1(n_29),
.B2(n_17),
.Y(n_242)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_159),
.B(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_190),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_17),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

OAI31xp33_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_163),
.A3(n_29),
.B(n_17),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_217),
.A2(n_219),
.B1(n_197),
.B2(n_188),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_196),
.B(n_198),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_223),
.B1(n_17),
.B2(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_29),
.Y(n_222)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_199),
.A2(n_37),
.B(n_36),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_182),
.B(n_184),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_231),
.B(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_234),
.C(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_178),
.C(n_194),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_181),
.C(n_175),
.Y(n_237)
);

XOR2x2_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_175),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_207),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_242),
.B1(n_223),
.B2(n_210),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_200),
.C(n_187),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_17),
.C(n_2),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_256),
.B1(n_238),
.B2(n_239),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_255),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_259),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_213),
.B1(n_209),
.B2(n_219),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_233),
.B1(n_235),
.B2(n_245),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_228),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_225),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_220),
.B1(n_208),
.B2(n_201),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_222),
.C(n_212),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.C(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_1),
.C(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_15),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_261),
.B(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_273),
.C(n_6),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_270),
.B1(n_274),
.B2(n_277),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_248),
.A2(n_232),
.B1(n_243),
.B2(n_4),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_278),
.B1(n_262),
.B2(n_260),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_271),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_1),
.C(n_3),
.Y(n_273)
);

NAND2x1_ASAP7_75t_SL g274 ( 
.A(n_253),
.B(n_3),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_13),
.B(n_15),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_11),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_278),
.Y(n_282)
);

OAI221xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_259),
.B1(n_257),
.B2(n_255),
.C(n_254),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_12),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_249),
.B1(n_11),
.B2(n_10),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_249),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_282),
.C(n_287),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_8),
.B1(n_290),
.B2(n_287),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_7),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_6),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_289),
.B(n_7),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_282),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_286),
.A2(n_264),
.B(n_273),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_293),
.B(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

INVx11_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_268),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_301),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_281),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_299),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_8),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_292),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_303),
.C(n_308),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_302),
.B(n_309),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_317),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_305),
.Y(n_320)
);


endmodule