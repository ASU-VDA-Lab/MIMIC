module real_aes_7430_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_85), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g447 ( .A(n_0), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_1), .A2(n_140), .B(n_143), .C(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_2), .A2(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g499 ( .A(n_3), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_4), .B(n_179), .Y(n_178) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_5), .A2(n_168), .B(n_477), .Y(n_476) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g243 ( .A(n_7), .Y(n_243) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_8), .B(n_40), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_9), .A2(n_267), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_10), .B(n_152), .Y(n_220) );
INVx1_ASAP7_75t_L g481 ( .A(n_11), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_12), .B(n_173), .Y(n_532) );
INVx1_ASAP7_75t_L g132 ( .A(n_13), .Y(n_132) );
INVx1_ASAP7_75t_L g544 ( .A(n_14), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_15), .A2(n_187), .B(n_228), .C(n_230), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_16), .B(n_179), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_17), .B(n_470), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_18), .B(n_168), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_19), .B(n_275), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_173), .B(n_204), .C(n_207), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_21), .B(n_179), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_22), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_23), .A2(n_206), .B(n_230), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_24), .B(n_152), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_25), .Y(n_134) );
INVx1_ASAP7_75t_L g185 ( .A(n_26), .Y(n_185) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_28), .Y(n_216) );
AOI222xp33_ASAP7_75t_L g451 ( .A1(n_29), .A2(n_43), .B1(n_452), .B2(n_740), .C1(n_741), .C2(n_744), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_30), .B(n_152), .Y(n_500) );
INVx1_ASAP7_75t_L g272 ( .A(n_31), .Y(n_272) );
INVx1_ASAP7_75t_L g489 ( .A(n_32), .Y(n_489) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_34), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_35), .A2(n_173), .B(n_174), .C(n_176), .Y(n_172) );
INVxp67_ASAP7_75t_L g273 ( .A(n_36), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g170 ( .A(n_37), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_38), .A2(n_143), .B(n_184), .C(n_191), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_39), .A2(n_140), .B(n_143), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_40), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g488 ( .A(n_41), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_42), .A2(n_118), .B1(n_439), .B2(n_440), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_42), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_43), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_44), .A2(n_154), .B(n_241), .C(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_45), .B(n_152), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_47), .Y(n_269) );
INVx1_ASAP7_75t_L g202 ( .A(n_48), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_49), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_50), .B(n_168), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_51), .A2(n_143), .B1(n_207), .B2(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_52), .Y(n_515) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_53), .Y(n_496) );
CKINVDCx14_ASAP7_75t_R g239 ( .A(n_54), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_55), .A2(n_176), .B(n_241), .C(n_480), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_56), .Y(n_524) );
INVx1_ASAP7_75t_L g478 ( .A(n_57), .Y(n_478) );
INVx1_ASAP7_75t_L g141 ( .A(n_58), .Y(n_141) );
INVx1_ASAP7_75t_L g131 ( .A(n_59), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_60), .A2(n_100), .B1(n_111), .B2(n_748), .Y(n_99) );
INVx1_ASAP7_75t_SL g175 ( .A(n_61), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_62), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_63), .B(n_179), .Y(n_209) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_SL g469 ( .A1(n_65), .A2(n_176), .B(n_470), .C(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_L g472 ( .A(n_66), .Y(n_472) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_68), .A2(n_168), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_69), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_70), .A2(n_168), .B(n_225), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_71), .Y(n_492) );
INVx1_ASAP7_75t_L g518 ( .A(n_72), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_73), .B(n_443), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_74), .A2(n_267), .B(n_268), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_75), .Y(n_182) );
INVx1_ASAP7_75t_L g226 ( .A(n_76), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_77), .A2(n_140), .B(n_143), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_78), .A2(n_168), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g229 ( .A(n_79), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_80), .B(n_186), .Y(n_512) );
INVx2_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
INVx1_ASAP7_75t_L g219 ( .A(n_82), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_83), .B(n_470), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_84), .A2(n_140), .B(n_143), .C(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g444 ( .A(n_85), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g456 ( .A(n_85), .Y(n_456) );
OR2x2_ASAP7_75t_L g739 ( .A(n_85), .B(n_446), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_86), .A2(n_143), .B(n_146), .C(n_156), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_87), .B(n_161), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_88), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_89), .A2(n_140), .B(n_143), .C(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_90), .Y(n_536) );
INVx1_ASAP7_75t_L g468 ( .A(n_91), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_92), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_93), .B(n_186), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_94), .B(n_127), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_95), .B(n_127), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g205 ( .A(n_97), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_98), .A2(n_168), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_103), .Y(n_749) );
CKINVDCx9p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_450), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g747 ( .A(n_113), .Y(n_747) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_441), .B(n_449), .Y(n_116) );
INVx3_ASAP7_75t_L g440 ( .A(n_118), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_118), .A2(n_454), .B1(n_738), .B2(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_SL g118 ( .A(n_119), .B(n_394), .Y(n_118) );
NOR4xp25_ASAP7_75t_L g119 ( .A(n_120), .B(n_331), .C(n_365), .D(n_381), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_257), .C(n_295), .D(n_311), .Y(n_120) );
AOI222xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_194), .B1(n_232), .B2(n_245), .C1(n_250), .C2(n_256), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI31xp33_ASAP7_75t_L g427 ( .A1(n_123), .A2(n_428), .A3(n_429), .B(n_431), .Y(n_427) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_162), .Y(n_123) );
AND2x2_ASAP7_75t_L g402 ( .A(n_124), .B(n_164), .Y(n_402) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_SL g249 ( .A(n_125), .Y(n_249) );
AND2x2_ASAP7_75t_L g256 ( .A(n_125), .B(n_180), .Y(n_256) );
AND2x2_ASAP7_75t_L g316 ( .A(n_125), .B(n_165), .Y(n_316) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
INVx3_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_126), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g514 ( .A(n_126), .B(n_515), .Y(n_514) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_127), .A2(n_466), .B(n_473), .Y(n_465) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g265 ( .A(n_128), .Y(n_265) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_129), .B(n_130), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_142), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_135), .A2(n_161), .B(n_182), .C(n_183), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_135), .A2(n_216), .B(n_217), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_135), .A2(n_157), .B1(n_486), .B2(n_490), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_135), .A2(n_496), .B(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_135), .A2(n_518), .B(n_519), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g168 ( .A(n_136), .B(n_140), .Y(n_168) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g208 ( .A(n_138), .Y(n_208) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
INVx3_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g470 ( .A(n_139), .Y(n_470) );
INVx4_ASAP7_75t_SL g157 ( .A(n_140), .Y(n_157) );
BUFx3_ASAP7_75t_L g191 ( .A(n_140), .Y(n_191) );
INVx5_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_151), .C(n_153), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_148), .A2(n_153), .B(n_219), .C(n_220), .Y(n_218) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_149), .A2(n_150), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
INVx4_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
INVx2_ASAP7_75t_L g241 ( .A(n_152), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_153), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_153), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_157), .A2(n_170), .B(n_171), .C(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g201 ( .A1(n_157), .A2(n_171), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_SL g225 ( .A1(n_157), .A2(n_171), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_157), .A2(n_171), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g268 ( .A1(n_157), .A2(n_171), .B(n_269), .C(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_157), .A2(n_171), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_157), .A2(n_171), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_157), .A2(n_171), .B(n_541), .C(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx1_ASAP7_75t_L g275 ( .A(n_160), .Y(n_275) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_160), .A2(n_528), .B(n_535), .Y(n_527) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g214 ( .A(n_161), .Y(n_214) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_161), .A2(n_237), .B(n_244), .Y(n_236) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_539), .B(n_545), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_162), .B(n_346), .Y(n_345) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_163), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_163), .B(n_260), .Y(n_306) );
AND2x2_ASAP7_75t_L g399 ( .A(n_163), .B(n_339), .Y(n_399) );
OAI321xp33_ASAP7_75t_L g433 ( .A1(n_163), .A2(n_249), .A3(n_406), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_163), .B(n_235), .C(n_346), .D(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
AND2x2_ASAP7_75t_L g301 ( .A(n_164), .B(n_247), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_164), .B(n_249), .Y(n_320) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g248 ( .A(n_165), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g276 ( .A(n_165), .B(n_180), .Y(n_276) );
AND2x2_ASAP7_75t_L g362 ( .A(n_165), .B(n_247), .Y(n_362) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_178), .Y(n_165) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_200), .B(n_209), .Y(n_199) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_224), .B(n_231), .Y(n_223) );
BUFx2_ASAP7_75t_L g267 ( .A(n_168), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_173), .B(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_177), .Y(n_533) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_179), .A2(n_476), .B(n_482), .Y(n_475) );
INVx3_ASAP7_75t_SL g247 ( .A(n_180), .Y(n_247) );
AND2x2_ASAP7_75t_L g294 ( .A(n_180), .B(n_281), .Y(n_294) );
OR2x2_ASAP7_75t_L g327 ( .A(n_180), .B(n_249), .Y(n_327) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_180), .Y(n_334) );
AND2x2_ASAP7_75t_L g363 ( .A(n_180), .B(n_248), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_180), .B(n_336), .Y(n_378) );
AND2x2_ASAP7_75t_L g410 ( .A(n_180), .B(n_402), .Y(n_410) );
AND2x2_ASAP7_75t_L g419 ( .A(n_180), .B(n_261), .Y(n_419) );
OR2x6_ASAP7_75t_L g180 ( .A(n_181), .B(n_192), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_189), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_186), .A2(n_206), .B1(n_272), .B2(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_186), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
INVx5_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_187), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_187), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_187), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_190), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_210), .Y(n_195) );
INVx1_ASAP7_75t_SL g387 ( .A(n_196), .Y(n_387) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g252 ( .A(n_197), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g234 ( .A(n_198), .B(n_212), .Y(n_234) );
AND2x2_ASAP7_75t_L g323 ( .A(n_198), .B(n_236), .Y(n_323) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g293 ( .A(n_199), .B(n_223), .Y(n_293) );
OR2x2_ASAP7_75t_L g304 ( .A(n_199), .B(n_236), .Y(n_304) );
AND2x2_ASAP7_75t_L g330 ( .A(n_199), .B(n_236), .Y(n_330) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_199), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_206), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_206), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g501 ( .A(n_207), .Y(n_501) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_210), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_210), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g303 ( .A(n_211), .B(n_304), .Y(n_303) );
AOI322xp5_ASAP7_75t_L g389 ( .A1(n_211), .A2(n_293), .A3(n_299), .B1(n_330), .B2(n_380), .C1(n_390), .C2(n_392), .Y(n_389) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_212), .B(n_235), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_212), .B(n_236), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_212), .B(n_253), .Y(n_310) );
AND2x2_ASAP7_75t_L g364 ( .A(n_212), .B(n_330), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_212), .Y(n_368) );
AND2x2_ASAP7_75t_L g380 ( .A(n_212), .B(n_223), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_212), .B(n_252), .Y(n_412) );
INVx4_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g277 ( .A(n_213), .B(n_223), .Y(n_277) );
BUFx3_ASAP7_75t_L g291 ( .A(n_213), .Y(n_291) );
AND3x2_ASAP7_75t_L g373 ( .A(n_213), .B(n_353), .C(n_374), .Y(n_373) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_214), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_214), .B(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_214), .B(n_536), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g233 ( .A(n_223), .B(n_234), .C(n_235), .Y(n_233) );
INVx1_ASAP7_75t_SL g253 ( .A(n_223), .Y(n_253) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_223), .Y(n_358) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g352 ( .A(n_234), .B(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g359 ( .A(n_234), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_235), .B(n_375), .Y(n_397) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
BUFx3_ASAP7_75t_L g278 ( .A(n_236), .Y(n_278) );
AND2x2_ASAP7_75t_L g353 ( .A(n_236), .B(n_253), .Y(n_353) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
OR2x2_ASAP7_75t_L g297 ( .A(n_247), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g416 ( .A(n_247), .B(n_316), .Y(n_416) );
AND2x2_ASAP7_75t_L g430 ( .A(n_247), .B(n_249), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_248), .B(n_261), .Y(n_371) );
AND2x2_ASAP7_75t_L g418 ( .A(n_248), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g281 ( .A(n_249), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g298 ( .A(n_249), .B(n_261), .Y(n_298) );
INVx1_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
AND2x2_ASAP7_75t_L g339 ( .A(n_249), .B(n_261), .Y(n_339) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI221xp5_ASAP7_75t_L g381 ( .A1(n_251), .A2(n_382), .B1(n_386), .B2(n_388), .C(n_389), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g285 ( .A(n_252), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_255), .B(n_292), .Y(n_435) );
AOI322xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_277), .A3(n_278), .B1(n_279), .B2(n_285), .C1(n_287), .C2(n_294), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_276), .Y(n_259) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_260), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_260), .B(n_326), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_260), .A2(n_276), .B(n_350), .C(n_351), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_260), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_260), .B(n_320), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_260), .B(n_402), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_260), .B(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_261), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_261), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g391 ( .A(n_261), .B(n_278), .Y(n_391) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_266), .B(n_274), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_263), .A2(n_283), .B(n_284), .Y(n_282) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_263), .A2(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_SL g508 ( .A1(n_264), .A2(n_509), .B(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_265), .A2(n_485), .B(n_491), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_265), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_265), .A2(n_495), .B(n_502), .Y(n_494) );
INVx1_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_274), .Y(n_284) );
INVx1_ASAP7_75t_L g366 ( .A(n_276), .Y(n_366) );
OAI31xp33_ASAP7_75t_L g376 ( .A1(n_276), .A2(n_301), .A3(n_377), .B(n_379), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_276), .B(n_282), .Y(n_428) );
INVx1_ASAP7_75t_SL g289 ( .A(n_277), .Y(n_289) );
AND2x2_ASAP7_75t_L g322 ( .A(n_277), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g403 ( .A(n_277), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g288 ( .A(n_278), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g313 ( .A(n_278), .Y(n_313) );
AND2x2_ASAP7_75t_L g340 ( .A(n_278), .B(n_293), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_278), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g432 ( .A(n_278), .B(n_380), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_280), .B(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g337 ( .A(n_282), .Y(n_337) );
NAND2xp33_ASAP7_75t_SL g287 ( .A(n_288), .B(n_290), .Y(n_287) );
OAI211xp5_ASAP7_75t_SL g331 ( .A1(n_289), .A2(n_332), .B(n_338), .C(n_354), .Y(n_331) );
OR2x2_ASAP7_75t_L g406 ( .A(n_289), .B(n_387), .Y(n_406) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g343 ( .A(n_291), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_291), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_313), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B(n_302), .C(n_305), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g346 ( .A(n_298), .Y(n_346) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_301), .B(n_339), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_301), .Y(n_350) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g309 ( .A(n_304), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g342 ( .A(n_304), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
AOI21xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_307), .B(n_309), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_307), .A2(n_318), .B(n_321), .Y(n_317) );
AOI211xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B(n_317), .C(n_324), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_312), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_315), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_SL g328 ( .A(n_316), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_318), .A2(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_323), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g348 ( .A(n_323), .Y(n_348) );
AOI21xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_328), .B(n_329), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_336), .B(n_362), .Y(n_388) );
AND2x2_ASAP7_75t_L g401 ( .A(n_336), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g415 ( .A(n_336), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g425 ( .A(n_336), .B(n_363), .Y(n_425) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI211xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_341), .C(n_349), .Y(n_338) );
INVx1_ASAP7_75t_L g385 ( .A(n_339), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_345), .B2(n_347), .Y(n_341) );
OR2x2_ASAP7_75t_L g347 ( .A(n_343), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_343), .B(n_404), .Y(n_426) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g420 ( .A(n_353), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B1(n_363), .B2(n_364), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g438 ( .A(n_358), .Y(n_438) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_369), .C(n_376), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_384), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR5xp2_ASAP7_75t_L g394 ( .A(n_395), .B(n_413), .C(n_421), .D(n_427), .E(n_433), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_398), .B(n_400), .C(n_407), .Y(n_395) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_405), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_410), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_420), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g436 ( .A(n_416), .Y(n_436) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_440), .A2(n_454), .B1(n_457), .B2(n_738), .Y(n_453) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_445), .B(n_456), .Y(n_743) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g455 ( .A(n_446), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AOI21xp33_ASAP7_75t_L g450 ( .A1(n_449), .A2(n_451), .B(n_747), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g746 ( .A(n_457), .Y(n_746) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND4x1_ASAP7_75t_L g458 ( .A(n_459), .B(n_656), .C(n_703), .D(n_723), .Y(n_458) );
NOR3xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_586), .C(n_611), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_504), .B(n_546), .C(n_576), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_483), .Y(n_462) );
INVx3_ASAP7_75t_SL g628 ( .A(n_463), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_463), .B(n_559), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_463), .B(n_493), .Y(n_709) );
AND2x2_ASAP7_75t_L g732 ( .A(n_463), .B(n_598), .Y(n_732) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g550 ( .A(n_465), .B(n_475), .Y(n_550) );
INVx3_ASAP7_75t_L g563 ( .A(n_465), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_465), .B(n_474), .Y(n_568) );
OR2x2_ASAP7_75t_L g619 ( .A(n_465), .B(n_560), .Y(n_619) );
BUFx2_ASAP7_75t_L g639 ( .A(n_465), .Y(n_639) );
AND2x2_ASAP7_75t_L g649 ( .A(n_465), .B(n_560), .Y(n_649) );
AND2x2_ASAP7_75t_L g655 ( .A(n_465), .B(n_484), .Y(n_655) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_475), .B(n_560), .Y(n_574) );
INVx2_ASAP7_75t_L g584 ( .A(n_475), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_475), .B(n_563), .Y(n_597) );
OR2x2_ASAP7_75t_L g608 ( .A(n_475), .B(n_560), .Y(n_608) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_475), .B(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g666 ( .A(n_475), .Y(n_666) );
AND2x2_ASAP7_75t_L g712 ( .A(n_475), .B(n_484), .Y(n_712) );
INVx3_ASAP7_75t_SL g585 ( .A(n_483), .Y(n_585) );
OR2x2_ASAP7_75t_L g638 ( .A(n_483), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
INVx3_ASAP7_75t_L g560 ( .A(n_484), .Y(n_560) );
AND2x2_ASAP7_75t_L g627 ( .A(n_484), .B(n_494), .Y(n_627) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_484), .Y(n_695) );
AOI33xp33_ASAP7_75t_L g699 ( .A1(n_484), .A2(n_628), .A3(n_635), .B1(n_644), .B2(n_700), .B3(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g548 ( .A(n_493), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_493), .B(n_563), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_493), .B(n_623), .C(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g648 ( .A(n_493), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_493), .B(n_655), .Y(n_658) );
AND2x2_ASAP7_75t_L g711 ( .A(n_493), .B(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g567 ( .A(n_494), .Y(n_567) );
OR2x2_ASAP7_75t_L g661 ( .A(n_494), .B(n_560), .Y(n_661) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_525), .Y(n_504) );
AOI32xp33_ASAP7_75t_L g612 ( .A1(n_505), .A2(n_613), .A3(n_615), .B1(n_617), .B2(n_620), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_505), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g715 ( .A(n_505), .Y(n_715) );
INVx4_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g647 ( .A(n_506), .B(n_631), .Y(n_647) );
AND2x2_ASAP7_75t_L g667 ( .A(n_506), .B(n_593), .Y(n_667) );
AND2x2_ASAP7_75t_L g735 ( .A(n_506), .B(n_653), .Y(n_735) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
INVx3_ASAP7_75t_L g556 ( .A(n_507), .Y(n_556) );
AND2x2_ASAP7_75t_L g570 ( .A(n_507), .B(n_554), .Y(n_570) );
OR2x2_ASAP7_75t_L g575 ( .A(n_507), .B(n_553), .Y(n_575) );
INVx1_ASAP7_75t_L g582 ( .A(n_507), .Y(n_582) );
AND2x2_ASAP7_75t_L g590 ( .A(n_507), .B(n_564), .Y(n_590) );
AND2x2_ASAP7_75t_L g592 ( .A(n_507), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_507), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g645 ( .A(n_507), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_507), .B(n_730), .Y(n_729) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx2_ASAP7_75t_L g554 ( .A(n_516), .Y(n_554) );
AND2x2_ASAP7_75t_L g600 ( .A(n_516), .B(n_526), .Y(n_600) );
AND2x2_ASAP7_75t_L g610 ( .A(n_516), .B(n_538), .Y(n_610) );
INVx2_ASAP7_75t_L g730 ( .A(n_525), .Y(n_730) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_526), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
AND2x2_ASAP7_75t_L g615 ( .A(n_526), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g631 ( .A(n_526), .B(n_594), .Y(n_631) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g579 ( .A(n_527), .Y(n_579) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g644 ( .A(n_527), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_527), .B(n_554), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g555 ( .A(n_537), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g616 ( .A(n_537), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_537), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g653 ( .A(n_537), .Y(n_653) );
INVx1_ASAP7_75t_L g686 ( .A(n_537), .Y(n_686) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g564 ( .A(n_538), .B(n_554), .Y(n_564) );
INVx1_ASAP7_75t_L g594 ( .A(n_538), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_551), .B1(n_557), .B2(n_564), .C(n_565), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_548), .B(n_568), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_548), .B(n_631), .Y(n_708) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_550), .B(n_598), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_550), .B(n_559), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_550), .B(n_573), .Y(n_702) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g624 ( .A(n_554), .Y(n_624) );
AND2x2_ASAP7_75t_L g599 ( .A(n_555), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g677 ( .A(n_555), .Y(n_677) );
AND2x2_ASAP7_75t_L g609 ( .A(n_556), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_556), .B(n_579), .Y(n_625) );
AND2x2_ASAP7_75t_L g689 ( .A(n_556), .B(n_615), .Y(n_689) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g598 ( .A(n_560), .B(n_567), .Y(n_598) );
AND2x2_ASAP7_75t_L g694 ( .A(n_561), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_563), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_564), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_564), .B(n_571), .Y(n_659) );
AND2x2_ASAP7_75t_L g679 ( .A(n_564), .B(n_579), .Y(n_679) );
AND2x2_ASAP7_75t_L g700 ( .A(n_564), .B(n_644), .Y(n_700) );
OAI32xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .A3(n_571), .B1(n_572), .B2(n_575), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_SL g573 ( .A(n_567), .Y(n_573) );
NAND2x1_ASAP7_75t_L g614 ( .A(n_567), .B(n_597), .Y(n_614) );
OR2x2_ASAP7_75t_L g618 ( .A(n_567), .B(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_567), .B(n_666), .Y(n_719) );
INVx1_ASAP7_75t_L g587 ( .A(n_568), .Y(n_587) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_569), .A2(n_660), .B1(n_706), .B2(n_709), .C(n_710), .Y(n_705) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g577 ( .A(n_570), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g620 ( .A(n_570), .B(n_593), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_570), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g698 ( .A(n_570), .B(n_631), .Y(n_698) );
INVxp67_ASAP7_75t_L g634 ( .A(n_571), .Y(n_634) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g704 ( .A(n_573), .B(n_691), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_573), .B(n_654), .Y(n_727) );
INVx1_ASAP7_75t_L g602 ( .A(n_575), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_575), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g720 ( .A(n_575), .B(n_721), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_580), .B(n_583), .Y(n_576) );
AND2x2_ASAP7_75t_L g589 ( .A(n_578), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g673 ( .A(n_582), .B(n_593), .Y(n_673) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND2x2_ASAP7_75t_L g691 ( .A(n_584), .B(n_649), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_584), .B(n_648), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_585), .B(n_597), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_591), .C(n_601), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_587), .A2(n_622), .B1(n_626), .B2(n_629), .C(n_632), .Y(n_621) );
AOI31xp33_ASAP7_75t_L g716 ( .A1(n_587), .A2(n_717), .A3(n_718), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_595), .B1(n_597), .B2(n_599), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g717 ( .A(n_597), .Y(n_717) );
INVx1_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_L g723 ( .A1(n_600), .A2(n_724), .B(n_726), .C(n_728), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_605), .B2(n_609), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_606), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_SL g696 ( .A1(n_608), .A2(n_642), .B1(n_661), .B2(n_697), .C(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g692 ( .A(n_609), .Y(n_692) );
INVx1_ASAP7_75t_L g646 ( .A(n_610), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_621), .C(n_636), .Y(n_611) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_613), .A2(n_663), .B(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_615), .B(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g722 ( .A(n_616), .Y(n_722) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g660 ( .A(n_623), .B(n_643), .Y(n_660) );
INVx1_ASAP7_75t_L g635 ( .A(n_624), .Y(n_635) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g633 ( .A(n_627), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_627), .B(n_665), .Y(n_664) );
NOR4xp25_ASAP7_75t_L g632 ( .A(n_628), .B(n_633), .C(n_634), .D(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B1(n_647), .B2(n_648), .C1(n_650), .C2(n_654), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g734 ( .A(n_638), .Y(n_734) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_650), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g710 ( .A1(n_655), .A2(n_711), .B(n_713), .Y(n_710) );
NOR4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_668), .C(n_681), .D(n_696), .Y(n_656) );
OAI221xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B1(n_660), .B2(n_661), .C(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g737 ( .A(n_658), .Y(n_737) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_665), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
OAI222xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_674), .B2(n_675), .C1(n_678), .C2(n_680), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_673), .A2(n_704), .B(n_705), .C(n_716), .Y(n_703) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
OAI222xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_687), .B1(n_688), .B2(n_690), .C1(n_692), .C2(n_693), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_698), .A2(n_701), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI211xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_731), .B(n_733), .C(n_736), .Y(n_728) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
endmodule