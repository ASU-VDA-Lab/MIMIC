module fake_jpeg_1837_n_680 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g228 ( 
.A(n_63),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_30),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_68),
.B(n_70),
.Y(n_140)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_71),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_76),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_82),
.Y(n_185)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_111),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_91),
.Y(n_209)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

BUFx12f_ASAP7_75t_SL g93 ( 
.A(n_20),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_93),
.B(n_40),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_20),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_96),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_97),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_0),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_20),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_43),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_46),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_129),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_21),
.B(n_1),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_29),
.B(n_2),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_58),
.Y(n_161)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_123),
.Y(n_222)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_37),
.Y(n_124)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx11_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_21),
.B(n_18),
.Y(n_129)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_29),
.Y(n_130)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_27),
.B(n_28),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_131),
.B(n_59),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_68),
.B(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_132),
.B(n_147),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_44),
.B1(n_26),
.B2(n_25),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_135),
.A2(n_152),
.B1(n_190),
.B2(n_15),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_27),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_78),
.A2(n_44),
.B1(n_26),
.B2(n_25),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_161),
.B(n_167),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_28),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_169),
.A2(n_194),
.B(n_199),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_118),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_170),
.B(n_184),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_114),
.A2(n_49),
.B1(n_38),
.B2(n_53),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_183),
.A2(n_211),
.B1(n_224),
.B2(n_57),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_38),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_126),
.A2(n_51),
.B1(n_43),
.B2(n_53),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_187),
.B(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_100),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_64),
.Y(n_192)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_51),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_196),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_49),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_76),
.B(n_59),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_77),
.B(n_59),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_214),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_81),
.A2(n_48),
.B1(n_52),
.B2(n_40),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_86),
.B(n_48),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_87),
.B(n_48),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_215),
.B(n_221),
.Y(n_263)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_88),
.Y(n_216)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_95),
.Y(n_217)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_98),
.B(n_52),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_63),
.B(n_52),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_223),
.B(n_4),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_104),
.A2(n_36),
.B1(n_40),
.B2(n_54),
.Y(n_224)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_61),
.Y(n_227)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_230),
.B(n_238),
.Y(n_316)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_164),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_231),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_137),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_232),
.B(n_257),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_45),
.B1(n_54),
.B2(n_57),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_235),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_236),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_237),
.B(n_245),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_138),
.B(n_2),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_137),
.B(n_3),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g355 ( 
.A(n_239),
.B(n_244),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_153),
.Y(n_242)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_242),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_54),
.B1(n_57),
.B2(n_23),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_243),
.A2(n_273),
.B1(n_289),
.B2(n_295),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_139),
.B(n_4),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_149),
.A2(n_57),
.B(n_23),
.C(n_6),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_246),
.A2(n_244),
.B(n_268),
.C(n_239),
.Y(n_353)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_134),
.Y(n_247)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_251),
.Y(n_354)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_253),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_184),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_254),
.B(n_272),
.Y(n_369)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

BUFx4f_ASAP7_75t_SL g358 ( 
.A(n_258),
.Y(n_358)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_154),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_260),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_145),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_264),
.B(n_267),
.Y(n_342)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_225),
.Y(n_265)
);

BUFx4f_ASAP7_75t_SL g367 ( 
.A(n_265),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_194),
.A2(n_57),
.B1(n_23),
.B2(n_6),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_266),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_160),
.B(n_4),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_143),
.B(n_4),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_171),
.C(n_207),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_202),
.Y(n_269)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_197),
.B(n_5),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_149),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_180),
.Y(n_274)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_160),
.B(n_166),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_278),
.Y(n_313)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_155),
.Y(n_277)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_151),
.B(n_156),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_282),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_140),
.B(n_167),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_198),
.Y(n_286)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_168),
.Y(n_288)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_140),
.A2(n_23),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_221),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_312),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_135),
.A2(n_162),
.B1(n_199),
.B2(n_209),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_292),
.A2(n_298),
.B1(n_304),
.B2(n_305),
.Y(n_322)
);

NAND2xp67_ASAP7_75t_SL g293 ( 
.A(n_136),
.B(n_5),
.Y(n_293)
);

OR2x4_ASAP7_75t_L g350 ( 
.A(n_293),
.B(n_301),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_218),
.B(n_8),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_144),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_179),
.Y(n_297)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_174),
.A2(n_219),
.B1(n_185),
.B2(n_203),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_177),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_302),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_300),
.A2(n_306),
.B1(n_285),
.B2(n_296),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_144),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_301),
.A2(n_311),
.B1(n_295),
.B2(n_235),
.Y(n_321)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_141),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_148),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_307),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_159),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_304)
);

AOI22x1_ASAP7_75t_SL g306 ( 
.A1(n_175),
.A2(n_182),
.B1(n_178),
.B2(n_150),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_172),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_157),
.B(n_163),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_308),
.B(n_309),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_158),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_211),
.A2(n_190),
.B1(n_152),
.B2(n_204),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_310),
.A2(n_188),
.B1(n_193),
.B2(n_212),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_182),
.A2(n_181),
.B1(n_207),
.B2(n_165),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_133),
.B(n_201),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_315),
.B(n_331),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_328),
.B1(n_340),
.B2(n_239),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_305),
.A2(n_226),
.B1(n_148),
.B2(n_188),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_324),
.A2(n_345),
.B1(n_349),
.B2(n_269),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_280),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_325),
.B(n_307),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_133),
.B1(n_201),
.B2(n_212),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_229),
.B(n_226),
.C(n_193),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_333),
.A2(n_344),
.B1(n_259),
.B2(n_346),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_233),
.C(n_246),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_337),
.B(n_343),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_305),
.A2(n_243),
.B1(n_311),
.B2(n_312),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_256),
.B(n_290),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_290),
.A2(n_291),
.B1(n_306),
.B2(n_271),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_258),
.A2(n_265),
.B1(n_274),
.B2(n_232),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_247),
.A2(n_252),
.B1(n_287),
.B2(n_281),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_350),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_353),
.B(n_297),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_293),
.A2(n_300),
.B(n_262),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_255),
.B(n_241),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_260),
.B(n_286),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_244),
.B(n_268),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_231),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_374),
.A2(n_381),
.B1(n_390),
.B2(n_394),
.Y(n_459)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_331),
.B(n_336),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_375),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_376),
.B(n_358),
.Y(n_430)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_341),
.A2(n_333),
.B1(n_336),
.B2(n_322),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_313),
.B(n_240),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_387),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_323),
.A2(n_251),
.B(n_282),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_386),
.A2(n_412),
.B(n_414),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_288),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_388),
.A2(n_406),
.B(n_326),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_341),
.A2(n_279),
.B1(n_253),
.B2(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_248),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_392),
.B(n_407),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_340),
.A2(n_250),
.B1(n_248),
.B2(n_270),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_393),
.A2(n_401),
.B1(n_404),
.B2(n_411),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_341),
.A2(n_270),
.B1(n_277),
.B2(n_249),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_361),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_354),
.Y(n_396)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_396),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_398),
.Y(n_456)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_338),
.Y(n_399)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_399),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_337),
.A2(n_236),
.B1(n_283),
.B2(n_249),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_402),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_314),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_328),
.A2(n_321),
.B1(n_318),
.B2(n_350),
.Y(n_404)
);

MAJx3_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_276),
.C(n_302),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_276),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_359),
.A2(n_303),
.B1(n_261),
.B2(n_242),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_409),
.A2(n_413),
.B1(n_418),
.B2(n_406),
.Y(n_443)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_338),
.Y(n_410)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_359),
.A2(n_323),
.B1(n_315),
.B2(n_343),
.Y(n_411)
);

NAND2x1p5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_303),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_362),
.A2(n_330),
.B(n_326),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_335),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_332),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_320),
.B1(n_316),
.B2(n_342),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_416),
.A2(n_417),
.B1(n_419),
.B2(n_367),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_316),
.A2(n_342),
.B1(n_319),
.B2(n_347),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_319),
.A2(n_347),
.B1(n_360),
.B2(n_370),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_339),
.B(n_365),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_380),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_358),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_421),
.B(n_332),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_334),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_426),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_351),
.C(n_365),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_427),
.B(n_437),
.C(n_461),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_400),
.B(n_339),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_428),
.B(n_436),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_409),
.A2(n_334),
.B1(n_317),
.B2(n_325),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_429),
.A2(n_396),
.B1(n_408),
.B2(n_456),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_430),
.B(n_448),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_442),
.B(n_443),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_416),
.B(n_373),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_373),
.C(n_317),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_441),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_439),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_387),
.B(n_329),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_388),
.A2(n_329),
.B(n_356),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_374),
.A2(n_360),
.B1(n_367),
.B2(n_370),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_447),
.A2(n_462),
.B1(n_390),
.B2(n_419),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_348),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_460),
.Y(n_501)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_377),
.B(n_367),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_375),
.B(n_363),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_404),
.A2(n_368),
.B1(n_363),
.B2(n_348),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_459),
.A2(n_393),
.B1(n_406),
.B2(n_418),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_465),
.A2(n_473),
.B1(n_448),
.B2(n_462),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_461),
.B(n_385),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_466),
.B(n_450),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_385),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_472),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_440),
.A2(n_384),
.B(n_411),
.Y(n_470)
);

AOI21x1_ASAP7_75t_SL g518 ( 
.A1(n_470),
.A2(n_464),
.B(n_496),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_425),
.B(n_395),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_471),
.B(n_488),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_389),
.Y(n_472)
);

OAI22x1_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_381),
.B1(n_412),
.B2(n_397),
.Y(n_473)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_389),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_440),
.A2(n_386),
.B(n_412),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_476),
.A2(n_496),
.B(n_442),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_463),
.B(n_376),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_481),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_478),
.A2(n_484),
.B1(n_486),
.B2(n_493),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_460),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_423),
.Y(n_482)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_433),
.A2(n_417),
.B1(n_389),
.B2(n_401),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_424),
.B(n_392),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_430),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_425),
.B(n_405),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_454),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_491),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_490),
.B(n_492),
.Y(n_510)
);

OA22x2_ASAP7_75t_L g491 ( 
.A1(n_459),
.A2(n_422),
.B1(n_394),
.B2(n_379),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_383),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_433),
.A2(n_407),
.B1(n_414),
.B2(n_420),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_454),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_498),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_434),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_499),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_448),
.A2(n_382),
.B(n_403),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_441),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_424),
.B(n_356),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_438),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_447),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_503),
.B(n_481),
.Y(n_557)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_506),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_508),
.A2(n_529),
.B1(n_537),
.B2(n_538),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_471),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_509),
.B(n_524),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_469),
.B(n_446),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g565 ( 
.A(n_511),
.B(n_525),
.C(n_526),
.Y(n_565)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_515),
.B(n_534),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_476),
.A2(n_446),
.B(n_456),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g554 ( 
.A1(n_516),
.A2(n_517),
.B(n_503),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_464),
.A2(n_458),
.B(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_518),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_501),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_520),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_501),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_522),
.Y(n_567)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_480),
.Y(n_523)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_477),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_472),
.B(n_432),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_466),
.B(n_497),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_500),
.A2(n_432),
.B1(n_431),
.B2(n_450),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_533),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_474),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_531),
.B(n_498),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_489),
.B(n_431),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_497),
.B(n_445),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_SL g568 ( 
.A(n_535),
.B(n_511),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_536),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_485),
.A2(n_445),
.B1(n_452),
.B2(n_455),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_491),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_505),
.B(n_475),
.C(n_470),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_540),
.B(n_544),
.C(n_547),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_505),
.B(n_475),
.C(n_467),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_468),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_545),
.B(n_560),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_507),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_546),
.A2(n_563),
.B1(n_506),
.B2(n_491),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_467),
.C(n_487),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_486),
.C(n_473),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_555),
.C(n_564),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_554),
.A2(n_557),
.B(n_518),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_525),
.B(n_473),
.C(n_494),
.Y(n_555)
);

BUFx12_ASAP7_75t_L g556 ( 
.A(n_515),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_556),
.Y(n_595)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_528),
.Y(n_558)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_558),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_527),
.A2(n_483),
.B1(n_485),
.B2(n_478),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_559),
.A2(n_508),
.B1(n_507),
.B2(n_514),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_528),
.B(n_483),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_514),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_566),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_502),
.B(n_465),
.C(n_491),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_455),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_568),
.B(n_534),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_519),
.B(n_449),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_569),
.B(n_452),
.Y(n_594)
);

XNOR2x1_ASAP7_75t_SL g604 ( 
.A(n_572),
.B(n_568),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_557),
.A2(n_550),
.B(n_552),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g610 ( 
.A1(n_573),
.A2(n_554),
.B(n_564),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_513),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_577),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_539),
.Y(n_578)
);

CKINVDCx14_ASAP7_75t_R g613 ( 
.A(n_578),
.Y(n_613)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_579),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_542),
.A2(n_504),
.B1(n_536),
.B2(n_538),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_581),
.A2(n_583),
.B1(n_587),
.B2(n_589),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_582),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_552),
.A2(n_530),
.B1(n_513),
.B2(n_520),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_549),
.Y(n_584)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_585),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_502),
.C(n_517),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_586),
.B(n_550),
.C(n_561),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_567),
.A2(n_516),
.B1(n_522),
.B2(n_533),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_539),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_588),
.B(n_590),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_567),
.A2(n_523),
.B1(n_521),
.B2(n_512),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_543),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_540),
.B(n_491),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_591),
.B(n_551),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_592),
.A2(n_593),
.B1(n_594),
.B2(n_596),
.Y(n_606)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_541),
.Y(n_593)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_541),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_565),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_599),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_580),
.B(n_555),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_586),
.B(n_547),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_601),
.B(n_607),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_602),
.B(n_604),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_591),
.B(n_544),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_609),
.B(n_614),
.Y(n_621)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_610),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_576),
.B(n_554),
.C(n_561),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_612),
.B(n_617),
.C(n_595),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_556),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_556),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_616),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_572),
.B(n_570),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_618),
.B(n_604),
.Y(n_647)
);

INVx11_ASAP7_75t_L g620 ( 
.A(n_613),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_620),
.A2(n_629),
.B1(n_590),
.B2(n_574),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_581),
.C(n_573),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_622),
.B(n_624),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_577),
.C(n_587),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_611),
.A2(n_578),
.B1(n_588),
.B2(n_579),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_625),
.A2(n_608),
.B1(n_628),
.B2(n_619),
.Y(n_636)
);

FAx1_ASAP7_75t_SL g626 ( 
.A(n_612),
.B(n_577),
.CI(n_583),
.CON(n_626),
.SN(n_626)
);

MAJIxp5_ASAP7_75t_R g643 ( 
.A(n_626),
.B(n_600),
.C(n_616),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_584),
.C(n_589),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_627),
.B(n_630),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_615),
.A2(n_598),
.B(n_605),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_571),
.C(n_575),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_606),
.Y(n_631)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_631),
.Y(n_640)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_603),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_630),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_615),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_634),
.B(n_596),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_636),
.B(n_643),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g638 ( 
.A(n_618),
.B(n_627),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_638),
.B(n_644),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_639),
.Y(n_652)
);

MAJx2_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_607),
.C(n_609),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_642),
.B(n_646),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_617),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g645 ( 
.A(n_626),
.Y(n_645)
);

BUFx24_ASAP7_75t_SL g655 ( 
.A(n_645),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_631),
.A2(n_608),
.B1(n_571),
.B2(n_558),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_647),
.B(n_649),
.Y(n_658)
);

OAI321xp33_ASAP7_75t_L g657 ( 
.A1(n_648),
.A2(n_640),
.A3(n_620),
.B1(n_548),
.B2(n_570),
.C(n_553),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_622),
.B(n_593),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_619),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_621),
.C(n_623),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_654),
.B(n_656),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_623),
.C(n_621),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_657),
.B(n_659),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_643),
.B(n_624),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_661),
.B(n_642),
.Y(n_668)
);

AND2x4_ASAP7_75t_SL g662 ( 
.A(n_655),
.B(n_641),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_662),
.Y(n_672)
);

XOR2x2_ASAP7_75t_L g663 ( 
.A(n_653),
.B(n_644),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_663),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_656),
.B(n_658),
.C(n_660),
.Y(n_665)
);

A2O1A1O1Ixp25_ASAP7_75t_L g671 ( 
.A1(n_665),
.A2(n_635),
.B(n_660),
.C(n_633),
.D(n_553),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_651),
.A2(n_652),
.B(n_625),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g669 ( 
.A1(n_666),
.A2(n_668),
.B(n_626),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_SL g674 ( 
.A1(n_669),
.A2(n_671),
.B(n_667),
.Y(n_674)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_670),
.B(n_664),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_SL g675 ( 
.A1(n_673),
.A2(n_674),
.B(n_666),
.Y(n_675)
);

AOI322xp5_ASAP7_75t_L g676 ( 
.A1(n_675),
.A2(n_672),
.A3(n_548),
.B1(n_633),
.B2(n_444),
.C1(n_449),
.C2(n_421),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_444),
.C(n_451),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_677),
.B(n_422),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_451),
.B(n_402),
.Y(n_679)
);

MAJx2_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_399),
.C(n_410),
.Y(n_680)
);


endmodule