module fake_jpeg_20354_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_12),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_19),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_51),
.B1(n_62),
.B2(n_30),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_28),
.B1(n_25),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_50),
.B1(n_59),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_35),
.B1(n_22),
.B2(n_32),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_34),
.B(n_18),
.C(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_R g86 ( 
.A(n_53),
.B(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_20),
.B1(n_34),
.B2(n_18),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_19),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_52),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_35),
.B1(n_23),
.B2(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_43),
.B1(n_23),
.B2(n_35),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_97),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_69),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_71),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_78),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_43),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_80),
.C(n_89),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_38),
.B1(n_36),
.B2(n_41),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_76),
.B1(n_94),
.B2(n_100),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_36),
.B(n_18),
.C(n_34),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_31),
.B1(n_32),
.B2(n_22),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_82),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_31),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_88),
.Y(n_126)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_26),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_30),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_24),
.B1(n_39),
.B2(n_41),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_24),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_102),
.B1(n_39),
.B2(n_17),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_24),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_62),
.B(n_36),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_127),
.B(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_75),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_39),
.B1(n_26),
.B2(n_17),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_121),
.B1(n_128),
.B2(n_6),
.Y(n_147)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_93),
.C(n_83),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_104),
.Y(n_180)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_72),
.B(n_86),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_137),
.B(n_138),
.Y(n_182)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_66),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_96),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_99),
.B1(n_92),
.B2(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_80),
.B1(n_66),
.B2(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_70),
.B1(n_68),
.B2(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_85),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_6),
.C(n_7),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_7),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_117),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_121),
.B1(n_115),
.B2(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_147),
.B1(n_132),
.B2(n_158),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_188),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_174),
.B(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_133),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_178),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_126),
.B(n_107),
.C(n_115),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_104),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_185),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_107),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_150),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_204),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_139),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_201),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_103),
.B(n_145),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_209),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_132),
.B1(n_127),
.B2(n_152),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_213),
.C(n_215),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_127),
.B(n_155),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_165),
.A2(n_108),
.B1(n_128),
.B2(n_116),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_157),
.B1(n_110),
.B2(n_111),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_172),
.A2(n_118),
.A3(n_111),
.B1(n_157),
.B2(n_113),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_197),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_118),
.C(n_85),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_113),
.C(n_67),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_179),
.C(n_166),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_229),
.C(n_231),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_176),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_178),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_196),
.B(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_163),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_188),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_227),
.A2(n_230),
.B1(n_195),
.B2(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_170),
.C(n_166),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_170),
.C(n_183),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_235),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_189),
.B1(n_162),
.B2(n_183),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_210),
.B1(n_209),
.B2(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_234),
.A2(n_192),
.B1(n_197),
.B2(n_233),
.Y(n_238)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_231),
.C(n_221),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_243),
.C(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_201),
.C(n_215),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_220),
.B(n_229),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_249),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_168),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_253),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_217),
.A2(n_168),
.B(n_190),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_224),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_181),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_163),
.C(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_174),
.C(n_169),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_164),
.C(n_10),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_164),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_252),
.B1(n_164),
.B2(n_12),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_216),
.B1(n_227),
.B2(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_249),
.B1(n_247),
.B2(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_251),
.B(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_253),
.C(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_244),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_266),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_258),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_271),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_259),
.A2(n_236),
.B1(n_237),
.B2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_273),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_16),
.B1(n_11),
.B2(n_13),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_276),
.B(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_258),
.C(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_279),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_284),
.C(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_274),
.Y(n_284)
);

A2O1A1O1Ixp25_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_271),
.B(n_272),
.C(n_267),
.D(n_261),
.Y(n_285)
);

OAI211xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_275),
.B(n_283),
.C(n_13),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_278),
.B(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_9),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_286),
.C(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_294),
.B(n_9),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.Y(n_296)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_9),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.C(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_14),
.Y(n_298)
);


endmodule