module fake_jpeg_27073_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_0),
.C(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

OAI221xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_20),
.B1(n_21),
.B2(n_9),
.C(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_19),
.B(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_2),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_24),
.B1(n_14),
.B2(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_11),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_11),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_17),
.B1(n_8),
.B2(n_21),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.Y(n_31)
);

OA21x2_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_12),
.B(n_4),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_16),
.B1(n_12),
.B2(n_7),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_27),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_22),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_37),
.B(n_26),
.Y(n_40)
);


endmodule