module real_jpeg_19668_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_52),
.B1(n_57),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_60),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_0),
.A2(n_36),
.B1(n_37),
.B2(n_60),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_68),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_1),
.A2(n_15),
.B(n_27),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_64),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_104),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_1),
.A2(n_57),
.B(n_165),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_2),
.A2(n_48),
.B1(n_52),
.B2(n_57),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_48),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_63),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_52),
.B1(n_57),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_71),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_5),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_5),
.A2(n_58),
.B1(n_63),
.B2(n_72),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_27),
.B1(n_29),
.B2(n_58),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_41),
.Y(n_108)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g159 ( 
.A1(n_13),
.A2(n_37),
.A3(n_57),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_15),
.A2(n_27),
.B1(n_29),
.B2(n_38),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_21),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_25),
.A2(n_28),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_25),
.A2(n_26),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_25),
.A2(n_89),
.B1(n_120),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_25),
.A2(n_26),
.B1(n_122),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_25),
.A2(n_26),
.B1(n_108),
.B2(n_152),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_26),
.B(n_64),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_29),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_34),
.A2(n_39),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_34),
.A2(n_39),
.B1(n_130),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_34),
.A2(n_39),
.B1(n_150),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_34),
.A2(n_39),
.B1(n_47),
.B2(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_36),
.B(n_53),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_37),
.A2(n_38),
.B(n_64),
.C(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_39),
.B(n_64),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_61),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_55),
.B1(n_59),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_51),
.A2(n_55),
.B1(n_101),
.B2(n_164),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_57),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_62),
.B1(n_67),
.B2(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_52),
.B(n_64),
.Y(n_161)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_66),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.CON(n_62),
.SN(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_84),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_81),
.B2(n_83),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_117)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_97),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_93),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.C(n_106),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_99),
.B(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_105),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_187),
.B(n_191),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_173),
.B(n_186),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_154),
.B(n_172),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_142),
.B(n_153),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_131),
.B(n_141),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_123),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_136),
.B(n_140),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_135),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_144),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_151),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_162),
.B1(n_170),
.B2(n_171),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_159),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_169),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_175),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_183),
.C(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_182),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);


endmodule