module fake_jpeg_4430_n_336 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_17),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_63),
.Y(n_113)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_65),
.B(n_70),
.Y(n_132)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_73),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_15),
.B1(n_29),
.B2(n_14),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_116)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_38),
.A2(n_15),
.B1(n_29),
.B2(n_14),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_25),
.Y(n_76)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_37),
.A2(n_17),
.B1(n_23),
.B2(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_37),
.A2(n_43),
.B1(n_45),
.B2(n_23),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_35),
.B1(n_30),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_84),
.B(n_87),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_54),
.B1(n_57),
.B2(n_53),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_6),
.B(n_104),
.C(n_84),
.Y(n_133)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_39),
.A2(n_22),
.B1(n_19),
.B2(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_46),
.A2(n_28),
.B1(n_22),
.B2(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_102),
.B1(n_33),
.B2(n_3),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_46),
.A2(n_22),
.B1(n_32),
.B2(n_34),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_33),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_26),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_28),
.B1(n_22),
.B2(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_33),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_127),
.B1(n_67),
.B2(n_95),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_125),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_130),
.B1(n_93),
.B2(n_68),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_13),
.B(n_10),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_134),
.B(n_62),
.C(n_61),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_128),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_10),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_9),
.B1(n_8),
.B2(n_4),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_90),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_2),
.C(n_6),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_83),
.B(n_63),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_101),
.B(n_105),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_71),
.A2(n_92),
.B1(n_97),
.B2(n_86),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_59),
.B(n_74),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_74),
.C(n_60),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_72),
.C(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_64),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_88),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_72),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_140),
.A2(n_149),
.B(n_173),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_176),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_87),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_147),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_150),
.B(n_156),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_58),
.Y(n_164)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

BUFx2_ASAP7_75t_SL g165 ( 
.A(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_124),
.B(n_58),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_171),
.Y(n_194)
);

INVx6_ASAP7_75t_SL g172 ( 
.A(n_107),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_158),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_108),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_134),
.B1(n_130),
.B2(n_112),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_122),
.B1(n_117),
.B2(n_120),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_122),
.A2(n_117),
.B1(n_113),
.B2(n_129),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_120),
.B1(n_171),
.B2(n_167),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_202),
.B1(n_203),
.B2(n_208),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_121),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_187),
.C(n_201),
.Y(n_232)
);

HAxp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_121),
.CON(n_184),
.SN(n_184)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_189),
.B(n_193),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_121),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_195),
.B1(n_161),
.B2(n_189),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_120),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_149),
.B(n_155),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_141),
.B1(n_143),
.B2(n_173),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_210),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_140),
.C(n_145),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_156),
.B1(n_159),
.B2(n_172),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_147),
.A2(n_153),
.B(n_166),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_152),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_146),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_142),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_146),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_161),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_210),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_219),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_146),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_204),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_177),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_230),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_196),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_243),
.C(n_185),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_198),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_188),
.A2(n_202),
.B1(n_214),
.B2(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_241),
.B(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_182),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_202),
.C(n_205),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_184),
.B(n_203),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_216),
.B(n_228),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_259),
.C(n_264),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_205),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_185),
.B(n_207),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_225),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_235),
.B1(n_241),
.B2(n_224),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_198),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_211),
.C(n_197),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_266),
.C(n_267),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_190),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_231),
.B(n_211),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_236),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_283),
.C(n_285),
.Y(n_295)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_237),
.B1(n_190),
.B2(n_263),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_273),
.B1(n_247),
.B2(n_260),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_226),
.B1(n_239),
.B2(n_243),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_279),
.B1(n_221),
.B2(n_197),
.Y(n_294)
);

OA21x2_ASAP7_75t_SL g276 ( 
.A1(n_266),
.A2(n_215),
.B(n_220),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_259),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_219),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_222),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_258),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_240),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_213),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_230),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_217),
.C(n_233),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_285),
.B(n_247),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_252),
.B1(n_244),
.B2(n_255),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_289),
.B1(n_299),
.B2(n_246),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_244),
.B1(n_255),
.B2(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_281),
.B(n_217),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_265),
.C(n_267),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_275),
.C(n_277),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_277),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_306),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_278),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_295),
.C(n_282),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_287),
.B(n_299),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_303),
.Y(n_319)
);

OA21x2_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_291),
.B(n_292),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_306),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_296),
.B1(n_289),
.B2(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_296),
.B1(n_288),
.B2(n_295),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_304),
.B1(n_249),
.B2(n_268),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_282),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.C(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_293),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_221),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_313),
.C(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_329),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_323),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_318),
.C(n_302),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_318),
.C(n_320),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_321),
.B1(n_331),
.B2(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_328),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_314),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_257),
.Y(n_336)
);


endmodule