module fake_jpeg_21041_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_46),
.B(n_47),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_49),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_50),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_29),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_57),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_23),
.B(n_1),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_69),
.Y(n_89)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_70),
.Y(n_130)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_2),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_28),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_77),
.Y(n_131)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_2),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_33),
.B(n_20),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_16),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_42),
.B1(n_39),
.B2(n_34),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_32),
.B1(n_40),
.B2(n_38),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_91),
.A2(n_101),
.B1(n_110),
.B2(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_84),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_26),
.B1(n_40),
.B2(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_96),
.A2(n_105),
.B1(n_108),
.B2(n_113),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_31),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g175 ( 
.A1(n_100),
.A2(n_12),
.B(n_124),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_18),
.B1(n_37),
.B2(n_36),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_69),
.A2(n_61),
.B1(n_74),
.B2(n_51),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_103),
.A2(n_50),
.B1(n_82),
.B2(n_12),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_18),
.B1(n_37),
.B2(n_36),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_57),
.A2(n_16),
.B1(n_26),
.B2(n_42),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_67),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_113)
);

OR2x4_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_45),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_71),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_122),
.A2(n_135),
.B1(n_129),
.B2(n_88),
.Y(n_181)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_127)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_49),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_44),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_83),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_147),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_55),
.B1(n_81),
.B2(n_63),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_142),
.B(n_164),
.Y(n_215)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_144),
.B(n_150),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_178),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_8),
.C(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_68),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_89),
.B(n_82),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_54),
.B1(n_64),
.B2(n_48),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_166),
.B1(n_125),
.B2(n_128),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_58),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_76),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_76),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_168),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_76),
.C(n_82),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g167 ( 
.A(n_112),
.Y(n_167)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_8),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_172),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_10),
.B(n_12),
.C(n_99),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_117),
.B(n_128),
.C(n_106),
.Y(n_207)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_99),
.B(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_177),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_116),
.B(n_98),
.Y(n_188)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_181),
.B1(n_129),
.B2(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_92),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_102),
.B(n_92),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_116),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_104),
.B(n_138),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_148),
.B1(n_166),
.B2(n_181),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_207),
.C(n_149),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_88),
.B1(n_114),
.B2(n_119),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_142),
.A2(n_159),
.B1(n_158),
.B2(n_140),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_114),
.B1(n_119),
.B2(n_97),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_104),
.B1(n_134),
.B2(n_106),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_195),
.A2(n_212),
.B1(n_208),
.B2(n_215),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_214),
.B1(n_173),
.B2(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_136),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_218),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_158),
.A2(n_117),
.B(n_90),
.C(n_111),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_210),
.B(n_149),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_144),
.A2(n_90),
.B(n_111),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_182),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_146),
.B1(n_172),
.B2(n_143),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_176),
.B1(n_165),
.B2(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_152),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_145),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_223),
.A2(n_233),
.B(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_225),
.B(n_231),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_254),
.B1(n_211),
.B2(n_203),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_228),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_153),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_229),
.B(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_235),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_153),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_170),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_237),
.A2(n_239),
.B(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_238),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_188),
.B(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_194),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_201),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_202),
.Y(n_273)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_204),
.B(n_206),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_189),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_207),
.B(n_186),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_250),
.B(n_187),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_215),
.A2(n_207),
.B1(n_190),
.B2(n_191),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_197),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_252),
.A2(n_206),
.B1(n_210),
.B2(n_189),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_199),
.A2(n_208),
.B1(n_192),
.B2(n_195),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_252),
.B1(n_248),
.B2(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_263),
.A2(n_265),
.B1(n_276),
.B2(n_277),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_220),
.C(n_213),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_234),
.C(n_240),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_230),
.A2(n_220),
.B1(n_213),
.B2(n_217),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_222),
.B1(n_245),
.B2(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_273),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_234),
.A2(n_187),
.B1(n_202),
.B2(n_184),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_237),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_247),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_274),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_279),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_203),
.B1(n_196),
.B2(n_217),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_200),
.B1(n_196),
.B2(n_184),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_200),
.B1(n_184),
.B2(n_198),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_232),
.Y(n_283)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_259),
.B(n_246),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_291),
.Y(n_321)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_295),
.Y(n_309)
);

OR2x2_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_233),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_275),
.B(n_272),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_288),
.B(n_281),
.C(n_278),
.Y(n_323)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_290),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_228),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_229),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_280),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_298),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_231),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_278),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_257),
.B(n_227),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_266),
.B(n_234),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_281),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_255),
.B1(n_267),
.B2(n_273),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_264),
.B(n_223),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_270),
.B1(n_282),
.B2(n_255),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_308),
.B(n_324),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_310),
.A2(n_287),
.B(n_283),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_263),
.B1(n_268),
.B2(n_269),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_316),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_327),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_258),
.B1(n_270),
.B2(n_223),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_289),
.A2(n_299),
.B1(n_226),
.B2(n_290),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_320),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_265),
.B1(n_279),
.B2(n_276),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_304),
.C(n_302),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_277),
.B1(n_261),
.B2(n_262),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_261),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_306),
.Y(n_346)
);

BUFx12_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_335),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_285),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_333),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_322),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_341),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_325),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_338),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

INVx11_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_328),
.B(n_297),
.C(n_295),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_308),
.C(n_313),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_298),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_287),
.B(n_293),
.C(n_297),
.D(n_296),
.Y(n_345)
);

AOI321xp33_ASAP7_75t_L g360 ( 
.A1(n_345),
.A2(n_294),
.A3(n_307),
.B1(n_291),
.B2(n_300),
.C(n_262),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_340),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_329),
.A2(n_311),
.B1(n_320),
.B2(n_319),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_352),
.B1(n_356),
.B2(n_332),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g351 ( 
.A1(n_342),
.A2(n_326),
.B(n_321),
.Y(n_351)
);

FAx1_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_360),
.CI(n_345),
.CON(n_363),
.SN(n_363)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_344),
.A2(n_312),
.B1(n_316),
.B2(n_305),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_330),
.A2(n_318),
.B(n_303),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_353),
.A2(n_336),
.B(n_330),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_344),
.A2(n_323),
.B1(n_327),
.B2(n_317),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_343),
.C(n_346),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_359),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_338),
.A2(n_324),
.B1(n_307),
.B2(n_286),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_354),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_366),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_364),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_365),
.B(n_367),
.Y(n_379)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_370),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g369 ( 
.A1(n_360),
.A2(n_332),
.B(n_235),
.C(n_242),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_349),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_337),
.C(n_286),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_356),
.C(n_358),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_376),
.C(n_377),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_369),
.A2(n_363),
.B1(n_347),
.B2(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_371),
.A2(n_359),
.B(n_355),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_355),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_378),
.A2(n_369),
.B1(n_363),
.B2(n_361),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_385),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g383 ( 
.A(n_379),
.B(n_367),
.C(n_369),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_238),
.C(n_241),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_372),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_374),
.B(n_380),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_387),
.Y(n_392)
);

AOI322xp5_ASAP7_75t_L g388 ( 
.A1(n_386),
.A2(n_362),
.A3(n_352),
.B1(n_377),
.B2(n_224),
.C1(n_337),
.C2(n_292),
.Y(n_388)
);

AOI322xp5_ASAP7_75t_L g393 ( 
.A1(n_388),
.A2(n_390),
.A3(n_244),
.B1(n_251),
.B2(n_292),
.C1(n_249),
.C2(n_200),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_384),
.C(n_385),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_393),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_251),
.C(n_249),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_395),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_394),
.Y(n_397)
);


endmodule