module real_jpeg_6410_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_0),
.A2(n_148),
.B1(n_151),
.B2(n_154),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_0),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_0),
.B(n_171),
.C(n_174),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_0),
.B(n_74),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_0),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_0),
.B(n_165),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_0),
.B(n_264),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_1),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_1),
.Y(n_237)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_1),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_1),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_2),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_2),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_53),
.B1(n_88),
.B2(n_128),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_2),
.A2(n_88),
.B1(n_384),
.B2(n_386),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_2),
.A2(n_88),
.B1(n_249),
.B2(n_417),
.Y(n_416)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_3),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_3),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_3),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_3),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_4),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_5),
.A2(n_118),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_5),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_5),
.A2(n_179),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_5),
.A2(n_179),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_5),
.A2(n_56),
.B1(n_179),
.B2(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_6),
.Y(n_333)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_7),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_8),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_8),
.A2(n_57),
.B1(n_224),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_8),
.A2(n_57),
.B1(n_164),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_8),
.A2(n_57),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_9),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_11),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_12),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_12),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_160),
.B1(n_192),
.B2(n_196),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_12),
.A2(n_160),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_12),
.A2(n_160),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_14),
.A2(n_157),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_206),
.B1(n_221),
.B2(n_225),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_14),
.A2(n_41),
.B1(n_206),
.B2(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_14),
.A2(n_32),
.B1(n_48),
.B2(n_206),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_15),
.A2(n_49),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_15),
.A2(n_49),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_15),
.A2(n_49),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_16),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_16),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_94),
.B1(n_100),
.B2(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_16),
.A2(n_32),
.B1(n_94),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_16),
.A2(n_94),
.B1(n_180),
.B2(n_388),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_17),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_17),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_17),
.A2(n_277),
.B1(n_371),
.B2(n_373),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_17),
.A2(n_277),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_17),
.A2(n_277),
.B1(n_330),
.B2(n_457),
.Y(n_456)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_531),
.B(n_534),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_137),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_135),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_132),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_132),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_126),
.C(n_129),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_24),
.A2(n_25),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_58),
.C(n_95),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_26),
.B(n_519),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_27),
.A2(n_50),
.B1(n_52),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_50),
.B1(n_127),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_27),
.A2(n_357),
.B(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_27),
.A2(n_50),
.B1(n_411),
.B2(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_27),
.A2(n_46),
.B1(n_50),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_28),
.A2(n_337),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_28),
.B(n_358),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_32),
.Y(n_359)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_41),
.B2(n_44),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_39),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_40),
.Y(n_409)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_45),
.Y(n_335)
);

INVx6_ASAP7_75t_L g412 ( 
.A(n_47),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_50),
.B(n_154),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_50),
.A2(n_431),
.B(n_458),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_51),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_51),
.B(n_456),
.Y(n_455)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_58),
.A2(n_95),
.B1(n_96),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_58),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_84),
.B1(n_89),
.B2(n_90),
.Y(n_58)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_59),
.A2(n_89),
.B1(n_301),
.B2(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_59),
.A2(n_89),
.B1(n_400),
.B2(n_405),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_59),
.A2(n_84),
.B1(n_89),
.B2(n_508),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_74),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_65),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_68),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_68),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_68),
.Y(n_329)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_68),
.Y(n_336)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_73),
.Y(n_303)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_73),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_74),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_74),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_74),
.A2(n_130),
.B1(n_305),
.B2(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_74),
.A2(n_130),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g372 ( 
.A(n_77),
.Y(n_372)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_77),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_78),
.Y(n_254)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_79),
.Y(n_397)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_82),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_86),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_87),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_89),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_89),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_95),
.A2(n_96),
.B1(n_506),
.B2(n_507),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_95),
.B(n_503),
.C(n_506),
.Y(n_514)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_110),
.B(n_121),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_97),
.A2(n_147),
.B(n_155),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_97),
.A2(n_110),
.B1(n_204),
.B2(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_97),
.A2(n_155),
.B(n_248),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_97),
.A2(n_110),
.B1(n_370),
.B2(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_98),
.B(n_156),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_98),
.A2(n_165),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_98),
.A2(n_165),
.B1(n_394),
.B2(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_98),
.A2(n_165),
.B1(n_416),
.B2(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_102),
.Y(n_251)
);

INVx6_ASAP7_75t_L g374 ( 
.A(n_102),
.Y(n_374)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_110),
.A2(n_204),
.B(n_207),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_110),
.A2(n_207),
.B(n_370),
.Y(n_369)
);

AOI22x1_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_118),
.B2(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_116),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_118),
.B(n_214),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_119),
.Y(n_314)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_119),
.Y(n_385)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_121),
.Y(n_447)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_125),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_126),
.B(n_129),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_130),
.A2(n_257),
.B(n_265),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_130),
.B(n_305),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_130),
.A2(n_265),
.B(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_525),
.B(n_530),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_497),
.B(n_522),
.Y(n_138)
);

OAI311xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_377),
.A3(n_473),
.B1(n_491),
.C1(n_496),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_320),
.B(n_376),
.Y(n_140)
);

AO21x2_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_292),
.B(n_319),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_242),
.B(n_291),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_210),
.B(n_241),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_176),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_166),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_146),
.A2(n_166),
.B1(n_167),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_154),
.A2(n_185),
.B(n_188),
.Y(n_217)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_154),
.A2(n_258),
.B(n_262),
.Y(n_257)
);

HAxp5_ASAP7_75t_SL g337 ( 
.A(n_154),
.B(n_338),
.CON(n_337),
.SN(n_337)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_SL g418 ( 
.A(n_169),
.Y(n_418)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_201),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_202),
.C(n_209),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_185),
.B(n_188),
.Y(n_177)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_185),
.A2(n_343),
.B1(n_344),
.B2(n_347),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_185),
.A2(n_280),
.B1(n_383),
.B2(n_387),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_185),
.A2(n_228),
.B(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_191),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_186),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_186),
.A2(n_275),
.B1(n_309),
.B2(n_315),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_186),
.A2(n_348),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_197),
.Y(n_310)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_199),
.Y(n_389)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_208),
.B2(n_209),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_232),
.B(n_240),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_218),
.B(n_231),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_230),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_230),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_228),
.B(n_229),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_274),
.B(n_280),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_238),
.Y(n_240)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_244),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_272),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_255),
.C(n_272),
.Y(n_293)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_251),
.Y(n_393)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_261),
.Y(n_406)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_261),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_283),
.A3(n_284),
.B1(n_287),
.B2(n_289),
.Y(n_282)
);

INVx8_ASAP7_75t_L g404 ( 
.A(n_264),
.Y(n_404)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_282),
.Y(n_298)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_279),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_293),
.B(n_294),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_318),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_298),
.C(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_306),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_307),
.C(n_308),
.Y(n_350)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_321),
.B(n_322),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_353),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_323)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_341),
.B2(n_342),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_326),
.B(n_341),
.Y(n_469)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_330),
.A3(n_332),
.B1(n_334),
.B2(n_337),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_350),
.B(n_352),
.C(n_353),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_362),
.B2(n_375),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_354),
.B(n_363),
.C(n_369),
.Y(n_482)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_360),
.Y(n_457)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_369),
.Y(n_362)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx8_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_459),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_SL g491 ( 
.A1(n_378),
.A2(n_459),
.B(n_492),
.C(n_495),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_434),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_379),
.B(n_434),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_413),
.C(n_421),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g472 ( 
.A(n_380),
.B(n_413),
.CI(n_421),
.CON(n_472),
.SN(n_472)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_398),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_381),
.B(n_399),
.C(n_410),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_390),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_382),
.B(n_390),
.Y(n_465)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_410),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_419),
.B2(n_420),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_419),
.Y(n_451)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_419),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_420),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_419),
.A2(n_451),
.B(n_454),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_429),
.C(n_432),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_423),
.B(n_425),
.Y(n_481)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_432),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_438),
.C(n_449),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_449),
.B2(n_450),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_445),
.B(n_448),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_446),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_442),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g499 ( 
.A(n_448),
.B(n_500),
.CI(n_501),
.CON(n_499),
.SN(n_499)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_448),
.B(n_500),
.C(n_501),
.Y(n_521)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_460),
.B(n_472),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_466),
.B(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.C(n_470),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_467),
.A2(n_468),
.B1(n_470),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_472),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_486),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_475),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_483),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_483),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.C(n_482),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_489),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_481),
.B1(n_482),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_488),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_511),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_510),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_499),
.B(n_510),
.Y(n_523)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_499),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_505),
.B2(n_509),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_502),
.A2(n_503),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_513),
.C(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_505),
.Y(n_509)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_523),
.B(n_524),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_521),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_512),
.B(n_521),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_529),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx4f_ASAP7_75t_SL g531 ( 
.A(n_532),
.Y(n_531)
);

INVx13_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx5_ASAP7_75t_L g536 ( 
.A(n_533),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);


endmodule