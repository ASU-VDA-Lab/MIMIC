module fake_jpeg_13057_n_74 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;
wire n_70;
wire n_66;

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_40),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_1),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_47),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_32),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_37),
.B1(n_31),
.B2(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_33),
.C(n_26),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_57),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_54),
.B1(n_59),
.B2(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_26),
.B1(n_3),
.B2(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_3),
.B(n_4),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_13),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_9),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_64),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_65),
.C(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_68),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.C(n_62),
.Y(n_70)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_63),
.B(n_66),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_66),
.B(n_19),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_18),
.Y(n_74)
);


endmodule