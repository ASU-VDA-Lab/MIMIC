module fake_netlist_5_1761_n_1751 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1751);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1751;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_14),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_69),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_126),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_63),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_30),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_64),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_55),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_22),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_58),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_59),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_118),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_34),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_23),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_110),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_89),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_56),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_98),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_54),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_44),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_146),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_12),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_23),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_62),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_151),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_6),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_102),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_74),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_32),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_161),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_96),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_86),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_28),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_38),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_50),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_145),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_12),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_28),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_16),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_54),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_43),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_152),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_143),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_1),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_81),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_45),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_137),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_112),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_123),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_1),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_18),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_117),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_77),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_133),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_160),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_13),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_106),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_79),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_108),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_144),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_157),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_124),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_84),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_16),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_158),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_87),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_66),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_49),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_128),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_7),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_51),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_90),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_24),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_50),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_107),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_41),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_91),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_61),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_17),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_42),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_147),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_40),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_2),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_76),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_125),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_30),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_136),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_65),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_10),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_71),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_9),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_105),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_19),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_58),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_20),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_47),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_88),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_29),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_24),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_35),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_57),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_94),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_29),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_78),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_67),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_4),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_103),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_14),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_35),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_113),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_48),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_26),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_20),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_36),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_41),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_249),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_213),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_187),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_175),
.B(n_266),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_217),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_188),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_221),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_223),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_225),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_316),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_226),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_227),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_232),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_236),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_240),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_199),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_197),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_250),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_299),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_197),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_307),
.B(n_0),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_172),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_208),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_189),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_176),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_177),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_236),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_274),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_211),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_257),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_210),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_177),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_236),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_236),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_216),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_218),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_229),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_264),
.B(n_2),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_258),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_234),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_267),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_236),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_237),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_261),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_177),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_264),
.B(n_3),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_268),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_238),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_262),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_254),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_271),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_272),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_276),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_260),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_269),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_167),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_185),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_185),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_167),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_277),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_282),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_212),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_185),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_170),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_275),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_279),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_252),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_287),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_169),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_252),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_181),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_169),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_373),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_373),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_339),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_343),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_374),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

NAND2xp33_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_181),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_345),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_341),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_382),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_380),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_418),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_346),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_342),
.B(n_171),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_369),
.B(n_293),
.Y(n_452)
);

CKINVDCx6p67_ASAP7_75t_R g453 ( 
.A(n_369),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_347),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_386),
.B(n_170),
.Y(n_456)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_350),
.B(n_264),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_400),
.B(n_173),
.Y(n_459)
);

AND3x1_ASAP7_75t_L g460 ( 
.A(n_394),
.B(n_308),
.C(n_306),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_355),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_350),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_336),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_336),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_349),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_337),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_344),
.A2(n_334),
.B1(n_219),
.B2(n_331),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_352),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_173),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_353),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_356),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_357),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_337),
.B(n_179),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_361),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_419),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_340),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_371),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_340),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_348),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_348),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_351),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_377),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_351),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_380),
.B(n_393),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_387),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_364),
.B(n_288),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_354),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_392),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_397),
.B(n_179),
.Y(n_493)
);

NAND2x1_ASAP7_75t_L g494 ( 
.A(n_354),
.B(n_270),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_358),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_407),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_358),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_399),
.Y(n_498)
);

INVx4_ASAP7_75t_SL g499 ( 
.A(n_457),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_435),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_459),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_465),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_450),
.A2(n_222),
.B1(n_174),
.B2(n_297),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_445),
.B(n_401),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_464),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_445),
.B(n_409),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_470),
.B(n_412),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_435),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_465),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_432),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_436),
.B(n_288),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_436),
.B(n_184),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_490),
.B(n_398),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_467),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_398),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_457),
.B(n_270),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_410),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_464),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_456),
.A2(n_222),
.B1(n_183),
.B2(n_297),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_470),
.B(n_448),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_375),
.Y(n_524)
);

BUFx8_ASAP7_75t_SL g525 ( 
.A(n_437),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_463),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_483),
.B(n_174),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_475),
.B(n_273),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_464),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_432),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_484),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_479),
.B(n_393),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_463),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_485),
.A2(n_183),
.B1(n_324),
.B2(n_312),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_479),
.B(n_416),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_460),
.B(n_270),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_485),
.B(n_416),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_495),
.B(n_270),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_495),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_419),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_422),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_497),
.B(n_168),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_474),
.B(n_338),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_457),
.A2(n_317),
.B1(n_415),
.B2(n_414),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_448),
.B(n_384),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_461),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_452),
.A2(n_333),
.B1(n_304),
.B2(n_309),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_460),
.A2(n_433),
.B1(n_452),
.B2(n_424),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_497),
.B(n_270),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_461),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_480),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_464),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_429),
.B(n_404),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_422),
.B(n_384),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_451),
.B(n_367),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_480),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_494),
.Y(n_563)
);

INVx4_ASAP7_75t_SL g564 ( 
.A(n_457),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_429),
.B(n_364),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_482),
.B(n_178),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_496),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_482),
.B(n_180),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_496),
.B(n_366),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_482),
.B(n_190),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_457),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_457),
.A2(n_417),
.B1(n_415),
.B2(n_414),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_487),
.B(n_200),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_491),
.B(n_201),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_472),
.B(n_366),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_457),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_451),
.B(n_417),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_493),
.B(n_202),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_491),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_476),
.B(n_220),
.C(n_214),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_476),
.B(n_367),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_494),
.A2(n_403),
.B1(n_402),
.B2(n_396),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_454),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_447),
.B(n_370),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_455),
.B(n_370),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_427),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_466),
.B(n_403),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_440),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_454),
.A2(n_402),
.B1(n_396),
.B2(n_391),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_372),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_427),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_453),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_462),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_488),
.B(n_233),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

INVx4_ASAP7_75t_SL g602 ( 
.A(n_427),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_469),
.B(n_209),
.Y(n_603)
);

OR2x2_ASAP7_75t_SL g604 ( 
.A(n_423),
.B(n_231),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_427),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_458),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_441),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_423),
.B(n_372),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_376),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_SL g610 ( 
.A1(n_468),
.A2(n_242),
.B1(n_292),
.B2(n_251),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_458),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_425),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_453),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_425),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_428),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_441),
.B(n_235),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_428),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_430),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_453),
.B(n_311),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_444),
.B(n_376),
.Y(n_620)
);

NOR2x1p5_ASAP7_75t_L g621 ( 
.A(n_473),
.B(n_193),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_441),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_441),
.B(n_243),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_444),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_441),
.B(n_245),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_477),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_440),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_441),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_481),
.B(n_379),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_443),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_430),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_431),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_486),
.B(n_489),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_478),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_478),
.B(n_379),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_431),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_443),
.B(n_256),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_492),
.B(n_383),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_443),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_449),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_498),
.B(n_263),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_449),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_525),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_590),
.B(n_182),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_529),
.A2(n_305),
.B(n_325),
.C(n_319),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_552),
.A2(n_359),
.B1(n_378),
.B2(n_368),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_620),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_524),
.B(n_182),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_591),
.B(n_389),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_520),
.B(n_278),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_590),
.B(n_186),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_584),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_L g655 ( 
.A(n_527),
.B(n_186),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_533),
.B(n_294),
.Y(n_656)
);

CKINVDCx14_ASAP7_75t_R g657 ( 
.A(n_624),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_504),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_523),
.B(n_191),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_509),
.B(n_191),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_533),
.B(n_298),
.Y(n_662)
);

NOR2x1p5_ASAP7_75t_L g663 ( 
.A(n_501),
.B(n_193),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_502),
.B(n_322),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_563),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_629),
.B(n_192),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_522),
.A2(n_310),
.B1(n_205),
.B2(n_286),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_522),
.A2(n_395),
.B1(n_207),
.B2(n_204),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_543),
.B(n_192),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_511),
.B(n_438),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_503),
.A2(n_205),
.B1(n_206),
.B2(n_286),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_506),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_582),
.Y(n_673)
);

OR2x6_ASAP7_75t_L g674 ( 
.A(n_620),
.B(n_383),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_505),
.B(n_194),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_508),
.B(n_194),
.Y(n_676)
);

INVx6_ASAP7_75t_L g677 ( 
.A(n_514),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_517),
.B(n_442),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_540),
.A2(n_206),
.B1(n_289),
.B2(n_295),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_516),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_582),
.Y(n_681)
);

O2A1O1Ixp5_ASAP7_75t_L g682 ( 
.A1(n_539),
.A2(n_449),
.B(n_446),
.C(n_391),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_596),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_629),
.B(n_196),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_542),
.B(n_446),
.Y(n_685)
);

BUFx6f_ASAP7_75t_SL g686 ( 
.A(n_566),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_620),
.B(n_385),
.Y(n_687)
);

OR2x6_ASAP7_75t_L g688 ( 
.A(n_635),
.B(n_385),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_196),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_503),
.A2(n_289),
.B1(n_295),
.B2(n_296),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_506),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_608),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_516),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_580),
.B(n_198),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_593),
.B(n_609),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_521),
.A2(n_388),
.B(n_290),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_SL g698 ( 
.A1(n_560),
.A2(n_300),
.B1(n_252),
.B2(n_296),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_589),
.B(n_599),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_526),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_526),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_638),
.B(n_388),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_539),
.A2(n_536),
.B1(n_527),
.B2(n_550),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_596),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_518),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_535),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_500),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_600),
.A2(n_309),
.B1(n_302),
.B2(n_304),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_501),
.B(n_203),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_535),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_580),
.B(n_207),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_594),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_512),
.B(n_285),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_612),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_622),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_574),
.B(n_290),
.Y(n_716)
);

AND2x6_ASAP7_75t_SL g717 ( 
.A(n_619),
.B(n_360),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_614),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_594),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_537),
.B(n_291),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_534),
.B(n_291),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_534),
.B(n_301),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_637),
.A2(n_363),
.B(n_360),
.C(n_301),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_615),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_601),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_617),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_558),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_618),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_631),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_601),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_512),
.B(n_303),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_528),
.B(n_303),
.Y(n_733)
);

AO22x1_ASAP7_75t_L g734 ( 
.A1(n_575),
.A2(n_302),
.B1(n_313),
.B2(n_315),
.Y(n_734)
);

OAI221xp5_ASAP7_75t_L g735 ( 
.A1(n_536),
.A2(n_595),
.B1(n_588),
.B2(n_587),
.C(n_571),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_626),
.B(n_300),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_627),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_574),
.B(n_314),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_632),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_528),
.B(n_314),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_571),
.B(n_321),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_574),
.B(n_321),
.Y(n_742)
);

O2A1O1Ixp5_ASAP7_75t_L g743 ( 
.A1(n_545),
.A2(n_363),
.B(n_300),
.C(n_329),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_530),
.B(n_329),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_530),
.B(n_224),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_532),
.B(n_228),
.Y(n_746)
);

OAI221xp5_ASAP7_75t_L g747 ( 
.A1(n_595),
.A2(n_335),
.B1(n_230),
.B2(n_239),
.C(n_241),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_546),
.B(n_244),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_603),
.B(n_246),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_636),
.B(n_515),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_581),
.B(n_247),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_515),
.B(n_253),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_640),
.B(n_259),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_635),
.B(n_3),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_585),
.B(n_92),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_640),
.B(n_265),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_642),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_548),
.B(n_280),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_641),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_569),
.B(n_328),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_606),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_603),
.B(n_328),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_641),
.A2(n_327),
.B1(n_326),
.B2(n_323),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_587),
.B(n_327),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_556),
.B(n_326),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_562),
.B(n_323),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_567),
.B(n_320),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_565),
.B(n_320),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_611),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_600),
.A2(n_318),
.B1(n_315),
.B2(n_313),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_579),
.B(n_318),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_510),
.B(n_5),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_165),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_538),
.B(n_162),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_551),
.B(n_155),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_551),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_567),
.B(n_5),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_549),
.B(n_8),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_527),
.A2(n_9),
.B1(n_15),
.B2(n_21),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_639),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_567),
.B(n_15),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_627),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_555),
.B(n_21),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_507),
.B(n_138),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_550),
.B(n_25),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_600),
.A2(n_127),
.B1(n_122),
.B2(n_115),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_598),
.B(n_26),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_616),
.Y(n_789)
);

NOR2x1p5_ASAP7_75t_L g790 ( 
.A(n_544),
.B(n_27),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_507),
.B(n_101),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_785),
.A2(n_735),
.B(n_696),
.C(n_669),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_728),
.B(n_633),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_789),
.A2(n_750),
.B(n_751),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_648),
.B(n_583),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_751),
.A2(n_581),
.B(n_597),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_693),
.B(n_652),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_705),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_741),
.B(n_633),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_741),
.B(n_575),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_695),
.B(n_513),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_583),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_699),
.A2(n_581),
.B(n_597),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_658),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_680),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_779),
.A2(n_610),
.B1(n_527),
.B2(n_547),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_682),
.A2(n_577),
.B(n_568),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_680),
.B(n_566),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_680),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_675),
.B(n_588),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_675),
.A2(n_676),
.B1(n_749),
.B2(n_677),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_676),
.B(n_586),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_702),
.B(n_573),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_716),
.A2(n_572),
.B(n_570),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_695),
.B(n_586),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_711),
.B(n_607),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_658),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_669),
.A2(n_711),
.B(n_645),
.C(n_653),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_651),
.B(n_607),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_738),
.A2(n_578),
.B(n_623),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_779),
.A2(n_547),
.B1(n_576),
.B2(n_519),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_738),
.A2(n_554),
.B(n_625),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_703),
.A2(n_749),
.B1(n_764),
.B2(n_671),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_692),
.B(n_573),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_707),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_742),
.A2(n_554),
.B(n_576),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_661),
.B(n_557),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_644),
.B(n_531),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_742),
.A2(n_639),
.B(n_630),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_661),
.B(n_665),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_659),
.B(n_660),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_659),
.B(n_660),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_680),
.B(n_573),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_693),
.B(n_634),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_666),
.B(n_604),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_773),
.A2(n_628),
.B(n_592),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_654),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_703),
.B(n_736),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_SL g839 ( 
.A1(n_774),
.A2(n_630),
.B(n_553),
.C(n_499),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_753),
.A2(n_592),
.B(n_628),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_654),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_677),
.A2(n_621),
.B1(n_619),
.B2(n_613),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_670),
.A2(n_557),
.B(n_559),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_677),
.A2(n_619),
.B1(n_624),
.B2(n_559),
.Y(n_844)
);

BUFx4f_ASAP7_75t_L g845 ( 
.A(n_674),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_756),
.A2(n_628),
.B(n_592),
.Y(n_846)
);

O2A1O1Ixp5_ASAP7_75t_L g847 ( 
.A1(n_664),
.A2(n_637),
.B(n_553),
.C(n_541),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_684),
.B(n_668),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_650),
.B(n_602),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_673),
.B(n_553),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_646),
.B(n_525),
.C(n_31),
.Y(n_851)
);

NOR2x1_ASAP7_75t_R g852 ( 
.A(n_643),
.B(n_27),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_672),
.A2(n_553),
.B(n_541),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_658),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_649),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_681),
.B(n_553),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_772),
.A2(n_564),
.B(n_499),
.C(n_33),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_683),
.A2(n_564),
.B1(n_499),
.B2(n_541),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_745),
.A2(n_541),
.B(n_100),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_694),
.B(n_541),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_704),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_746),
.B(n_34),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_672),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_715),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_713),
.A2(n_97),
.B(n_95),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_714),
.A2(n_739),
.B1(n_730),
.B2(n_729),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_748),
.B(n_746),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_718),
.B(n_37),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_691),
.A2(n_93),
.B(n_75),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_732),
.A2(n_73),
.B(n_70),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_725),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_691),
.A2(n_68),
.B(n_60),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_733),
.A2(n_37),
.B(n_38),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_715),
.B(n_40),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_700),
.A2(n_42),
.B(n_45),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_727),
.B(n_46),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_740),
.A2(n_46),
.B(n_47),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_656),
.B(n_49),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_698),
.B(n_52),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_652),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_776),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_662),
.B(n_57),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_744),
.A2(n_791),
.B(n_784),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_709),
.B(n_679),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_752),
.A2(n_721),
.B1(n_722),
.B2(n_761),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_686),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_708),
.B(n_720),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_701),
.A2(n_780),
.B(n_757),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_769),
.B(n_737),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_678),
.A2(n_685),
.B(n_775),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_706),
.A2(n_757),
.B(n_731),
.Y(n_891)
);

AO21x1_ASAP7_75t_L g892 ( 
.A1(n_786),
.A2(n_723),
.B(n_762),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_655),
.A2(n_689),
.B(n_712),
.Y(n_893)
);

OAI321xp33_ASAP7_75t_L g894 ( 
.A1(n_667),
.A2(n_770),
.A3(n_690),
.B1(n_671),
.B2(n_763),
.C(n_747),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_706),
.A2(n_724),
.B(n_731),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_710),
.B(n_782),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_767),
.A2(n_781),
.B(n_777),
.C(n_743),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_712),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_667),
.B(n_688),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_719),
.A2(n_726),
.B(n_724),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_719),
.Y(n_901)
);

AOI21x1_ASAP7_75t_L g902 ( 
.A1(n_726),
.A2(n_780),
.B(n_766),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_674),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_765),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_768),
.B(n_771),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_767),
.B(n_781),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_697),
.A2(n_755),
.B(n_758),
.Y(n_907)
);

CKINVDCx10_ASAP7_75t_R g908 ( 
.A(n_754),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_777),
.Y(n_909)
);

OAI321xp33_ASAP7_75t_L g910 ( 
.A1(n_690),
.A2(n_759),
.A3(n_778),
.B1(n_783),
.B2(n_754),
.C(n_788),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_674),
.A2(n_687),
.B(n_688),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_647),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_687),
.B(n_688),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_760),
.B(n_787),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_754),
.A2(n_687),
.B(n_788),
.C(n_663),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_717),
.B(n_734),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_790),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_788),
.B(n_657),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_658),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_693),
.B(n_652),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_648),
.B(n_529),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_682),
.A2(n_789),
.B(n_751),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_648),
.B(n_529),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_749),
.A2(n_711),
.B(n_695),
.C(n_648),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_703),
.A2(n_735),
.B1(n_665),
.B2(n_661),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_702),
.B(n_728),
.Y(n_926)
);

AO21x1_ASAP7_75t_L g927 ( 
.A1(n_749),
.A2(n_539),
.B(n_695),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_648),
.B(n_529),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_749),
.A2(n_711),
.B(n_695),
.C(n_648),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_648),
.B(n_529),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_789),
.A2(n_521),
.B(n_750),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_789),
.A2(n_521),
.B(n_750),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_749),
.A2(n_711),
.B(n_695),
.C(n_648),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_789),
.A2(n_521),
.B(n_750),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_696),
.B(n_646),
.C(n_785),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_648),
.B(n_529),
.Y(n_936)
);

OAI321xp33_ASAP7_75t_L g937 ( 
.A1(n_785),
.A2(n_550),
.A3(n_450),
.B1(n_708),
.B2(n_779),
.C(n_711),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_728),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_696),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_785),
.A2(n_779),
.B1(n_735),
.B2(n_522),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_728),
.B(n_569),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_658),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_789),
.A2(n_521),
.B(n_750),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_648),
.B(n_529),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_648),
.B(n_529),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_702),
.B(n_728),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_728),
.B(n_626),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_785),
.A2(n_779),
.B1(n_735),
.B2(n_522),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_682),
.A2(n_789),
.B(n_751),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_789),
.A2(n_521),
.B(n_750),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_648),
.B(n_529),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_785),
.A2(n_735),
.B(n_539),
.C(n_696),
.Y(n_952)
);

OAI22x1_ASAP7_75t_L g953 ( 
.A1(n_800),
.A2(n_799),
.B1(n_801),
.B2(n_832),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_891),
.Y(n_955)
);

INVx6_ASAP7_75t_L g956 ( 
.A(n_886),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_832),
.B(n_831),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_825),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_938),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_940),
.A2(n_948),
.B(n_933),
.C(n_929),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_924),
.A2(n_823),
.B1(n_940),
.B2(n_948),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_926),
.B(n_946),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_794),
.A2(n_803),
.B(n_830),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_925),
.A2(n_812),
.B(n_820),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_938),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_799),
.A2(n_800),
.B(n_848),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_871),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_921),
.B(n_923),
.Y(n_968)
);

NOR2x1_ASAP7_75t_SL g969 ( 
.A(n_864),
.B(n_809),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_928),
.B(n_930),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_797),
.B(n_920),
.Y(n_971)
);

OAI21x1_ASAP7_75t_L g972 ( 
.A1(n_869),
.A2(n_949),
.B(n_922),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_889),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_888),
.A2(n_900),
.B(n_895),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_936),
.B(n_944),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_945),
.B(n_951),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_886),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_901),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_931),
.A2(n_934),
.B(n_932),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_867),
.B(n_904),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_823),
.B(n_905),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_864),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_795),
.B(n_802),
.Y(n_983)
);

AO31x2_ASAP7_75t_L g984 ( 
.A1(n_927),
.A2(n_892),
.A3(n_862),
.B(n_897),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_837),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_829),
.A2(n_836),
.B(n_840),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_943),
.A2(n_950),
.B(n_819),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_814),
.A2(n_822),
.B(n_821),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_810),
.A2(n_952),
.B(n_792),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_848),
.A2(n_937),
.B(n_862),
.C(n_894),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_903),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_811),
.B(n_939),
.Y(n_992)
);

AOI21x1_ASAP7_75t_SL g993 ( 
.A1(n_878),
.A2(n_882),
.B(n_849),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_939),
.B(n_793),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_846),
.A2(n_847),
.B(n_807),
.Y(n_995)
);

OAI21x1_ASAP7_75t_SL g996 ( 
.A1(n_875),
.A2(n_872),
.B(n_907),
.Y(n_996)
);

AND3x4_ASAP7_75t_L g997 ( 
.A(n_851),
.B(n_935),
.C(n_947),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_827),
.A2(n_826),
.B(n_896),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_909),
.B(n_855),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_818),
.A2(n_838),
.B(n_847),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_861),
.A2(n_877),
.A3(n_873),
.B(n_876),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_935),
.A2(n_887),
.B1(n_906),
.B2(n_835),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_813),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_841),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_797),
.B(n_920),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_941),
.B(n_909),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_912),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_850),
.A2(n_856),
.B(n_860),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_863),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_866),
.B(n_885),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_839),
.A2(n_809),
.B(n_805),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_806),
.B(n_910),
.C(n_835),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_805),
.A2(n_898),
.B(n_884),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_806),
.A2(n_828),
.B(n_879),
.C(n_851),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_881),
.A2(n_853),
.B(n_865),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_899),
.B(n_824),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_804),
.B(n_942),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_804),
.B(n_942),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_868),
.B(n_804),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_804),
.B(n_942),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_870),
.A2(n_859),
.B(n_858),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_898),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_817),
.B(n_942),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_824),
.B(n_914),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_898),
.A2(n_864),
.B(n_808),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_857),
.A2(n_911),
.B(n_833),
.Y(n_1026)
);

AO21x1_ASAP7_75t_L g1027 ( 
.A1(n_874),
.A2(n_880),
.B(n_842),
.Y(n_1027)
);

AOI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_916),
.A2(n_915),
.B(n_914),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_834),
.A2(n_913),
.B(n_844),
.Y(n_1029)
);

BUFx4_ASAP7_75t_SL g1030 ( 
.A(n_917),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_898),
.A2(n_918),
.B(n_864),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_817),
.A2(n_919),
.B(n_854),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_845),
.A2(n_852),
.B(n_908),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_940),
.A2(n_948),
.B(n_924),
.C(n_933),
.Y(n_1034)
);

CKINVDCx11_ASAP7_75t_R g1035 ( 
.A(n_886),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_804),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_938),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_832),
.B(n_831),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_799),
.B(n_525),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_924),
.A2(n_929),
.B1(n_933),
.B2(n_823),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_832),
.B(n_831),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_800),
.B(n_855),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_804),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_924),
.A2(n_929),
.B1(n_933),
.B2(n_823),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_864),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_797),
.B(n_920),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_832),
.B(n_831),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_798),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_797),
.B(n_920),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_924),
.A2(n_933),
.B(n_929),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_SL g1055 ( 
.A(n_924),
.B(n_933),
.C(n_929),
.Y(n_1055)
);

OA21x2_ASAP7_75t_L g1056 ( 
.A1(n_927),
.A2(n_949),
.B(n_922),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_SL g1057 ( 
.A1(n_952),
.A2(n_792),
.B(n_875),
.Y(n_1057)
);

AOI221x1_ASAP7_75t_L g1058 ( 
.A1(n_924),
.A2(n_929),
.B1(n_933),
.B2(n_832),
.C(n_862),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_801),
.B(n_926),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_825),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_800),
.A2(n_450),
.B(n_832),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_891),
.A2(n_843),
.B(n_902),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_940),
.A2(n_948),
.B(n_924),
.C(n_933),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_924),
.A2(n_933),
.B(n_929),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_843),
.A2(n_891),
.B(n_902),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_891),
.A2(n_843),
.B(n_902),
.Y(n_1068)
);

AND2x2_ASAP7_75t_SL g1069 ( 
.A(n_940),
.B(n_948),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_924),
.B(n_929),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_832),
.B(n_831),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_809),
.B(n_854),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_832),
.B(n_831),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_864),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_797),
.B(n_920),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_800),
.B(n_855),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_843),
.A2(n_891),
.B(n_902),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_864),
.Y(n_1081)
);

AOI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_832),
.A2(n_799),
.B(n_800),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_SL g1083 ( 
.A1(n_831),
.A2(n_816),
.B(n_815),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_864),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_941),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_891),
.A2(n_843),
.B(n_893),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_940),
.A2(n_948),
.B(n_924),
.C(n_933),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_883),
.A2(n_890),
.B(n_796),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_832),
.B(n_831),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_864),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_832),
.B(n_831),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_924),
.A2(n_933),
.B(n_929),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_957),
.B(n_1039),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_967),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1082),
.B(n_1063),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_971),
.B(n_1005),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_994),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1043),
.B(n_1051),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_982),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_1061),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_SL g1101 ( 
.A1(n_953),
.A2(n_1079),
.B(n_1044),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_958),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1089),
.B(n_1091),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_971),
.B(n_1005),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1069),
.A2(n_990),
.B1(n_1012),
.B2(n_961),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_1035),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_1042),
.A2(n_1046),
.A3(n_1058),
.B(n_990),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_954),
.A2(n_1060),
.B(n_1050),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_970),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_971),
.B(n_1005),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_985),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1070),
.A2(n_1088),
.B(n_1073),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1052),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_1007),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_1002),
.A2(n_1012),
.B(n_975),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_976),
.B(n_983),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1059),
.B(n_962),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1035),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_981),
.B(n_1069),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_965),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_1054),
.A2(n_1092),
.B(n_1066),
.C(n_1071),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_965),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_992),
.B(n_973),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_978),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_960),
.A2(n_1065),
.B(n_1087),
.C(n_1034),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1003),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1004),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_960),
.B(n_1034),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1004),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_979),
.A2(n_987),
.B(n_964),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1009),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_991),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1038),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1038),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_959),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_999),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1049),
.B(n_1053),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_1085),
.B(n_1024),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1065),
.A2(n_1087),
.B1(n_1014),
.B2(n_1010),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1090),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1049),
.B(n_1053),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_955),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_SL g1145 ( 
.A1(n_1040),
.A2(n_1016),
.B1(n_1006),
.B2(n_980),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1090),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1085),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_1090),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1030),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_988),
.A2(n_1071),
.B(n_963),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_999),
.B(n_1014),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1029),
.B(n_1049),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_989),
.B(n_1055),
.Y(n_1153)
);

AOI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_1057),
.A2(n_1000),
.B(n_1027),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1055),
.A2(n_998),
.B(n_1008),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1053),
.B(n_1078),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1019),
.B(n_984),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_997),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_1078),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1078),
.B(n_1031),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_969),
.B(n_1022),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1030),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_984),
.B(n_1022),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_977),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_996),
.A2(n_1017),
.B(n_972),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1017),
.A2(n_972),
.B(n_974),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1047),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1036),
.B(n_1045),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_984),
.B(n_1013),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_995),
.A2(n_1056),
.B(n_1015),
.Y(n_1170)
);

OR2x6_ASAP7_75t_L g1171 ( 
.A(n_956),
.B(n_977),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1047),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1018),
.A2(n_1023),
.B(n_1020),
.C(n_997),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_1033),
.A2(n_1025),
.B1(n_1011),
.B2(n_1018),
.C(n_1023),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1076),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_956),
.B(n_1074),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1001),
.B(n_984),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1076),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1001),
.B(n_1084),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1036),
.B(n_1045),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1056),
.A2(n_1021),
.B(n_986),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1001),
.B(n_1084),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_956),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1090),
.Y(n_1184)
);

INVx8_ASAP7_75t_L g1185 ( 
.A(n_1081),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1186)
);

O2A1O1Ixp5_ASAP7_75t_L g1187 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1068),
.C(n_1083),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1056),
.A2(n_1074),
.B1(n_1001),
.B2(n_993),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1037),
.A2(n_1077),
.B(n_1041),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_SL g1190 ( 
.A(n_993),
.B(n_1048),
.C(n_1062),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1067),
.B(n_1080),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1086),
.A2(n_972),
.B(n_1000),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_967),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_954),
.A2(n_1060),
.B(n_1050),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1082),
.B(n_1063),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1061),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_982),
.Y(n_1197)
);

BUFx2_ASAP7_75t_SL g1198 ( 
.A(n_958),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_967),
.Y(n_1199)
);

NAND2x1p5_ASAP7_75t_L g1200 ( 
.A(n_971),
.B(n_809),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_966),
.A2(n_800),
.B1(n_799),
.B2(n_832),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_957),
.B(n_1039),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_971),
.B(n_1005),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_L g1204 ( 
.A(n_1012),
.B(n_924),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1061),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_971),
.B(n_809),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_957),
.B(n_1039),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1063),
.A2(n_799),
.B1(n_800),
.B2(n_832),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1061),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_971),
.B(n_809),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_1035),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1035),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1067),
.A2(n_1080),
.B(n_1068),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_966),
.A2(n_924),
.B(n_933),
.C(n_929),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_982),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1063),
.A2(n_799),
.B1(n_800),
.B2(n_832),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_966),
.A2(n_924),
.B(n_933),
.C(n_929),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1044),
.B(n_1079),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_967),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1035),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1069),
.A2(n_948),
.B1(n_940),
.B2(n_823),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_982),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_971),
.B(n_1005),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_985),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_956),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_990),
.A2(n_1034),
.B(n_960),
.Y(n_1226)
);

HAxp5_ASAP7_75t_L g1227 ( 
.A(n_1030),
.B(n_621),
.CON(n_1227),
.SN(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1061),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_982),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_954),
.A2(n_1060),
.B(n_1050),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1061),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_966),
.A2(n_924),
.B(n_933),
.C(n_929),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_967),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1082),
.B(n_1063),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_985),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1061),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1231),
.Y(n_1237)
);

BUFx8_ASAP7_75t_SL g1238 ( 
.A(n_1107),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1144),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1134),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1201),
.A2(n_1216),
.B(n_1208),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1158),
.A2(n_1221),
.B1(n_1097),
.B2(n_1195),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1184),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1121),
.Y(n_1244)
);

AO21x1_ASAP7_75t_L g1245 ( 
.A1(n_1221),
.A2(n_1217),
.B(n_1214),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1112),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1151),
.A2(n_1110),
.B1(n_1104),
.B2(n_1093),
.Y(n_1247)
);

INVx6_ASAP7_75t_L g1248 ( 
.A(n_1184),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1123),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1130),
.Y(n_1250)
);

OR2x6_ASAP7_75t_L g1251 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1211),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1095),
.B(n_1234),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1190),
.A2(n_1113),
.B(n_1109),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1225),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1110),
.A2(n_1117),
.B1(n_1104),
.B2(n_1098),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1204),
.A2(n_1116),
.B1(n_1106),
.B2(n_1145),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1117),
.A2(n_1093),
.B1(n_1202),
.B2(n_1098),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1120),
.B(n_1226),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_R g1260 ( 
.A(n_1212),
.B(n_1119),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1225),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1155),
.A2(n_1150),
.B(n_1131),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1220),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1106),
.A2(n_1141),
.B1(n_1153),
.B2(n_1226),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1183),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1164),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1176),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1114),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1120),
.B(n_1124),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1127),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1102),
.A2(n_1207),
.B1(n_1202),
.B2(n_1137),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1193),
.Y(n_1272)
);

BUFx4f_ASAP7_75t_SL g1273 ( 
.A(n_1196),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1115),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1199),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1149),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1155),
.A2(n_1181),
.B(n_1170),
.Y(n_1277)
);

BUFx10_ASAP7_75t_L g1278 ( 
.A(n_1140),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1102),
.B(n_1207),
.Y(n_1279)
);

NAND2x1p5_ASAP7_75t_L g1280 ( 
.A(n_1179),
.B(n_1182),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1124),
.B(n_1126),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1219),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1223),
.B(n_1096),
.Y(n_1283)
);

NAND2x1p5_ASAP7_75t_L g1284 ( 
.A(n_1186),
.B(n_1160),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1157),
.B(n_1108),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1233),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1223),
.B(n_1096),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1160),
.B(n_1177),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1141),
.A2(n_1129),
.B1(n_1135),
.B2(n_1100),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1125),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1209),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1118),
.B(n_1218),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1132),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1198),
.A2(n_1129),
.B1(n_1147),
.B2(n_1228),
.Y(n_1294)
);

INVxp33_ASAP7_75t_L g1295 ( 
.A(n_1103),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1223),
.B(n_1105),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1161),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1162),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1176),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1171),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1192),
.B(n_1191),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1128),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1224),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1235),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1163),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1138),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1154),
.A2(n_1205),
.B1(n_1100),
.B2(n_1159),
.Y(n_1307)
);

INVx4_ASAP7_75t_L g1308 ( 
.A(n_1176),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1108),
.B(n_1122),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1115),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1133),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1101),
.A2(n_1236),
.B1(n_1136),
.B2(n_1171),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_1171),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1189),
.A2(n_1166),
.B(n_1165),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_1230),
.B(n_1194),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1232),
.A2(n_1173),
.B1(n_1111),
.B2(n_1174),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1178),
.Y(n_1317)
);

OAI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1111),
.A2(n_1154),
.B1(n_1210),
.B2(n_1206),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1167),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1172),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1156),
.A2(n_1105),
.B1(n_1143),
.B2(n_1203),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1139),
.A2(n_1143),
.B1(n_1203),
.B2(n_1157),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1175),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1099),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1108),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1139),
.A2(n_1161),
.B1(n_1210),
.B2(n_1206),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1169),
.B(n_1099),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1185),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1188),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1185),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1187),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1192),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1142),
.B(n_1148),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1200),
.A2(n_1180),
.B1(n_1168),
.B2(n_1222),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1229),
.A2(n_1227),
.B1(n_1222),
.B2(n_1148),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1215),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1138),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1146),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1197),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1220),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1134),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1097),
.B(n_1151),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1155),
.A2(n_1150),
.B(n_1131),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1103),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1201),
.A2(n_966),
.B1(n_799),
.B2(n_800),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1094),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1225),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_1184),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1094),
.Y(n_1349)
);

BUFx2_ASAP7_75t_R g1350 ( 
.A(n_1119),
.Y(n_1350)
);

CKINVDCx8_ASAP7_75t_R g1351 ( 
.A(n_1198),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1225),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1231),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1120),
.B(n_1153),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1115),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1285),
.B(n_1354),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1245),
.A2(n_1329),
.A3(n_1331),
.B(n_1325),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1292),
.B(n_1253),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1288),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1267),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1240),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1242),
.B(n_1345),
.C(n_1257),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1259),
.B(n_1280),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1342),
.B(n_1256),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1251),
.B(n_1267),
.Y(n_1365)
);

INVx5_ASAP7_75t_L g1366 ( 
.A(n_1267),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1285),
.B(n_1354),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1240),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1332),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1259),
.B(n_1280),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1305),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1270),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1309),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1309),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1327),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1239),
.Y(n_1376)
);

AO21x2_ASAP7_75t_L g1377 ( 
.A1(n_1314),
.A2(n_1315),
.B(n_1254),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1267),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1251),
.B(n_1342),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1301),
.A2(n_1277),
.B(n_1262),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1301),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1301),
.A2(n_1277),
.B(n_1262),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1279),
.B(n_1258),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1313),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1251),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1241),
.A2(n_1253),
.B(n_1316),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1251),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1302),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1288),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1288),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1284),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1269),
.B(n_1281),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1269),
.B(n_1281),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1268),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1272),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1341),
.Y(n_1396)
);

INVx2_ASAP7_75t_SL g1397 ( 
.A(n_1313),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1275),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1282),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1254),
.A2(n_1318),
.B(n_1247),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1286),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1244),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1312),
.A2(n_1349),
.B(n_1346),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1290),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1262),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1299),
.B(n_1308),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1293),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1317),
.A2(n_1335),
.B(n_1271),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1307),
.B(n_1343),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1264),
.A2(n_1322),
.B1(n_1294),
.B2(n_1321),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1297),
.B(n_1246),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1340),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1297),
.B(n_1250),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1238),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1341),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1244),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1297),
.A2(n_1304),
.B(n_1303),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1289),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1274),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1299),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1324),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1336),
.A2(n_1333),
.B(n_1319),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1337),
.A2(n_1338),
.B(n_1320),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1308),
.Y(n_1424)
);

NOR4xp25_ASAP7_75t_SL g1425 ( 
.A(n_1414),
.B(n_1252),
.C(n_1263),
.D(n_1330),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1356),
.B(n_1310),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1356),
.B(n_1291),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1367),
.B(n_1373),
.Y(n_1428)
);

INVx2_ASAP7_75t_SL g1429 ( 
.A(n_1391),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1381),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1373),
.B(n_1278),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1369),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1372),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1388),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1362),
.A2(n_1351),
.B1(n_1355),
.B2(n_1300),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1374),
.B(n_1375),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1375),
.B(n_1278),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1367),
.B(n_1291),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1381),
.B(n_1296),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1381),
.B(n_1323),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1383),
.B(n_1249),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1410),
.A2(n_1351),
.B1(n_1353),
.B2(n_1237),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1366),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1386),
.A2(n_1344),
.B1(n_1295),
.B2(n_1311),
.C(n_1298),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1377),
.A2(n_1296),
.B(n_1283),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1363),
.B(n_1370),
.Y(n_1446)
);

CKINVDCx16_ASAP7_75t_R g1447 ( 
.A(n_1412),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1409),
.B(n_1311),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1364),
.B(n_1295),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1363),
.B(n_1296),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1409),
.B(n_1287),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1358),
.B(n_1273),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1371),
.B(n_1326),
.Y(n_1453)
);

HB1xp67_ASAP7_75t_L g1454 ( 
.A(n_1422),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1392),
.B(n_1270),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1422),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1405),
.B(n_1306),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1379),
.B(n_1265),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1422),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1417),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1392),
.B(n_1298),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1379),
.B(n_1265),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1444),
.B(n_1442),
.C(n_1435),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1419),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1444),
.B(n_1418),
.C(n_1442),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

OAI221xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1435),
.A2(n_1418),
.B1(n_1387),
.B2(n_1385),
.C(n_1365),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1441),
.A2(n_1415),
.B1(n_1396),
.B2(n_1368),
.C(n_1361),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1449),
.B(n_1416),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1426),
.B(n_1402),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1452),
.A2(n_1393),
.B(n_1378),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1453),
.A2(n_1402),
.B1(n_1393),
.B2(n_1387),
.C(n_1385),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1453),
.B(n_1399),
.C(n_1407),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1446),
.B(n_1436),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1434),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1448),
.A2(n_1365),
.B1(n_1406),
.B2(n_1389),
.C(n_1390),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1426),
.B(n_1394),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1436),
.B(n_1400),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1461),
.A2(n_1378),
.B(n_1359),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1447),
.B(n_1378),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1451),
.B(n_1400),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1426),
.B(n_1395),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1455),
.A2(n_1365),
.B1(n_1378),
.B2(n_1408),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1427),
.B(n_1395),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1437),
.A2(n_1401),
.B1(n_1399),
.B2(n_1404),
.C(n_1398),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_L g1488 ( 
.A1(n_1448),
.A2(n_1260),
.B(n_1390),
.C(n_1263),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1425),
.B(n_1407),
.C(n_1404),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1431),
.B(n_1357),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1447),
.A2(n_1366),
.B1(n_1334),
.B2(n_1365),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1433),
.A2(n_1408),
.B1(n_1403),
.B2(n_1300),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1357),
.Y(n_1493)
);

OAI21xp33_ASAP7_75t_L g1494 ( 
.A1(n_1438),
.A2(n_1401),
.B(n_1398),
.Y(n_1494)
);

NAND3xp33_ASAP7_75t_L g1495 ( 
.A(n_1454),
.B(n_1424),
.C(n_1378),
.Y(n_1495)
);

OAI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1458),
.A2(n_1397),
.B1(n_1360),
.B2(n_1384),
.C(n_1252),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1437),
.B(n_1403),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1425),
.B(n_1421),
.C(n_1424),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1439),
.A2(n_1365),
.B1(n_1378),
.B2(n_1408),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1454),
.A2(n_1382),
.B(n_1380),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1440),
.B(n_1403),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1462),
.B(n_1376),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1462),
.A2(n_1360),
.B(n_1423),
.Y(n_1503)
);

NOR3xp33_ASAP7_75t_L g1504 ( 
.A(n_1443),
.B(n_1420),
.C(n_1397),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1456),
.B(n_1413),
.C(n_1411),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1460),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1477),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1501),
.B(n_1428),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1474),
.B(n_1443),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1480),
.B(n_1445),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1474),
.B(n_1459),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1469),
.B(n_1276),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1497),
.B(n_1428),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1475),
.B(n_1445),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1475),
.B(n_1483),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1500),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1445),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1484),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1470),
.B(n_1428),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1445),
.Y(n_1524)
);

AND2x2_ASAP7_75t_SL g1525 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1490),
.B(n_1357),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1493),
.B(n_1430),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1471),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1493),
.B(n_1357),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1486),
.B(n_1464),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1502),
.B(n_1457),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1494),
.B(n_1357),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1494),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1505),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1482),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1508),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_R g1538 ( 
.A(n_1516),
.B(n_1340),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1520),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1518),
.B(n_1492),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1525),
.B(n_1488),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1504),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1506),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1515),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1507),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1508),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1507),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1503),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1509),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1509),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1519),
.B(n_1450),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1534),
.B(n_1487),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1515),
.Y(n_1554)
);

NOR3x1_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1463),
.C(n_1465),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1520),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1533),
.B(n_1468),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1513),
.B(n_1495),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1524),
.B(n_1485),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1431),
.Y(n_1560)
);

INVxp33_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1463),
.B(n_1488),
.C(n_1481),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1533),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1531),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1508),
.B(n_1429),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1525),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1535),
.Y(n_1568)
);

NAND4xp25_ASAP7_75t_L g1569 ( 
.A(n_1532),
.B(n_1467),
.C(n_1473),
.D(n_1489),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1511),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1567),
.B(n_1508),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1568),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1537),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1539),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1539),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1537),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1539),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1544),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1567),
.B(n_1508),
.Y(n_1580)
);

NAND2x1_ASAP7_75t_L g1581 ( 
.A(n_1558),
.B(n_1527),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1569),
.B(n_1517),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1546),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1553),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1519),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1552),
.B(n_1519),
.Y(n_1587)
);

NAND2xp33_ASAP7_75t_L g1588 ( 
.A(n_1562),
.B(n_1535),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1472),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1557),
.B(n_1530),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_L g1591 ( 
.A(n_1557),
.B(n_1538),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1569),
.B(n_1517),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1555),
.B(n_1528),
.Y(n_1593)
);

NAND4xp75_ASAP7_75t_L g1594 ( 
.A(n_1555),
.B(n_1532),
.C(n_1521),
.D(n_1514),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1528),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1563),
.B(n_1512),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1568),
.B(n_1512),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1510),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1546),
.Y(n_1599)
);

NOR2x1_ASAP7_75t_L g1600 ( 
.A(n_1558),
.B(n_1498),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1560),
.B(n_1527),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1548),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1548),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1550),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1550),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1536),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1543),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1551),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1543),
.B(n_1510),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1543),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1551),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1564),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1559),
.B(n_1522),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1590),
.B(n_1559),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1578),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1581),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1588),
.A2(n_1545),
.B1(n_1554),
.B2(n_1559),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1600),
.B(n_1543),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1589),
.B(n_1540),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1590),
.B(n_1540),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1574),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1571),
.B(n_1545),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1589),
.B(n_1607),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1599),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1589),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1571),
.B(n_1540),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1575),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1613),
.B(n_1564),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1603),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1572),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1575),
.A2(n_1554),
.B(n_1556),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1579),
.B(n_1541),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1593),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1582),
.B(n_1592),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1571),
.B(n_1549),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1591),
.B(n_1238),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1610),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1580),
.B(n_1549),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1604),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1580),
.B(n_1586),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1580),
.B(n_1558),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1605),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1606),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1573),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1615),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1618),
.A2(n_1594),
.B1(n_1579),
.B2(n_1585),
.Y(n_1651)
);

OAI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1618),
.A2(n_1585),
.B1(n_1588),
.B2(n_1561),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1639),
.A2(n_1591),
.B(n_1596),
.C(n_1576),
.Y(n_1653)
);

AOI222xp33_ASAP7_75t_L g1654 ( 
.A1(n_1619),
.A2(n_1549),
.B1(n_1541),
.B2(n_1558),
.C1(n_1598),
.C2(n_1597),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1615),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1638),
.B(n_1541),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1638),
.B(n_1587),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1628),
.A2(n_1598),
.B1(n_1612),
.B2(n_1609),
.Y(n_1658)
);

AOI321xp33_ASAP7_75t_L g1659 ( 
.A1(n_1639),
.A2(n_1598),
.A3(n_1609),
.B1(n_1496),
.B2(n_1491),
.C(n_1478),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1635),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1641),
.A2(n_1266),
.B(n_1350),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

OAI22xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1628),
.A2(n_1606),
.B1(n_1609),
.B2(n_1536),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1625),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1614),
.A2(n_1526),
.B1(n_1529),
.B2(n_1601),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1624),
.Y(n_1670)
);

OAI32xp33_ASAP7_75t_L g1671 ( 
.A1(n_1614),
.A2(n_1529),
.A3(n_1526),
.B1(n_1570),
.B2(n_1536),
.Y(n_1671)
);

INVxp67_ASAP7_75t_L g1672 ( 
.A(n_1635),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1627),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1626),
.B(n_1266),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1616),
.B(n_1626),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1661),
.B(n_1642),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1670),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1672),
.B(n_1668),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1675),
.B(n_1620),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1670),
.B(n_1620),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1624),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1668),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1674),
.B(n_1621),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1652),
.A2(n_1616),
.B1(n_1637),
.B2(n_1646),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1669),
.B(n_1645),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1669),
.B(n_1645),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1653),
.A2(n_1646),
.B1(n_1629),
.B2(n_1643),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1658),
.B(n_1629),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1660),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1656),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1657),
.B(n_1646),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1651),
.B(n_1649),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_SL g1696 ( 
.A1(n_1695),
.A2(n_1659),
.B(n_1648),
.C(n_1663),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1687),
.A2(n_1654),
.B(n_1646),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1693),
.A2(n_1662),
.B1(n_1664),
.B2(n_1649),
.C(n_1634),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1684),
.B(n_1649),
.C(n_1665),
.Y(n_1699)
);

AOI21xp33_ASAP7_75t_L g1700 ( 
.A1(n_1686),
.A2(n_1673),
.B(n_1666),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1683),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1676),
.A2(n_1671),
.B1(n_1667),
.B2(n_1662),
.C(n_1627),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1679),
.A2(n_1647),
.B(n_1644),
.C(n_1631),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1691),
.A2(n_1640),
.B1(n_1643),
.B2(n_1648),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1690),
.A2(n_1640),
.B1(n_1634),
.B2(n_1632),
.Y(n_1705)
);

AOI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1691),
.A2(n_1647),
.B1(n_1644),
.B2(n_1631),
.C(n_1633),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1680),
.A2(n_1694),
.B(n_1689),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1699),
.B(n_1694),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1707),
.B(n_1680),
.Y(n_1709)
);

NOR3xp33_ASAP7_75t_L g1710 ( 
.A(n_1698),
.B(n_1681),
.C(n_1677),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1701),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1697),
.B(n_1678),
.Y(n_1712)
);

AOI211x1_ASAP7_75t_L g1713 ( 
.A1(n_1700),
.A2(n_1681),
.B(n_1682),
.C(n_1678),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_L g1714 ( 
.A(n_1696),
.B(n_1702),
.C(n_1706),
.Y(n_1714)
);

AND5x1_ASAP7_75t_L g1715 ( 
.A(n_1704),
.B(n_1688),
.C(n_1689),
.D(n_1682),
.E(n_1683),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1705),
.A2(n_1688),
.B(n_1685),
.Y(n_1716)
);

NOR2x1_ASAP7_75t_L g1717 ( 
.A(n_1703),
.B(n_1692),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1696),
.B(n_1692),
.C(n_1685),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1713),
.B(n_1633),
.Y(n_1719)
);

NAND4xp25_ASAP7_75t_L g1720 ( 
.A(n_1714),
.B(n_1632),
.C(n_1622),
.D(n_1630),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1622),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1708),
.B(n_1636),
.C(n_1623),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1718),
.A2(n_1622),
.B1(n_1630),
.B2(n_1623),
.C(n_1608),
.Y(n_1723)
);

NAND4xp25_ASAP7_75t_SL g1724 ( 
.A(n_1712),
.B(n_1630),
.C(n_1623),
.D(n_1611),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_L g1725 ( 
.A(n_1710),
.B(n_1636),
.C(n_1261),
.Y(n_1725)
);

NOR2x1_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1717),
.Y(n_1726)
);

AND3x4_ASAP7_75t_L g1727 ( 
.A(n_1725),
.B(n_1715),
.C(n_1716),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1721),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1719),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1723),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1720),
.Y(n_1731)
);

NAND4xp75_ASAP7_75t_L g1732 ( 
.A(n_1726),
.B(n_1711),
.C(n_1722),
.D(n_1577),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1728),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1727),
.B(n_1255),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1276),
.B1(n_1577),
.B2(n_1536),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1730),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1732),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1736),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1733),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1738),
.A2(n_1729),
.B1(n_1734),
.B2(n_1735),
.Y(n_1740)
);

AND3x1_ASAP7_75t_L g1741 ( 
.A(n_1740),
.B(n_1737),
.C(n_1739),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1737),
.B(n_1739),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1741),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1739),
.B(n_1261),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1743),
.A2(n_1347),
.B(n_1255),
.Y(n_1745)
);

AOI21xp33_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1352),
.B(n_1347),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1352),
.B1(n_1565),
.B2(n_1556),
.C(n_1570),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1746),
.A2(n_1747),
.B(n_1330),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_SL g1749 ( 
.A1(n_1748),
.A2(n_1547),
.B1(n_1556),
.B2(n_1248),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1749),
.A2(n_1339),
.B1(n_1547),
.B2(n_1566),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1328),
.B(n_1348),
.C(n_1243),
.Y(n_1751)
);


endmodule