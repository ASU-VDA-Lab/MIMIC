module fake_jpeg_3532_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_27),
.Y(n_47)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_34),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_29),
.B(n_33),
.C(n_31),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_27),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_27),
.B1(n_41),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_57),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_41),
.B1(n_34),
.B2(n_28),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_28),
.B1(n_36),
.B2(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_30),
.B1(n_26),
.B2(n_2),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_26),
.C(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_2),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_13),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_74),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_45),
.B1(n_14),
.B2(n_15),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_75),
.A2(n_4),
.B(n_6),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_3),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_24),
.C(n_22),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_83),
.B(n_7),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_82),
.B1(n_75),
.B2(n_8),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_6),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_71),
.A3(n_78),
.B1(n_69),
.B2(n_72),
.C(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_82),
.B(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_88),
.Y(n_92)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_17),
.B(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_19),
.Y(n_96)
);


endmodule