module real_jpeg_17616_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_50;
wire n_33;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_47;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_20),
.Y(n_31)
);

OR2x4_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_2),
.B(n_11),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_2),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_15),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_3),
.B(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_15),
.Y(n_16)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_37),
.C(n_39),
.Y(n_7)
);

INVxp67_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_17),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NAND3xp33_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_14),
.C(n_16),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_15),
.B(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_21),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_38),
.Y(n_37)
);

OR2x4_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_38),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);


endmodule