module fake_netlist_6_1626_n_1068 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1068);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1068;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1027;
wire n_875;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_184;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_964;
wire n_802;
wire n_831;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_970;
wire n_849;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_960;
wire n_841;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_18),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_31),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_75),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_14),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_26),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_38),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_93),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_81),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_90),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_116),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_8),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_137),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_17),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_67),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_136),
.Y(n_210)
);

BUFx8_ASAP7_75t_SL g211 ( 
.A(n_108),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_22),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_100),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_97),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_102),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_96),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_141),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_89),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_24),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_158),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_64),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_83),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_42),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_85),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_71),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_111),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_84),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_157),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_95),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_154),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_12),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_126),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_24),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_8),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_124),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_114),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_182),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_194),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_204),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_247),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_192),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_191),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_205),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_192),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_203),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_203),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_218),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_222),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_220),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_220),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_246),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_189),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_222),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_189),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_202),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_202),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_243),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_273),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_268),
.A2(n_296),
.B(n_223),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_243),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_256),
.B(n_186),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_245),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_223),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_187),
.Y(n_317)
);

CKINVDCx6p67_ASAP7_75t_R g318 ( 
.A(n_279),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_196),
.B(n_193),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_267),
.A2(n_198),
.B(n_197),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_254),
.B(n_187),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_281),
.A2(n_200),
.B(n_199),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_259),
.B(n_201),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_261),
.A2(n_244),
.B1(n_208),
.B2(n_240),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_206),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_287),
.B(n_248),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_257),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_251),
.B(n_214),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_244),
.B1(n_239),
.B2(n_237),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_289),
.C(n_291),
.Y(n_355)
);

BUFx6f_ASAP7_75t_SL g356 ( 
.A(n_348),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_303),
.B(n_336),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_301),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_349),
.B(n_270),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_290),
.Y(n_364)
);

INVxp67_ASAP7_75t_R g365 ( 
.A(n_321),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_351),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_348),
.B(n_290),
.Y(n_374)
);

NOR2x1p5_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_294),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_301),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_302),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_310),
.B(n_294),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_348),
.B(n_216),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_302),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_348),
.B(n_228),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_303),
.B(n_333),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_350),
.B(n_229),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_303),
.B(n_231),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_350),
.B(n_232),
.Y(n_393)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_350),
.B(n_234),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_319),
.Y(n_400)
);

OA22x2_ASAP7_75t_L g401 ( 
.A1(n_335),
.A2(n_354),
.B1(n_349),
.B2(n_303),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g404 ( 
.A(n_306),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_338),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_354),
.A2(n_236),
.B1(n_280),
.B2(n_265),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_333),
.B(n_310),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_350),
.B(n_265),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_343),
.B(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_352),
.B(n_280),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_211),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_343),
.B(n_211),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_352),
.B(n_353),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_369),
.Y(n_426)
);

XNOR2x2_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_288),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_367),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_353),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_387),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_383),
.B(n_353),
.Y(n_432)
);

OR2x6_ASAP7_75t_L g433 ( 
.A(n_375),
.B(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_382),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_306),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_399),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_417),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_346),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_408),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_304),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_352),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_366),
.B(n_324),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_369),
.B(n_308),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_394),
.B(n_308),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_394),
.B(n_344),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_404),
.B(n_347),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_416),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_419),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_327),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_419),
.Y(n_474)
);

NAND2x1p5_ASAP7_75t_L g475 ( 
.A(n_425),
.B(n_344),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_395),
.A2(n_316),
.B(n_326),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_424),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_385),
.B(n_345),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_421),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_402),
.B(n_345),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_385),
.B(n_344),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_370),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_370),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_371),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_422),
.B(n_344),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_402),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_371),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_402),
.Y(n_492)
);

AOI21x1_ASAP7_75t_L g493 ( 
.A1(n_395),
.A2(n_320),
.B(n_321),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_391),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_288),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_364),
.B(n_322),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_388),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_400),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_356),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_400),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_360),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_449),
.B(n_356),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_427),
.A2(n_410),
.B1(n_403),
.B2(n_356),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_472),
.A2(n_410),
.B1(n_403),
.B2(n_316),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_364),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_484),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_463),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_485),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_432),
.B(n_374),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_472),
.B(n_394),
.Y(n_516)
);

INVx8_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_374),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_499),
.B(n_380),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_451),
.B(n_410),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_430),
.B(n_390),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_452),
.B(n_355),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_473),
.B(n_390),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_393),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_468),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_426),
.B(n_393),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_481),
.B(n_426),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_470),
.B(n_397),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_498),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_429),
.B(n_397),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_322),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_316),
.B1(n_362),
.B2(n_384),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_448),
.B(n_380),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_461),
.B(n_347),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_434),
.B(n_409),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_489),
.Y(n_538)
);

INVx8_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_409),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_460),
.A2(n_365),
.B1(n_380),
.B2(n_384),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_454),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_436),
.B(n_409),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_439),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_455),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_440),
.B(n_361),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_503),
.A2(n_316),
.B1(n_362),
.B2(n_384),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_441),
.B(n_361),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_442),
.B(n_361),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_443),
.B(n_413),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_475),
.A2(n_372),
.B1(n_379),
.B2(n_378),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_447),
.B(n_413),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_492),
.B(n_326),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_495),
.B(n_413),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_450),
.B(n_372),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_477),
.B(n_339),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_457),
.A2(n_332),
.B1(n_320),
.B2(n_331),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_456),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_502),
.B(n_373),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_479),
.B(n_373),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_510),
.A2(n_474),
.B1(n_445),
.B2(n_444),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_528),
.B(n_483),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_507),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

AOI22x1_ASAP7_75t_L g574 ( 
.A1(n_542),
.A2(n_475),
.B1(n_476),
.B2(n_469),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_514),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_524),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_505),
.B(n_467),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_517),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_512),
.B(n_497),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_529),
.A2(n_474),
.B1(n_465),
.B2(n_483),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

AND2x6_ASAP7_75t_SL g583 ( 
.A(n_530),
.B(n_438),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_561),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_525),
.B(n_471),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_518),
.B(n_458),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_532),
.B(n_480),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_530),
.B(n_488),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_539),
.Y(n_592)
);

AO22x1_ASAP7_75t_L g593 ( 
.A1(n_535),
.A2(n_347),
.B1(n_446),
.B2(n_491),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_548),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_490),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_531),
.B(n_522),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_531),
.B(n_494),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_523),
.Y(n_601)
);

NOR3xp33_ASAP7_75t_SL g602 ( 
.A(n_535),
.B(n_313),
.C(n_347),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_526),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_527),
.B(n_496),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_515),
.A2(n_466),
.B1(n_476),
.B2(n_478),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

BUFx4_ASAP7_75t_SL g609 ( 
.A(n_511),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_547),
.B(n_331),
.Y(n_610)
);

CKINVDCx8_ASAP7_75t_R g611 ( 
.A(n_539),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_513),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_538),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_549),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_553),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_514),
.B(n_331),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_559),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_554),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_541),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_541),
.B(n_378),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_L g626 ( 
.A(n_541),
.B(n_379),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_508),
.B(n_340),
.C(n_337),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_543),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_574),
.A2(n_544),
.B(n_556),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_541),
.Y(n_630)
);

AOI221xp5_ASAP7_75t_L g631 ( 
.A1(n_601),
.A2(n_508),
.B1(n_563),
.B2(n_340),
.C(n_509),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_570),
.Y(n_632)
);

AOI21x1_ASAP7_75t_L g633 ( 
.A1(n_593),
.A2(n_516),
.B(n_568),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_581),
.A2(n_509),
.B1(n_520),
.B2(n_533),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_573),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_599),
.B(n_546),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_571),
.A2(n_516),
.B(n_534),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_626),
.A2(n_534),
.B(n_506),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_570),
.Y(n_639)
);

AND3x4_ASAP7_75t_L g640 ( 
.A(n_587),
.B(n_230),
.C(n_566),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_585),
.A2(n_506),
.B(n_560),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_558),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_606),
.A2(n_560),
.B(n_519),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_572),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_621),
.B(n_519),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_580),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_584),
.A2(n_550),
.B(n_533),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_607),
.A2(n_493),
.B(n_550),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_609),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_610),
.A2(n_563),
.B(n_337),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_622),
.Y(n_652)
);

BUFx6f_ASAP7_75t_SL g653 ( 
.A(n_570),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_620),
.A2(n_313),
.B(n_32),
.Y(n_654)
);

OAI21xp33_ASAP7_75t_L g655 ( 
.A1(n_569),
.A2(n_230),
.B(n_0),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_598),
.B(n_1),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_627),
.A2(n_314),
.B(n_33),
.Y(n_657)
);

CKINVDCx8_ASAP7_75t_R g658 ( 
.A(n_583),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_582),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_598),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_660)
);

AOI21xp33_ASAP7_75t_L g661 ( 
.A1(n_591),
.A2(n_4),
.B(n_5),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_588),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_587),
.A2(n_314),
.B1(n_7),
.B2(n_9),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_594),
.Y(n_665)
);

AOI221x1_ASAP7_75t_L g666 ( 
.A1(n_619),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_666)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_600),
.A2(n_617),
.B(n_618),
.C(n_624),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_612),
.B(n_10),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_624),
.A2(n_35),
.B(n_34),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_614),
.Y(n_670)
);

OAI21x1_ASAP7_75t_SL g671 ( 
.A1(n_628),
.A2(n_39),
.B(n_36),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_615),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_628),
.A2(n_45),
.B(n_41),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_616),
.B(n_11),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_604),
.B(n_13),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_608),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_575),
.A2(n_314),
.B(n_48),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_613),
.A2(n_49),
.B(n_47),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_589),
.A2(n_314),
.B(n_51),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_595),
.A2(n_314),
.B(n_52),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_605),
.B(n_13),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_596),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_589),
.A2(n_597),
.B(n_613),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_649),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_646),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_651),
.A2(n_597),
.B(n_613),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_648),
.A2(n_603),
.B(n_625),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_629),
.A2(n_625),
.B(n_602),
.Y(n_688)
);

AO22x2_ASAP7_75t_L g689 ( 
.A1(n_666),
.A2(n_578),
.B1(n_611),
.B2(n_625),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_661),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_690)
);

O2A1O1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_655),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_654),
.A2(n_625),
.B(n_623),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_647),
.A2(n_623),
.B(n_579),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_659),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_665),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_637),
.A2(n_19),
.A3(n_20),
.B(n_21),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_633),
.A2(n_579),
.B(n_576),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_644),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_635),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_641),
.A2(n_592),
.B(n_576),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_632),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_650),
.B(n_592),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_592),
.B(n_122),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_670),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_682),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_645),
.A2(n_21),
.B(n_23),
.C(n_25),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_653),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_676),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_SL g709 ( 
.A(n_640),
.B(n_26),
.C(n_27),
.Y(n_709)
);

O2A1O1Ixp5_ASAP7_75t_L g710 ( 
.A1(n_657),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_710)
);

O2A1O1Ixp33_ASAP7_75t_SL g711 ( 
.A1(n_667),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_681),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_SL g714 ( 
.A1(n_664),
.A2(n_30),
.B(n_31),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_658),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_50),
.Y(n_716)
);

BUFx2_ASAP7_75t_R g717 ( 
.A(n_630),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_672),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_674),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_643),
.A2(n_181),
.B(n_55),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_669),
.A2(n_54),
.B(n_56),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_642),
.Y(n_722)
);

OA21x2_ASAP7_75t_L g723 ( 
.A1(n_673),
.A2(n_57),
.B(n_58),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_653),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_675),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_636),
.B(n_656),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_680),
.A2(n_59),
.B(n_60),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_663),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_634),
.A2(n_66),
.B(n_68),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_677),
.A2(n_679),
.B(n_683),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_631),
.A2(n_180),
.B(n_70),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_645),
.A2(n_179),
.B(n_72),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_671),
.A2(n_69),
.B(n_74),
.Y(n_733)
);

AO31x2_ASAP7_75t_L g734 ( 
.A1(n_660),
.A2(n_639),
.A3(n_678),
.B(n_668),
.Y(n_734)
);

A2O1A1Ixp33_ASAP7_75t_L g735 ( 
.A1(n_632),
.A2(n_77),
.B(n_79),
.C(n_82),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_662),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_639),
.B(n_91),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_662),
.A2(n_92),
.B(n_94),
.C(n_99),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_662),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_632),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_649),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_639),
.B(n_101),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_648),
.A2(n_103),
.B(n_104),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_644),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_655),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_725),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_684),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_701),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_695),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_704),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_708),
.Y(n_751)
);

CKINVDCx11_ASAP7_75t_R g752 ( 
.A(n_724),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_715),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_714),
.A2(n_113),
.B1(n_115),
.B2(n_117),
.Y(n_754)
);

CKINVDCx11_ASAP7_75t_R g755 ( 
.A(n_724),
.Y(n_755)
);

INVx6_ASAP7_75t_L g756 ( 
.A(n_707),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_726),
.B(n_118),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_719),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_722),
.B(n_712),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_685),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_731),
.A2(n_128),
.B(n_129),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_701),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_701),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_709),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_764)
);

INVx8_ASAP7_75t_L g765 ( 
.A(n_702),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_699),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_744),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_694),
.B(n_138),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_740),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_702),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_689),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_741),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_698),
.Y(n_774)
);

BUFx4_ASAP7_75t_R g775 ( 
.A(n_717),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_705),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_713),
.Y(n_777)
);

BUFx2_ASAP7_75t_R g778 ( 
.A(n_739),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_696),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_745),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_740),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_706),
.A2(n_150),
.B(n_151),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_716),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_740),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_696),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_742),
.B(n_160),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_696),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_691),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_742),
.Y(n_789)
);

INVx6_ASAP7_75t_L g790 ( 
.A(n_700),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_687),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_697),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_SL g793 ( 
.A1(n_737),
.A2(n_723),
.B1(n_690),
.B2(n_711),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_735),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_723),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_720),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_693),
.Y(n_797)
);

INVx1_ASAP7_75t_SL g798 ( 
.A(n_686),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_734),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_736),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

INVx6_ASAP7_75t_L g802 ( 
.A(n_734),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_765),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_789),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_765),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_749),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_751),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_772),
.Y(n_809)
);

OAI21x1_ASAP7_75t_L g810 ( 
.A1(n_799),
.A2(n_688),
.B(n_730),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_789),
.B(n_729),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_797),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_779),
.Y(n_813)
);

OAI21x1_ASAP7_75t_L g814 ( 
.A1(n_801),
.A2(n_692),
.B(n_721),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_785),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_792),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_787),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_791),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_754),
.A2(n_710),
.B(n_728),
.C(n_738),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_790),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_802),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_802),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_773),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_750),
.B(n_733),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_759),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_777),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_774),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_798),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_790),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_767),
.Y(n_830)
);

BUFx8_ASAP7_75t_L g831 ( 
.A(n_766),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_795),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_752),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_795),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_793),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_760),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_780),
.A2(n_703),
.A3(n_732),
.B(n_727),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_768),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_748),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_762),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_770),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_757),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_789),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_753),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_763),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_763),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_761),
.A2(n_169),
.B(n_170),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

OAI21x1_ASAP7_75t_L g851 ( 
.A1(n_796),
.A2(n_171),
.B(n_173),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_769),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_771),
.B(n_174),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_786),
.B(n_175),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_781),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_805),
.B(n_782),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_836),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_845),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_809),
.B(n_769),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_813),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_816),
.B(n_784),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_818),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_813),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_832),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_815),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_828),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_825),
.B(n_764),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_845),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_809),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_832),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_823),
.B(n_800),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_815),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_804),
.B(n_800),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_817),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_817),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_810),
.A2(n_788),
.B(n_758),
.Y(n_876)
);

AO21x2_ASAP7_75t_L g877 ( 
.A1(n_814),
.A2(n_783),
.B(n_746),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_808),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_807),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_808),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_844),
.B(n_794),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_805),
.B(n_756),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_834),
.B(n_794),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_826),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_812),
.B(n_778),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_821),
.B(n_177),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_839),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_824),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_862),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_878),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_862),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_862),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_860),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_858),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_860),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_883),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_858),
.B(n_889),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_889),
.B(n_888),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_889),
.B(n_827),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_863),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_866),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_857),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_883),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_868),
.B(n_830),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_868),
.B(n_821),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_888),
.B(n_885),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_881),
.B(n_844),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_863),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_869),
.B(n_880),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_883),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_865),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_880),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_908),
.B(n_873),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_897),
.A2(n_835),
.B1(n_856),
.B2(n_904),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_901),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_901),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_902),
.B(n_910),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_905),
.B(n_859),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_901),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_890),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_905),
.B(n_859),
.Y(n_922)
);

NOR3xp33_ASAP7_75t_L g923 ( 
.A(n_903),
.B(n_867),
.C(n_819),
.Y(n_923)
);

AOI211xp5_ASAP7_75t_SL g924 ( 
.A1(n_891),
.A2(n_884),
.B(n_871),
.C(n_886),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_894),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_894),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_903),
.B(n_884),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_896),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_896),
.B(n_833),
.C(n_855),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_897),
.B(n_883),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_907),
.B(n_873),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_930),
.B(n_897),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_923),
.B(n_914),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_930),
.B(n_904),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_927),
.B(n_907),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_916),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_925),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_916),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_925),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_926),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_928),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_917),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_919),
.B(n_904),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_920),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_918),
.B(n_911),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_937),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_932),
.B(n_922),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_937),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_940),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_934),
.B(n_924),
.Y(n_950)
);

AOI211xp5_ASAP7_75t_SL g951 ( 
.A1(n_945),
.A2(n_915),
.B(n_853),
.C(n_887),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_933),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_952),
.B(n_935),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_953),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_953),
.B(n_941),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_950),
.B(n_833),
.Y(n_957)
);

NOR2xp67_ASAP7_75t_L g958 ( 
.A(n_950),
.B(n_945),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_951),
.B(n_943),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_947),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_960),
.B(n_946),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_957),
.B(n_756),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_956),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_955),
.B(n_948),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_949),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_954),
.B(n_947),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_958),
.B(n_939),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_960),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_960),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_960),
.B(n_929),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_958),
.B(n_843),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_942),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_964),
.B(n_755),
.Y(n_973)
);

AOI32xp33_ASAP7_75t_L g974 ( 
.A1(n_970),
.A2(n_911),
.A3(n_853),
.B1(n_886),
.B2(n_895),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_969),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_961),
.Y(n_976)
);

NAND3x2_ASAP7_75t_L g977 ( 
.A(n_965),
.B(n_861),
.C(n_929),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_967),
.B(n_931),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_966),
.A2(n_911),
.B1(n_846),
.B2(n_895),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_973),
.A2(n_971),
.B1(n_962),
.B2(n_963),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_977),
.A2(n_962),
.B1(n_856),
.B2(n_877),
.Y(n_981)
);

AOI21xp33_ASAP7_75t_L g982 ( 
.A1(n_976),
.A2(n_944),
.B(n_938),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_974),
.A2(n_843),
.B(n_846),
.C(n_944),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_972),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_975),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

OAI31xp33_ASAP7_75t_SL g987 ( 
.A1(n_984),
.A2(n_979),
.A3(n_831),
.B(n_775),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_980),
.A2(n_938),
.B1(n_936),
.B2(n_917),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_986),
.B(n_831),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_985),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_983),
.B(n_936),
.Y(n_991)
);

INVxp33_ASAP7_75t_SL g992 ( 
.A(n_989),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_990),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_988),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_987),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_991),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_990),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_981),
.B(n_982),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_996),
.B(n_831),
.C(n_776),
.Y(n_999)
);

OAI211xp5_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_806),
.B(n_803),
.C(n_855),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_993),
.B(n_806),
.C(n_803),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_992),
.A2(n_887),
.B(n_854),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_997),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_1003),
.B(n_992),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_998),
.Y(n_1005)
);

AOI211xp5_ASAP7_75t_L g1006 ( 
.A1(n_1000),
.A2(n_887),
.B(n_805),
.C(n_861),
.Y(n_1006)
);

AOI211xp5_ASAP7_75t_L g1007 ( 
.A1(n_1001),
.A2(n_887),
.B(n_805),
.C(n_838),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1002),
.B(n_921),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_1004),
.A2(n_999),
.B1(n_883),
.B2(n_829),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1005),
.A2(n_854),
.B1(n_906),
.B2(n_921),
.Y(n_1010)
);

AOI221xp5_ASAP7_75t_L g1011 ( 
.A1(n_1006),
.A2(n_849),
.B1(n_913),
.B2(n_852),
.C(n_920),
.Y(n_1011)
);

OAI211xp5_ASAP7_75t_SL g1012 ( 
.A1(n_1008),
.A2(n_820),
.B(n_829),
.C(n_850),
.Y(n_1012)
);

AOI211xp5_ASAP7_75t_L g1013 ( 
.A1(n_1007),
.A2(n_805),
.B(n_851),
.C(n_906),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_1005),
.B(n_848),
.C(n_854),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_1004),
.A2(n_854),
.B1(n_820),
.B2(n_829),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_1004),
.A2(n_820),
.B1(n_848),
.B2(n_898),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_SL g1017 ( 
.A(n_1012),
.B(n_1011),
.C(n_1014),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_1009),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1015),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_1016),
.Y(n_1020)
);

AOI221xp5_ASAP7_75t_L g1021 ( 
.A1(n_1013),
.A2(n_849),
.B1(n_909),
.B2(n_912),
.C(n_893),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_900),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_1015),
.B(n_840),
.Y(n_1023)
);

NOR2x1_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_849),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1009),
.A2(n_899),
.B1(n_910),
.B2(n_847),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_1023),
.B(n_899),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1022),
.Y(n_1027)
);

XNOR2x1_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_178),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_SL g1029 ( 
.A(n_1019),
.B(n_1020),
.C(n_1017),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1024),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1021),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_1018),
.Y(n_1033)
);

NOR2x1_ASAP7_75t_L g1034 ( 
.A(n_1019),
.B(n_912),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_1018),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_1019),
.B(n_840),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1018),
.B(n_890),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1036),
.Y(n_1038)
);

OAI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_1035),
.A2(n_856),
.B1(n_909),
.B2(n_893),
.C(n_892),
.Y(n_1039)
);

AOI221xp5_ASAP7_75t_L g1040 ( 
.A1(n_1029),
.A2(n_892),
.B1(n_900),
.B2(n_890),
.C(n_879),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1033),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_1028),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1034),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1037),
.A2(n_851),
.B(n_876),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1031),
.A2(n_847),
.B1(n_877),
.B2(n_781),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1043),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1041),
.A2(n_1027),
.B1(n_1032),
.B2(n_1030),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_1038),
.A2(n_1026),
.B1(n_839),
.B2(n_898),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1042),
.A2(n_842),
.B1(n_841),
.B2(n_877),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_SL g1050 ( 
.A1(n_1039),
.A2(n_856),
.B1(n_811),
.B2(n_822),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1040),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_1046),
.A2(n_1047),
.B1(n_1051),
.B2(n_1048),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1050),
.A2(n_1045),
.B1(n_1044),
.B2(n_856),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_1049),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1052),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1055),
.Y(n_1056)
);

AO22x2_ASAP7_75t_L g1057 ( 
.A1(n_1056),
.A2(n_1053),
.B1(n_1054),
.B2(n_842),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1056),
.A2(n_879),
.B(n_841),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1057),
.A2(n_870),
.B1(n_864),
.B2(n_822),
.Y(n_1059)
);

NAND4xp25_ASAP7_75t_L g1060 ( 
.A(n_1058),
.B(n_870),
.C(n_864),
.D(n_824),
.Y(n_1060)
);

AOI22x1_ASAP7_75t_L g1061 ( 
.A1(n_1057),
.A2(n_811),
.B1(n_870),
.B2(n_864),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_870),
.C(n_864),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1061),
.B(n_837),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1060),
.B(n_837),
.Y(n_1064)
);

AO21x2_ASAP7_75t_L g1065 ( 
.A1(n_1063),
.A2(n_876),
.B(n_874),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1062),
.A2(n_872),
.B(n_875),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_1064),
.B1(n_874),
.B2(n_875),
.C(n_865),
.Y(n_1067)
);

AOI211xp5_ASAP7_75t_L g1068 ( 
.A1(n_1067),
.A2(n_1066),
.B(n_872),
.C(n_882),
.Y(n_1068)
);


endmodule