module fake_ariane_643_n_1411 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1411);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1411;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_1063;
wire n_537;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_38),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_77),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_249),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_66),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_261),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_96),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_142),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_109),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_12),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_164),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_14),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_262),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_19),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_299),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_42),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_337),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_318),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_224),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_103),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_185),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_296),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_300),
.Y(n_366)
);

BUFx2_ASAP7_75t_SL g367 ( 
.A(n_174),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_64),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_254),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_43),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_313),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_336),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_248),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

BUFx2_ASAP7_75t_R g375 ( 
.A(n_331),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_306),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_288),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_43),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_312),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_259),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_209),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_82),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_214),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_202),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_12),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_135),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_90),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_141),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_218),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_200),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_105),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_36),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_154),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_228),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_294),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_89),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_271),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_231),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_32),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_152),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_80),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_307),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_60),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_35),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_268),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_150),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_58),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_277),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_315),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_9),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_6),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_92),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_204),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_65),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_49),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_289),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_258),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_134),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_6),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_206),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_229),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_107),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_130),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_78),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_263),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_175),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_243),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_37),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_309),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_280),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_301),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_68),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_217),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_88),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_76),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_168),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_180),
.B(n_100),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_129),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_113),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_111),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_334),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_155),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_58),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_255),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_241),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_32),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_138),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_115),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_324),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_215),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_276),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_335),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_128),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_310),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_252),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_0),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_56),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_67),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_44),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_220),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_20),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_193),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_163),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_10),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_9),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_240),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_226),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_339),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_298),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_21),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_279),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_3),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_44),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_34),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_110),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_94),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_160),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_219),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_338),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_287),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_316),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_208),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_292),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_146),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_330),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_327),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_33),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_17),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_30),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_95),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_156),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_101),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_8),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_137),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_56),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_314),
.Y(n_499)
);

BUFx10_ASAP7_75t_L g500 ( 
.A(n_212),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_171),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_176),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_37),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_13),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_178),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_72),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_30),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_247),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_60),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_328),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_321),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_260),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_293),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_232),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_151),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_7),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_184),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_131),
.Y(n_518)
);

BUFx8_ASAP7_75t_SL g519 ( 
.A(n_281),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_183),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_283),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_140),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_305),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_234),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_274),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_233),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_238),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_75),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_179),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_221),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_99),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_322),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_282),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_326),
.Y(n_534)
);

INVx5_ASAP7_75t_L g535 ( 
.A(n_348),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_398),
.B(n_0),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_348),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_1),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_348),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_348),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_360),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_1),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_370),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_464),
.B(n_2),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_360),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_415),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_407),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_360),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_501),
.B(n_446),
.Y(n_555)
);

BUFx12f_ASAP7_75t_L g556 ( 
.A(n_474),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_360),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_476),
.B(n_2),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_421),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_3),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_509),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_404),
.B(n_4),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_404),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_509),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_509),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_358),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_349),
.B(n_4),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_474),
.B(n_480),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_405),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_371),
.B(n_5),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_368),
.B(n_5),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_405),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_440),
.B(n_63),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_399),
.B(n_7),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_405),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_480),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_473),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_369),
.B(n_8),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

BUFx12f_ASAP7_75t_L g582 ( 
.A(n_500),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_500),
.B(n_10),
.Y(n_584)
);

NOR2x1_ASAP7_75t_L g585 ( 
.A(n_400),
.B(n_69),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_471),
.B(n_11),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_11),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_430),
.B(n_13),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_379),
.B(n_14),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_352),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_381),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_463),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_392),
.B(n_15),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_383),
.B(n_15),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_463),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_354),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_384),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_70),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_387),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_402),
.B(n_16),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_512),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_481),
.B(n_16),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_357),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_533),
.B(n_17),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_461),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_359),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_394),
.B(n_18),
.Y(n_612)
);

CKINVDCx6p67_ASAP7_75t_R g613 ( 
.A(n_372),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_378),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_469),
.B(n_531),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_512),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_416),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_417),
.B(n_18),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_344),
.B(n_19),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_418),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_385),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_419),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_374),
.B(n_466),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_423),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_403),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_410),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_411),
.B(n_449),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_343),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_425),
.Y(n_629)
);

BUFx8_ASAP7_75t_SL g630 ( 
.A(n_342),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_534),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_426),
.B(n_428),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_431),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_460),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_436),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_539),
.A2(n_467),
.B1(n_468),
.B2(n_462),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_567),
.B(n_375),
.Y(n_638)
);

OAI22xp33_ASAP7_75t_L g639 ( 
.A1(n_596),
.A2(n_503),
.B1(n_376),
.B2(n_408),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_569),
.B(n_475),
.Y(n_640)
);

INVx8_ASAP7_75t_L g641 ( 
.A(n_549),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_377),
.B1(n_455),
.B2(n_445),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_551),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_578),
.B(n_477),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_543),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_578),
.B(n_490),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_578),
.B(n_615),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_545),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_548),
.B(n_491),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_628),
.B(n_555),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_550),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_552),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

AOI22x1_ASAP7_75t_SL g654 ( 
.A1(n_538),
.A2(n_492),
.B1(n_516),
.B2(n_498),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_627),
.B(n_361),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_536),
.A2(n_581),
.B1(n_583),
.B2(n_564),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_626),
.B(n_437),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_556),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_561),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_L g661 ( 
.A1(n_536),
.A2(n_514),
.B1(n_521),
.B2(n_489),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_607),
.A2(n_523),
.B1(n_517),
.B2(n_458),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_609),
.A2(n_517),
.B1(n_482),
.B2(n_439),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_SL g664 ( 
.A1(n_539),
.A2(n_482),
.B1(n_447),
.B2(n_451),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_559),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_560),
.A2(n_443),
.B1(n_454),
.B2(n_452),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_626),
.B(n_592),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_581),
.B(n_470),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_634),
.B(n_367),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_SL g671 ( 
.A1(n_564),
.A2(n_532),
.B1(n_478),
.B2(n_479),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_584),
.A2(n_483),
.B1(n_485),
.B2(n_472),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_603),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_615),
.B(n_499),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_565),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_619),
.A2(n_511),
.B1(n_522),
.B2(n_505),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_566),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_544),
.A2(n_528),
.B1(n_529),
.B2(n_524),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_571),
.A2(n_502),
.B1(n_520),
.B2(n_487),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_546),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_540),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_SL g682 ( 
.A1(n_544),
.A2(n_346),
.B1(n_347),
.B2(n_345),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_608),
.A2(n_351),
.B1(n_353),
.B2(n_350),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_608),
.B(n_355),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_621),
.B(n_356),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_540),
.Y(n_686)
);

OA22x2_ASAP7_75t_L g687 ( 
.A1(n_591),
.A2(n_363),
.B1(n_364),
.B2(n_362),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_628),
.B(n_365),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_621),
.A2(n_373),
.B1(n_380),
.B2(n_366),
.Y(n_689)
);

OAI22xp33_ASAP7_75t_R g690 ( 
.A1(n_586),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_625),
.A2(n_386),
.B1(n_388),
.B2(n_382),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

OR2x6_ASAP7_75t_L g693 ( 
.A(n_582),
.B(n_519),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_625),
.A2(n_390),
.B1(n_393),
.B2(n_391),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_395),
.B1(n_397),
.B2(n_396),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_611),
.B(n_401),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_558),
.A2(n_406),
.B1(n_412),
.B2(n_409),
.Y(n_697)
);

AO22x2_ASAP7_75t_L g698 ( 
.A1(n_558),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_SL g699 ( 
.A1(n_632),
.A2(n_414),
.B1(n_420),
.B2(n_413),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_576),
.B(n_424),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_632),
.A2(n_429),
.B1(n_432),
.B2(n_427),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_L g702 ( 
.A1(n_613),
.A2(n_435),
.B1(n_438),
.B2(n_433),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_546),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_611),
.B(n_441),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_614),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_563),
.A2(n_530),
.B1(n_527),
.B2(n_526),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_599),
.A2(n_518),
.B1(n_515),
.B2(n_513),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_568),
.A2(n_510),
.B1(n_508),
.B2(n_506),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_576),
.A2(n_497),
.B1(n_495),
.B2(n_494),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_588),
.A2(n_493),
.B1(n_488),
.B2(n_486),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_568),
.A2(n_484),
.B1(n_465),
.B2(n_457),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_572),
.A2(n_456),
.B1(n_453),
.B2(n_450),
.Y(n_713)
);

AO22x2_ASAP7_75t_L g714 ( 
.A1(n_572),
.A2(n_590),
.B1(n_597),
.B2(n_580),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_610),
.A2(n_448),
.B1(n_442),
.B2(n_434),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_541),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_SL g717 ( 
.A1(n_591),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_610),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_541),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_574),
.A2(n_434),
.B1(n_389),
.B2(n_28),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_636),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_651),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_666),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_703),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_658),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_668),
.B(n_624),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_714),
.A2(n_623),
.B(n_590),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_645),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_642),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_652),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_650),
.B(n_593),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_674),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_669),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_660),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_696),
.B(n_600),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_655),
.B(n_629),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_640),
.B(n_602),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_680),
.Y(n_740)
);

XOR2xp5_ASAP7_75t_L g741 ( 
.A(n_638),
.B(n_630),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_714),
.B(n_574),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_665),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_647),
.Y(n_744)
);

XOR2xp5_ASAP7_75t_L g745 ( 
.A(n_639),
.B(n_585),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_675),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_677),
.Y(n_747)
);

INVxp67_ASAP7_75t_SL g748 ( 
.A(n_657),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_657),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_681),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_644),
.B(n_575),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_646),
.B(n_617),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_641),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_716),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_656),
.B(n_580),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_719),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_680),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_649),
.B(n_620),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_653),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_653),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_673),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_673),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_705),
.B(n_620),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_670),
.B(n_620),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

NAND2x1_ASAP7_75t_L g768 ( 
.A(n_720),
.B(n_574),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_686),
.Y(n_769)
);

XOR2xp5_ASAP7_75t_L g770 ( 
.A(n_708),
.B(n_597),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_684),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_700),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_685),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_676),
.Y(n_774)
);

NOR2x1p5_ASAP7_75t_L g775 ( 
.A(n_641),
.B(n_612),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_678),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_679),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_679),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_688),
.B(n_622),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_718),
.B(n_622),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_695),
.B(n_622),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_659),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_706),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_671),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_687),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_672),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_664),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_710),
.B(n_631),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_663),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_667),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_698),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_698),
.Y(n_792)
);

XNOR2x2_ASAP7_75t_L g793 ( 
.A(n_662),
.B(n_612),
.Y(n_793)
);

XOR2x2_ASAP7_75t_L g794 ( 
.A(n_637),
.B(n_618),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_704),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_707),
.B(n_631),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_704),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_711),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_715),
.B(n_618),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_683),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_689),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_691),
.B(n_631),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_713),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_699),
.Y(n_806)
);

INVxp33_ASAP7_75t_L g807 ( 
.A(n_717),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_701),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_702),
.B(n_586),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_712),
.A2(n_587),
.B(n_547),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_799),
.B(n_690),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_733),
.B(n_709),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_735),
.B(n_693),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_727),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_735),
.B(n_693),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_727),
.B(n_633),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_795),
.B(n_574),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_749),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_809),
.A2(n_733),
.B1(n_770),
.B2(n_800),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_754),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_734),
.B(n_587),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_734),
.B(n_682),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_633),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_738),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_782),
.B(n_633),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_783),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_737),
.B(n_635),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_737),
.B(n_635),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_765),
.B(n_744),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_758),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_739),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_769),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_782),
.B(n_635),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_783),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_736),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_765),
.B(n_744),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_740),
.B(n_731),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_774),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_783),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_772),
.B(n_690),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_748),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_772),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_768),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_771),
.B(n_773),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_779),
.B(n_661),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_810),
.A2(n_601),
.B(n_589),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_748),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_779),
.B(n_547),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_730),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_722),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_721),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_SL g852 ( 
.A(n_756),
.B(n_601),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_766),
.B(n_589),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_750),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_732),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_766),
.B(n_601),
.Y(n_856)
);

INVxp33_ASAP7_75t_L g857 ( 
.A(n_796),
.Y(n_857)
);

AND2x2_ASAP7_75t_SL g858 ( 
.A(n_797),
.B(n_601),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_801),
.B(n_654),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_760),
.B(n_598),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_772),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_781),
.B(n_598),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_723),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_780),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_791),
.B(n_26),
.Y(n_865)
);

AND2x6_ASAP7_75t_L g866 ( 
.A(n_742),
.B(n_541),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_767),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_743),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_753),
.B(n_27),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_753),
.B(n_28),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_803),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_803),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_802),
.A2(n_804),
.B1(n_798),
.B2(n_805),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_724),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_792),
.B(n_29),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_781),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_776),
.B(n_29),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_752),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_789),
.B(n_31),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_788),
.B(n_598),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_725),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_788),
.B(n_729),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_777),
.B(n_31),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_729),
.B(n_542),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_752),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_790),
.B(n_33),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_786),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_787),
.B(n_542),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_746),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_806),
.B(n_654),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_778),
.B(n_34),
.Y(n_892)
);

AND2x6_ASAP7_75t_L g893 ( 
.A(n_742),
.B(n_542),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_747),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_784),
.B(n_557),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_759),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_761),
.B(n_71),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_810),
.A2(n_434),
.B(n_389),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_793),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_808),
.B(n_557),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_SL g901 ( 
.A(n_762),
.B(n_535),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_785),
.B(n_35),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_763),
.B(n_36),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_755),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_775),
.B(n_38),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_818),
.Y(n_907)
);

AND2x6_ASAP7_75t_L g908 ( 
.A(n_817),
.B(n_764),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_818),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_849),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_861),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_861),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_861),
.B(n_757),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_820),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_861),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_835),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_842),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_849),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_857),
.B(n_876),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_871),
.B(n_794),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_825),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_842),
.B(n_872),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_835),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_831),
.B(n_807),
.Y(n_924)
);

CKINVDCx6p67_ASAP7_75t_R g925 ( 
.A(n_840),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_843),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_831),
.B(n_745),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_883),
.B(n_741),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_837),
.B(n_39),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_812),
.B(n_389),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_820),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_855),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_855),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_868),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_868),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_814),
.B(n_39),
.Y(n_937)
);

OR2x6_ASAP7_75t_L g938 ( 
.A(n_883),
.B(n_557),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_826),
.B(n_40),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_889),
.Y(n_940)
);

BUFx4f_ASAP7_75t_L g941 ( 
.A(n_895),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_883),
.B(n_570),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_876),
.B(n_389),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_899),
.B(n_389),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_843),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_841),
.B(n_389),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_857),
.B(n_40),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_843),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_889),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_878),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_814),
.B(n_41),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_826),
.B(n_41),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_824),
.B(n_42),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_878),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_894),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_824),
.B(n_45),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_894),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_834),
.Y(n_958)
);

BUFx8_ASAP7_75t_L g959 ( 
.A(n_813),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_847),
.B(n_434),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_903),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_834),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_850),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_850),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_833),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_892),
.B(n_570),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_888),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_811),
.B(n_819),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_882),
.B(n_434),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_839),
.B(n_45),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_863),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_903),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_899),
.B(n_434),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_905),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_900),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_811),
.B(n_46),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_823),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_974),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_948),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_908),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_922),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_948),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_922),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_948),
.Y(n_984)
);

INVx6_ASAP7_75t_L g985 ( 
.A(n_963),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_931),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_948),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_932),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_926),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_917),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_920),
.A2(n_859),
.B1(n_840),
.B2(n_895),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_968),
.B(n_865),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_914),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_926),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_963),
.B(n_829),
.Y(n_995)
);

INVx8_ASAP7_75t_L g996 ( 
.A(n_908),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_917),
.Y(n_997)
);

OR2x6_ASAP7_75t_L g998 ( 
.A(n_938),
.B(n_892),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_959),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_959),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_974),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_910),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_919),
.B(n_887),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_932),
.Y(n_1004)
);

BUFx2_ASAP7_75t_R g1005 ( 
.A(n_927),
.Y(n_1005)
);

AO22x1_ASAP7_75t_L g1006 ( 
.A1(n_920),
.A2(n_859),
.B1(n_815),
.B2(n_890),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_908),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_918),
.Y(n_1008)
);

BUFx12f_ASAP7_75t_L g1009 ( 
.A(n_928),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_958),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_924),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_911),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_925),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_976),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_961),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_937),
.Y(n_1016)
);

CKINVDCx11_ASAP7_75t_R g1017 ( 
.A(n_928),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_945),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_961),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_938),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_938),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_941),
.B(n_865),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_911),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_942),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_958),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_908),
.B(n_839),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_915),
.B(n_945),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_933),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_962),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_919),
.B(n_840),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_928),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_951),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_941),
.A2(n_885),
.B1(n_887),
.B2(n_845),
.Y(n_1033)
);

BUFx4_ASAP7_75t_SL g1034 ( 
.A(n_942),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_965),
.B(n_838),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_962),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_935),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_911),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_963),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_940),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1030),
.A2(n_947),
.B1(n_890),
.B2(n_908),
.Y(n_1041)
);

INVx6_ASAP7_75t_L g1042 ( 
.A(n_986),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1003),
.B(n_967),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_995),
.A2(n_898),
.B(n_943),
.Y(n_1044)
);

INVx8_ASAP7_75t_L g1045 ( 
.A(n_996),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_SL g1046 ( 
.A1(n_1014),
.A2(n_973),
.B1(n_944),
.B2(n_879),
.Y(n_1046)
);

CKINVDCx6p67_ASAP7_75t_R g1047 ( 
.A(n_986),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_978),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_980),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_993),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_1017),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_992),
.A2(n_947),
.B1(n_973),
.B2(n_944),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_992),
.B(n_975),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1001),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_991),
.B(n_929),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1002),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1008),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1011),
.A2(n_877),
.B1(n_886),
.B2(n_921),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_998),
.A2(n_902),
.B1(n_966),
.B2(n_942),
.Y(n_1059)
);

CKINVDCx11_ASAP7_75t_R g1060 ( 
.A(n_999),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_1000),
.Y(n_1061)
);

BUFx10_ASAP7_75t_L g1062 ( 
.A(n_1013),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1028),
.B(n_838),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_1013),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_981),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1009),
.A2(n_864),
.B1(n_874),
.B2(n_863),
.Y(n_1066)
);

CKINVDCx11_ASAP7_75t_R g1067 ( 
.A(n_1017),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1037),
.Y(n_1068)
);

CKINVDCx14_ASAP7_75t_R g1069 ( 
.A(n_1031),
.Y(n_1069)
);

INVx6_ASAP7_75t_L g1070 ( 
.A(n_1009),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1016),
.A2(n_874),
.B1(n_881),
.B2(n_844),
.Y(n_1071)
);

OAI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1032),
.A2(n_966),
.B1(n_822),
.B2(n_881),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_SL g1073 ( 
.A1(n_1031),
.A2(n_902),
.B1(n_892),
.B2(n_875),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_981),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_988),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_980),
.Y(n_1076)
);

INVx3_ASAP7_75t_SL g1077 ( 
.A(n_985),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_980),
.Y(n_1078)
);

BUFx2_ASAP7_75t_SL g1079 ( 
.A(n_983),
.Y(n_1079)
);

OAI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_998),
.A2(n_966),
.B1(n_852),
.B2(n_965),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1034),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_988),
.Y(n_1082)
);

BUFx4f_ASAP7_75t_SL g1083 ( 
.A(n_997),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1033),
.A2(n_972),
.B1(n_936),
.B2(n_977),
.Y(n_1084)
);

NAND2x1p5_ASAP7_75t_L g1085 ( 
.A(n_1007),
.B(n_915),
.Y(n_1085)
);

CKINVDCx11_ASAP7_75t_R g1086 ( 
.A(n_997),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_983),
.Y(n_1087)
);

INVx6_ASAP7_75t_L g1088 ( 
.A(n_1021),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_1010),
.Y(n_1089)
);

INVx6_ASAP7_75t_L g1090 ( 
.A(n_1021),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1010),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1040),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1022),
.A2(n_955),
.B1(n_957),
.B2(n_949),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_1022),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1035),
.A2(n_909),
.B1(n_907),
.B2(n_865),
.Y(n_1095)
);

CKINVDCx6p67_ASAP7_75t_R g1096 ( 
.A(n_1025),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1006),
.A2(n_875),
.B1(n_858),
.B2(n_906),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_1083),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1044),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1041),
.A2(n_906),
.B(n_870),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1055),
.A2(n_875),
.B1(n_998),
.B2(n_816),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1052),
.A2(n_998),
.B1(n_939),
.B2(n_970),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1056),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1043),
.B(n_873),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1045),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1073),
.A2(n_1097),
.B1(n_1046),
.B2(n_1071),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1048),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1069),
.B(n_953),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1058),
.A2(n_916),
.B1(n_923),
.B2(n_963),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1059),
.A2(n_956),
.B1(n_971),
.B2(n_964),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1043),
.A2(n_939),
.B1(n_970),
.B2(n_952),
.Y(n_1111)
);

AOI222xp33_ASAP7_75t_L g1112 ( 
.A1(n_1053),
.A2(n_869),
.B1(n_906),
.B2(n_904),
.C1(n_858),
.C2(n_930),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_1067),
.Y(n_1113)
);

OAI21xp33_ASAP7_75t_L g1114 ( 
.A1(n_1063),
.A2(n_821),
.B(n_943),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1059),
.A2(n_952),
.B(n_846),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_SL g1116 ( 
.A(n_1051),
.B(n_897),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1072),
.A2(n_971),
.B1(n_964),
.B2(n_1004),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1057),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1080),
.A2(n_930),
.B(n_897),
.C(n_827),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1053),
.A2(n_1007),
.B1(n_996),
.B2(n_1005),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1086),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1095),
.A2(n_964),
.B1(n_971),
.B2(n_996),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_1077),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1094),
.A2(n_971),
.B1(n_964),
.B2(n_1004),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1094),
.B(n_1021),
.Y(n_1125)
);

OAI222xp33_ASAP7_75t_L g1126 ( 
.A1(n_1063),
.A2(n_1015),
.B1(n_1019),
.B2(n_1007),
.C1(n_1024),
.C2(n_836),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1068),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1066),
.A2(n_1015),
.B1(n_1019),
.B2(n_854),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1084),
.A2(n_854),
.B1(n_996),
.B2(n_851),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_1089),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1070),
.A2(n_851),
.B1(n_891),
.B2(n_1026),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1050),
.A2(n_896),
.B1(n_954),
.B2(n_950),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1092),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1091),
.B(n_1025),
.Y(n_1134)
);

INVx4_ASAP7_75t_L g1135 ( 
.A(n_1096),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1070),
.A2(n_891),
.B1(n_1026),
.B2(n_995),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1054),
.Y(n_1137)
);

BUFx4f_ASAP7_75t_SL g1138 ( 
.A(n_1047),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1093),
.A2(n_828),
.B1(n_1026),
.B2(n_1024),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1081),
.A2(n_1007),
.B1(n_1024),
.B2(n_1020),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1081),
.B(n_1065),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1064),
.A2(n_848),
.B(n_946),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1075),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1061),
.A2(n_896),
.B1(n_1007),
.B2(n_990),
.Y(n_1144)
);

CKINVDCx11_ASAP7_75t_R g1145 ( 
.A(n_1060),
.Y(n_1145)
);

AOI211xp5_ASAP7_75t_L g1146 ( 
.A1(n_1074),
.A2(n_901),
.B(n_1036),
.C(n_1029),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1079),
.B(n_1029),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1082),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1087),
.A2(n_1036),
.B1(n_990),
.B2(n_969),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1049),
.A2(n_985),
.B1(n_989),
.B2(n_994),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1045),
.A2(n_817),
.B1(n_860),
.B2(n_830),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1042),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1088),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1062),
.B(n_1039),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1088),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1090),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1090),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1062),
.B(n_1039),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1049),
.B(n_989),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1042),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1106),
.A2(n_1045),
.B1(n_1078),
.B2(n_1076),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1103),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1112),
.A2(n_1078),
.B1(n_1076),
.B2(n_934),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1100),
.A2(n_985),
.B1(n_1018),
.B2(n_989),
.Y(n_1164)
);

OAI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1115),
.A2(n_960),
.B1(n_946),
.B2(n_1044),
.C(n_853),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1101),
.A2(n_934),
.B1(n_969),
.B2(n_817),
.Y(n_1166)
);

AOI222xp33_ASAP7_75t_L g1167 ( 
.A1(n_1104),
.A2(n_1101),
.B1(n_1111),
.B2(n_1102),
.C1(n_1116),
.C2(n_1114),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1120),
.A2(n_830),
.B1(n_832),
.B2(n_893),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1130),
.B(n_46),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1120),
.A2(n_832),
.B1(n_893),
.B2(n_866),
.Y(n_1170)
);

CKINVDCx14_ASAP7_75t_R g1171 ( 
.A(n_1145),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1109),
.A2(n_893),
.B1(n_866),
.B2(n_880),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1139),
.A2(n_893),
.B1(n_866),
.B2(n_862),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1139),
.A2(n_893),
.B1(n_866),
.B2(n_994),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1110),
.A2(n_994),
.B1(n_1018),
.B2(n_982),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1110),
.A2(n_1018),
.B1(n_982),
.B2(n_984),
.Y(n_1176)
);

OAI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1121),
.A2(n_979),
.B1(n_987),
.B2(n_911),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1149),
.A2(n_982),
.B1(n_984),
.B2(n_979),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1129),
.A2(n_866),
.B1(n_960),
.B2(n_867),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1142),
.A2(n_867),
.B1(n_912),
.B2(n_984),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1149),
.A2(n_912),
.B1(n_1027),
.B2(n_1038),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1136),
.A2(n_987),
.B1(n_979),
.B2(n_1023),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1132),
.B(n_1038),
.C(n_1023),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1125),
.A2(n_912),
.B1(n_856),
.B2(n_1027),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1118),
.B(n_1127),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_912),
.B1(n_884),
.B2(n_913),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1146),
.B(n_1012),
.C(n_987),
.Y(n_1187)
);

OAI211xp5_ASAP7_75t_SL g1188 ( 
.A1(n_1133),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1188)
);

OAI211xp5_ASAP7_75t_L g1189 ( 
.A1(n_1099),
.A2(n_898),
.B(n_1012),
.C(n_987),
.Y(n_1189)
);

OAI222xp33_ASAP7_75t_L g1190 ( 
.A1(n_1117),
.A2(n_1085),
.B1(n_913),
.B2(n_987),
.C1(n_979),
.C2(n_52),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1121),
.A2(n_979),
.B1(n_1085),
.B2(n_1012),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1131),
.A2(n_1012),
.B1(n_48),
.B2(n_50),
.Y(n_1192)
);

OAI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1147),
.A2(n_616),
.B1(n_605),
.B2(n_595),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1141),
.B(n_47),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1123),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1122),
.A2(n_616),
.B1(n_570),
.B2(n_605),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1107),
.A2(n_616),
.B1(n_605),
.B2(n_595),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1137),
.A2(n_1108),
.B1(n_1122),
.B2(n_1128),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1143),
.A2(n_577),
.B1(n_573),
.B2(n_595),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1148),
.A2(n_573),
.B1(n_577),
.B2(n_594),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1135),
.A2(n_573),
.B1(n_577),
.B2(n_594),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1134),
.B(n_51),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1140),
.A2(n_594),
.B1(n_604),
.B2(n_606),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1140),
.A2(n_606),
.B1(n_604),
.B2(n_554),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1153),
.B(n_53),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1124),
.A2(n_606),
.B1(n_604),
.B2(n_554),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1154),
.B(n_53),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1151),
.A2(n_606),
.B1(n_604),
.B2(n_554),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_SL g1209 ( 
.A1(n_1119),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.C(n_59),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1144),
.A2(n_554),
.B1(n_537),
.B2(n_535),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1155),
.A2(n_537),
.B1(n_535),
.B2(n_57),
.Y(n_1211)
);

OAI211xp5_ASAP7_75t_L g1212 ( 
.A1(n_1099),
.A2(n_54),
.B(n_55),
.C(n_59),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1158),
.B(n_61),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1156),
.A2(n_537),
.B1(n_535),
.B2(n_61),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1157),
.B(n_1159),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1113),
.A2(n_62),
.B1(n_537),
.B2(n_74),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1152),
.A2(n_62),
.B(n_73),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1162),
.B(n_1123),
.Y(n_1218)
);

AND2x2_ASAP7_75t_SL g1219 ( 
.A(n_1216),
.B(n_1135),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1209),
.B(n_1150),
.C(n_1098),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1194),
.B(n_1098),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1215),
.B(n_1160),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1161),
.A2(n_1105),
.B1(n_1138),
.B2(n_1126),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1185),
.B(n_1105),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1167),
.B(n_1105),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1207),
.B(n_1213),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1198),
.B(n_1105),
.Y(n_1227)
);

NAND3xp33_ASAP7_75t_L g1228 ( 
.A(n_1212),
.B(n_1126),
.C(n_1138),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1217),
.B(n_79),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1202),
.B(n_341),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1216),
.B(n_81),
.C(n_83),
.Y(n_1231)
);

OAI221xp5_ASAP7_75t_L g1232 ( 
.A1(n_1161),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1188),
.A2(n_91),
.B1(n_93),
.B2(n_97),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1169),
.B(n_340),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1198),
.B(n_98),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1183),
.B(n_333),
.Y(n_1236)
);

NAND3xp33_ASAP7_75t_L g1237 ( 
.A(n_1195),
.B(n_102),
.C(n_104),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1181),
.B(n_106),
.Y(n_1238)
);

OAI221xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1163),
.A2(n_108),
.B1(n_112),
.B2(n_114),
.C(n_116),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1205),
.B(n_332),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_L g1241 ( 
.A(n_1180),
.B(n_117),
.C(n_118),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_SL g1242 ( 
.A(n_1187),
.B(n_1190),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1171),
.A2(n_119),
.B(n_120),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1211),
.A2(n_121),
.B(n_122),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1163),
.B(n_1178),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1189),
.A2(n_123),
.B(n_124),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1164),
.B(n_1175),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1165),
.B(n_125),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1214),
.A2(n_126),
.B1(n_127),
.B2(n_132),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1191),
.B(n_133),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1176),
.B(n_1177),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1184),
.B(n_329),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1186),
.B(n_136),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1192),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1166),
.B(n_145),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1170),
.A2(n_147),
.B(n_148),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1166),
.B(n_323),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1203),
.A2(n_149),
.B(n_153),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1168),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1182),
.B(n_320),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1204),
.B(n_161),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1173),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1174),
.B(n_167),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1196),
.B(n_169),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1179),
.B(n_170),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1224),
.Y(n_1266)
);

OR2x2_ASAP7_75t_SL g1267 ( 
.A(n_1228),
.B(n_1201),
.Y(n_1267)
);

OAI211xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1218),
.A2(n_1210),
.B(n_1208),
.C(n_1172),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1242),
.A2(n_1193),
.B1(n_1197),
.B2(n_1206),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1222),
.B(n_172),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_L g1271 ( 
.A(n_1246),
.B(n_1197),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_L g1272 ( 
.A(n_1248),
.B(n_1200),
.C(n_1199),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1224),
.B(n_173),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1221),
.B(n_319),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1248),
.B(n_177),
.C(n_181),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1247),
.B(n_182),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1226),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1227),
.Y(n_1278)
);

NAND3xp33_ASAP7_75t_L g1279 ( 
.A(n_1231),
.B(n_186),
.C(n_187),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_L g1280 ( 
.A(n_1233),
.B(n_188),
.C(n_190),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1225),
.B(n_191),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1245),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1251),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1238),
.Y(n_1284)
);

NAND4xp75_ASAP7_75t_L g1285 ( 
.A(n_1219),
.B(n_192),
.C(n_194),
.D(n_195),
.Y(n_1285)
);

OA211x2_ASAP7_75t_L g1286 ( 
.A1(n_1223),
.A2(n_1236),
.B(n_1220),
.C(n_1229),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1235),
.Y(n_1287)
);

OAI211xp5_ASAP7_75t_L g1288 ( 
.A1(n_1243),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_1288)
);

NAND4xp75_ASAP7_75t_L g1289 ( 
.A(n_1219),
.B(n_199),
.C(n_201),
.D(n_205),
.Y(n_1289)
);

OAI211xp5_ASAP7_75t_L g1290 ( 
.A1(n_1244),
.A2(n_207),
.B(n_210),
.C(n_211),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1240),
.B(n_216),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_1223),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1266),
.B(n_1230),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1282),
.B(n_1234),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1278),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1277),
.B(n_1246),
.Y(n_1296)
);

OAI31xp33_ASAP7_75t_L g1297 ( 
.A1(n_1288),
.A2(n_1229),
.A3(n_1239),
.B(n_1256),
.Y(n_1297)
);

XNOR2x2_ASAP7_75t_L g1298 ( 
.A(n_1271),
.B(n_1255),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1283),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1287),
.B(n_1257),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1284),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1276),
.B(n_1233),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1292),
.B(n_1260),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1276),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1237),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1270),
.B(n_1252),
.Y(n_1306)
);

NAND4xp75_ASAP7_75t_SL g1307 ( 
.A(n_1274),
.B(n_1263),
.C(n_1253),
.D(n_1261),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1281),
.B(n_1263),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1279),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1267),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1309),
.Y(n_1311)
);

XOR2x2_ASAP7_75t_L g1312 ( 
.A(n_1298),
.B(n_1285),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1295),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1300),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1304),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1304),
.B(n_1291),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1300),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1299),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1303),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1293),
.Y(n_1320)
);

XOR2x2_ASAP7_75t_L g1321 ( 
.A(n_1298),
.B(n_1289),
.Y(n_1321)
);

OA22x2_ASAP7_75t_L g1322 ( 
.A1(n_1311),
.A2(n_1310),
.B1(n_1309),
.B2(n_1296),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1313),
.Y(n_1323)
);

OA22x2_ASAP7_75t_L g1324 ( 
.A1(n_1311),
.A2(n_1310),
.B1(n_1296),
.B2(n_1308),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1318),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1314),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1316),
.Y(n_1327)
);

OA22x2_ASAP7_75t_L g1328 ( 
.A1(n_1312),
.A2(n_1321),
.B1(n_1319),
.B2(n_1320),
.Y(n_1328)
);

XNOR2xp5_ASAP7_75t_L g1329 ( 
.A(n_1312),
.B(n_1321),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1317),
.A2(n_1286),
.B1(n_1302),
.B2(n_1308),
.Y(n_1330)
);

XOR2x2_ASAP7_75t_L g1331 ( 
.A(n_1315),
.B(n_1307),
.Y(n_1331)
);

AOI22x1_ASAP7_75t_L g1332 ( 
.A1(n_1311),
.A2(n_1302),
.B1(n_1297),
.B2(n_1290),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1313),
.Y(n_1333)
);

OA22x2_ASAP7_75t_L g1334 ( 
.A1(n_1311),
.A2(n_1294),
.B1(n_1306),
.B2(n_1301),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1327),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1329),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1325),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1323),
.Y(n_1338)
);

XOR2x2_ASAP7_75t_L g1339 ( 
.A(n_1329),
.B(n_1305),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1333),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_SL g1341 ( 
.A(n_1326),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1328),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1322),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1338),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1336),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1340),
.Y(n_1346)
);

OAI22x1_ASAP7_75t_L g1347 ( 
.A1(n_1342),
.A2(n_1332),
.B1(n_1330),
.B2(n_1331),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1337),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1341),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1345),
.A2(n_1332),
.B1(n_1335),
.B2(n_1341),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1345),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1349),
.A2(n_1334),
.B1(n_1343),
.B2(n_1324),
.Y(n_1352)
);

NOR2x1_ASAP7_75t_L g1353 ( 
.A(n_1348),
.B(n_1336),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1344),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1347),
.A2(n_1339),
.B1(n_1275),
.B2(n_1280),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1351),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1350),
.B(n_1346),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1353),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1352),
.A2(n_1280),
.B1(n_1279),
.B2(n_1268),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1354),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1355),
.A2(n_1272),
.B1(n_1249),
.B2(n_1254),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1351),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1353),
.B(n_1232),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1358),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1363),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1360),
.Y(n_1366)
);

NOR3xp33_ASAP7_75t_L g1367 ( 
.A(n_1357),
.B(n_1250),
.C(n_1241),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1356),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1359),
.A2(n_1272),
.B1(n_1269),
.B2(n_1258),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1362),
.Y(n_1370)
);

AO22x2_ASAP7_75t_L g1371 ( 
.A1(n_1365),
.A2(n_1361),
.B1(n_1259),
.B2(n_1261),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1364),
.A2(n_1262),
.B1(n_1265),
.B2(n_1264),
.Y(n_1372)
);

AND4x1_ASAP7_75t_L g1373 ( 
.A(n_1367),
.B(n_1262),
.C(n_1264),
.D(n_225),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1366),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1369),
.A2(n_222),
.B1(n_223),
.B2(n_227),
.Y(n_1375)
);

AO22x2_ASAP7_75t_L g1376 ( 
.A1(n_1370),
.A2(n_230),
.B1(n_235),
.B2(n_236),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1374),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1371),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1375),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1373),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1372),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1376),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1376),
.Y(n_1383)
);

NOR2x1_ASAP7_75t_L g1384 ( 
.A(n_1374),
.B(n_1368),
.Y(n_1384)
);

OAI22x1_ASAP7_75t_L g1385 ( 
.A1(n_1380),
.A2(n_1384),
.B1(n_1378),
.B2(n_1381),
.Y(n_1385)
);

OAI22x1_ASAP7_75t_L g1386 ( 
.A1(n_1377),
.A2(n_237),
.B1(n_239),
.B2(n_242),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1382),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1383),
.A2(n_1379),
.B1(n_245),
.B2(n_246),
.Y(n_1388)
);

XOR2x2_ASAP7_75t_L g1389 ( 
.A(n_1379),
.B(n_244),
.Y(n_1389)
);

OAI211xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1384),
.A2(n_250),
.B(n_251),
.C(n_253),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1380),
.A2(n_256),
.B1(n_257),
.B2(n_264),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1384),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1392),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1386),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1389),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1385),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1387),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1397),
.A2(n_1388),
.B1(n_1391),
.B2(n_1390),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1394),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1393),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1396),
.A2(n_273),
.B1(n_275),
.B2(n_278),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1398),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1399),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1401),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1404),
.A2(n_1395),
.B1(n_1402),
.B2(n_1403),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1403),
.A2(n_1400),
.B1(n_285),
.B2(n_286),
.Y(n_1406)
);

AO22x2_ASAP7_75t_L g1407 ( 
.A1(n_1402),
.A2(n_284),
.B1(n_290),
.B2(n_291),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1405),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1407),
.Y(n_1409)
);

AOI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1409),
.A2(n_1406),
.B1(n_1408),
.B2(n_302),
.C(n_303),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1410),
.A2(n_295),
.B1(n_297),
.B2(n_304),
.Y(n_1411)
);


endmodule