module fake_jpeg_28444_n_46 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_2),
.B(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.B(n_19),
.Y(n_27)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_19),
.B1(n_20),
.B2(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_27),
.B1(n_29),
.B2(n_3),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_18),
.C(n_19),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_28),
.C(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_38),
.Y(n_40)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_10),
.C(n_2),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_34),
.C(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_1),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_43),
.B1(n_7),
.B2(n_8),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_42),
.C2(n_38),
.Y(n_46)
);


endmodule