module fake_jpeg_13039_n_466 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_466);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_466;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_17),
.B(n_9),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_61),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_66),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_8),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_86),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_78),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_30),
.B(n_20),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_23),
.B(n_10),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_10),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_90),
.Y(n_123)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_18),
.A2(n_6),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_0),
.Y(n_95)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_95),
.B(n_129),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_96),
.A2(n_143),
.B1(n_109),
.B2(n_97),
.Y(n_180)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_138),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_121),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_62),
.A2(n_39),
.B1(n_43),
.B2(n_42),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_98),
.B1(n_134),
.B2(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_26),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_54),
.B(n_44),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_131),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_147),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_84),
.Y(n_138)
);

CKINVDCx10_ASAP7_75t_R g139 ( 
.A(n_65),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

BUFx4f_ASAP7_75t_SL g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_60),
.B(n_32),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_40),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_25),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_43),
.B1(n_87),
.B2(n_82),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_150),
.A2(n_164),
.B(n_110),
.Y(n_205)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_153),
.Y(n_244)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_156),
.Y(n_247)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_30),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_162),
.A2(n_167),
.B1(n_184),
.B2(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_19),
.B1(n_25),
.B2(n_38),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_102),
.A2(n_43),
.B1(n_88),
.B2(n_70),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_102),
.A2(n_30),
.B1(n_37),
.B2(n_34),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_118),
.B1(n_133),
.B2(n_124),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_96),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_31),
.B1(n_37),
.B2(n_34),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_172),
.B1(n_173),
.B2(n_185),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_38),
.C(n_33),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_176),
.Y(n_207)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_27),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_25),
.B1(n_19),
.B2(n_145),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_182),
.B1(n_192),
.B2(n_196),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_203),
.B1(n_137),
.B2(n_118),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_123),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_104),
.C(n_124),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_187),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_103),
.A2(n_19),
.B1(n_29),
.B2(n_3),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_128),
.A2(n_29),
.B1(n_2),
.B2(n_4),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_128),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_1),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_157),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_117),
.B(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_13),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_29),
.B1(n_6),
.B2(n_11),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_106),
.A2(n_92),
.B(n_135),
.C(n_114),
.Y(n_195)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_137),
.B1(n_119),
.B2(n_112),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_92),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_109),
.A2(n_16),
.B1(n_6),
.B2(n_12),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_197),
.A2(n_200),
.B1(n_185),
.B2(n_160),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_5),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_199),
.A2(n_151),
.B1(n_159),
.B2(n_177),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_143),
.A2(n_5),
.B1(n_12),
.B2(n_13),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_146),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_202),
.Y(n_232)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_116),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_205),
.B(n_214),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_208),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_211),
.B(n_212),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_117),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_213),
.A2(n_239),
.B(n_205),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_200),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_104),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_231),
.C(n_149),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_124),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_225),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_133),
.B1(n_104),
.B2(n_15),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_246),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_164),
.A2(n_133),
.B1(n_14),
.B2(n_16),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_152),
.B(n_13),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_150),
.A2(n_14),
.B1(n_16),
.B2(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_152),
.B(n_14),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_152),
.B(n_154),
.C(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_174),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_158),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_206),
.B(n_234),
.C(n_207),
.D(n_228),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_238),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_158),
.A2(n_181),
.B1(n_168),
.B2(n_172),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_197),
.B1(n_155),
.B2(n_166),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_240),
.A2(n_241),
.B1(n_204),
.B2(n_233),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_189),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_175),
.B(n_199),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_166),
.B(n_179),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_248),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_186),
.A2(n_195),
.B1(n_194),
.B2(n_170),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_171),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_153),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_221),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_201),
.B(n_156),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_149),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_260),
.Y(n_297)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_177),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_256),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_285),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_177),
.B(n_202),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_259),
.A2(n_247),
.B(n_244),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_183),
.C(n_175),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_219),
.B(n_175),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_263),
.A2(n_283),
.B(n_208),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_182),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_266),
.B(n_291),
.Y(n_305)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_182),
.B1(n_199),
.B2(n_227),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_272),
.A2(n_278),
.B1(n_277),
.B2(n_269),
.Y(n_321)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_288),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_243),
.B1(n_224),
.B2(n_226),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_252),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_281),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_206),
.C(n_215),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_225),
.B(n_229),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_204),
.B1(n_241),
.B2(n_236),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_284),
.A2(n_294),
.B1(n_223),
.B2(n_213),
.Y(n_304)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_209),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_232),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_287),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_211),
.A2(n_220),
.B(n_236),
.C(n_213),
.D(n_217),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_242),
.C(n_238),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_260),
.Y(n_325)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_230),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_233),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_238),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_247),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_302),
.A2(n_329),
.B(n_273),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_304),
.A2(n_278),
.B1(n_269),
.B2(n_272),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_230),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_309),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_264),
.B(n_214),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_307),
.B(n_310),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_208),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_279),
.B(n_244),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_311),
.B(n_320),
.Y(n_346)
);

OAI21xp33_ASAP7_75t_SL g332 ( 
.A1(n_312),
.A2(n_255),
.B(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_214),
.Y(n_318)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_289),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_321),
.A2(n_275),
.B1(n_285),
.B2(n_318),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_322),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_270),
.B(n_214),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_323),
.B(n_324),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_293),
.B(n_222),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_319),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_274),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_326),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_290),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_255),
.B(n_283),
.C(n_264),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_252),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_354),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_359),
.B1(n_361),
.B2(n_305),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_297),
.B(n_282),
.C(n_253),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_340),
.C(n_353),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_314),
.A2(n_284),
.B1(n_273),
.B2(n_258),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_337),
.A2(n_349),
.B(n_350),
.Y(n_375)
);

OA22x2_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_273),
.B1(n_271),
.B2(n_267),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_348),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_261),
.C(n_283),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_298),
.Y(n_342)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_347),
.B(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_295),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_314),
.A2(n_258),
.B(n_259),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_350),
.A2(n_329),
.B(n_301),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_352),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_307),
.B1(n_327),
.B2(n_316),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_325),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_327),
.A2(n_295),
.B1(n_320),
.B2(n_306),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_323),
.A2(n_295),
.B1(n_326),
.B2(n_328),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_362),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_309),
.B1(n_331),
.B2(n_302),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_296),
.Y(n_362)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_364),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_300),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_369),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_310),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_334),
.A2(n_305),
.B1(n_324),
.B2(n_322),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_372),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_317),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_339),
.B1(n_341),
.B2(n_356),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_373),
.A2(n_376),
.B1(n_382),
.B2(n_384),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_374),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_385),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_301),
.B1(n_315),
.B2(n_308),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_346),
.B(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_378),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_333),
.B(n_299),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_315),
.B1(n_308),
.B2(n_313),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_348),
.A2(n_299),
.B1(n_313),
.B2(n_333),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_357),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_356),
.B1(n_338),
.B2(n_352),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_340),
.B(n_359),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_343),
.Y(n_387)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_387),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_361),
.Y(n_391)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_349),
.C(n_351),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_401),
.C(n_403),
.Y(n_418)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_355),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_395),
.B(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_407),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_345),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_337),
.C(n_338),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_363),
.C(n_365),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_338),
.C(n_342),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_358),
.C(n_406),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_343),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_383),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_399),
.A2(n_396),
.B(n_374),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_412),
.B(n_413),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_408),
.A2(n_379),
.B(n_375),
.C(n_384),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_404),
.A2(n_379),
.B(n_370),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_402),
.B(n_344),
.Y(n_415)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_405),
.A2(n_380),
.B1(n_344),
.B2(n_376),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_421),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_382),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_417),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_380),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_419),
.B(n_416),
.Y(n_436)
);

INVx11_ASAP7_75t_L g422 ( 
.A(n_392),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_406),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_423),
.B(n_425),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_395),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_430),
.B(n_433),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_401),
.C(n_403),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_434),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_394),
.Y(n_433)
);

A2O1A1O1Ixp25_ASAP7_75t_L g434 ( 
.A1(n_411),
.A2(n_388),
.B(n_413),
.C(n_423),
.D(n_412),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_418),
.B(n_388),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_436),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_425),
.C(n_414),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_417),
.C(n_419),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_421),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_421),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_447),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_415),
.B1(n_410),
.B2(n_409),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_448),
.B1(n_427),
.B2(n_431),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_442),
.B(n_444),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_412),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_412),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_426),
.C(n_434),
.Y(n_453)
);

OAI321xp33_ASAP7_75t_L g447 ( 
.A1(n_431),
.A2(n_409),
.A3(n_410),
.B1(n_412),
.B2(n_420),
.C(n_429),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_440),
.A2(n_432),
.B(n_429),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_449),
.A2(n_443),
.B(n_444),
.Y(n_457)
);

BUFx12_ASAP7_75t_L g451 ( 
.A(n_439),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_445),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_446),
.A2(n_420),
.B(n_426),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_455),
.A2(n_442),
.B(n_453),
.Y(n_458)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_450),
.C(n_451),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_457),
.A2(n_458),
.B(n_455),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_460),
.A2(n_461),
.B(n_459),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_462),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_461),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_463),
.B(n_451),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_454),
.Y(n_466)
);


endmodule