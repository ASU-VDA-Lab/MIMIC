module fake_netlist_1_1364_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NOR2xp33_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
BUFx3_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_5), .B(n_0), .Y(n_6) );
OR2x6_ASAP7_75t_L g7 ( .A(n_3), .B(n_0), .Y(n_7) );
CKINVDCx8_ASAP7_75t_R g8 ( .A(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_7), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_8), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B1(n_4), .B2(n_3), .C(n_5), .Y(n_13) );
AOI211xp5_ASAP7_75t_L g14 ( .A1(n_11), .A2(n_10), .B(n_5), .C(n_2), .Y(n_14) );
NAND4xp25_ASAP7_75t_L g15 ( .A(n_13), .B(n_11), .C(n_1), .D(n_2), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_1), .Y(n_16) );
AOI21xp33_ASAP7_75t_SL g17 ( .A1(n_16), .A2(n_1), .B(n_2), .Y(n_17) );
NAND2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
endmodule