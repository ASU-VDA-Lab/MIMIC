module real_jpeg_4832_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_0),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_57),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_1),
.A2(n_73),
.B1(n_205),
.B2(n_309),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_1),
.A2(n_73),
.B1(n_160),
.B2(n_161),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_1),
.A2(n_73),
.B1(n_328),
.B2(n_393),
.Y(n_392)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_2),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_2),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_3),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_3),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_3),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_3),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_4),
.A2(n_53),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_4),
.A2(n_53),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_4),
.A2(n_53),
.B1(n_202),
.B2(n_377),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_5),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_5),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_5),
.A2(n_279),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_5),
.A2(n_279),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g443 ( 
.A1(n_5),
.A2(n_49),
.B1(n_279),
.B2(n_444),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_48),
.B1(n_57),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_60),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_6),
.A2(n_60),
.B1(n_278),
.B2(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_6),
.A2(n_60),
.B1(n_360),
.B2(n_403),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_46),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_7),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_7),
.A2(n_76),
.B1(n_219),
.B2(n_227),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_7),
.A2(n_76),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_7),
.A2(n_76),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_8),
.Y(n_326)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_9),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_10),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_10),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_10),
.A2(n_166),
.B1(n_201),
.B2(n_205),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_10),
.A2(n_166),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_10),
.A2(n_166),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_13),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_15),
.A2(n_181),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_15),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_15),
.A2(n_185),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_15),
.A2(n_185),
.B1(n_268),
.B2(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_15),
.A2(n_185),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_17),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_17),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_17),
.B(n_175),
.C(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_17),
.B(n_88),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_17),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_17),
.B(n_169),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_17),
.B(n_263),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_18),
.A2(n_93),
.B1(n_160),
.B2(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_18),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_18),
.A2(n_211),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_18),
.A2(n_32),
.B1(n_211),
.B2(n_270),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_18),
.A2(n_39),
.B1(n_40),
.B2(n_211),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_520),
.B(n_523),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_63),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_62),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_54),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_24),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_24),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_25),
.B(n_162),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_25),
.A2(n_55),
.B1(n_395),
.B2(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_25)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_27),
.Y(n_260)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_28),
.Y(n_428)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_30),
.Y(n_390)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_30),
.Y(n_431)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_36),
.A2(n_344),
.B(n_346),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_36),
.B(n_348),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_41),
.Y(n_323)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_49),
.B(n_162),
.Y(n_332)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_54),
.B(n_65),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_55),
.A2(n_61),
.B1(n_69),
.B2(n_74),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_74),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_55),
.A2(n_347),
.B(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_55),
.A2(n_61),
.B1(n_69),
.B2(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_61),
.A2(n_416),
.B(n_446),
.Y(n_456)
);

AO21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_149),
.B(n_519),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_145),
.C(n_146),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_66),
.A2(n_67),
.B1(n_515),
.B2(n_516),
.Y(n_514)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_77),
.C(n_112),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_68),
.B(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_72),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_77),
.A2(n_112),
.B1(n_113),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_77),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_78),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_78),
.A2(n_107),
.B1(n_302),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_78),
.A2(n_107),
.B1(n_387),
.B2(n_392),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_78),
.A2(n_100),
.B1(n_107),
.B2(n_496),
.Y(n_495)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_88),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_80),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_87),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_87),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_87),
.Y(n_354)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

AOI22x1_ASAP7_75t_L g417 ( 
.A1(n_88),
.A2(n_147),
.B1(n_304),
.B2(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_88),
.A2(n_147),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_91),
.Y(n_289)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_93),
.B(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_93),
.Y(n_382)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_94),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_96),
.Y(n_359)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_96),
.Y(n_362)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_102),
.Y(n_269)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_106),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_107),
.B(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_107),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_109),
.Y(n_393)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_112),
.A2(n_113),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_112),
.B(n_491),
.C(n_494),
.Y(n_502)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_130),
.B(n_139),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_159),
.B(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_114),
.A2(n_130),
.B1(n_210),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_114),
.A2(n_163),
.B(n_253),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_114),
.A2(n_130),
.B1(n_356),
.B2(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_115),
.B(n_164),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_115),
.A2(n_169),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_115),
.A2(n_169),
.B1(n_381),
.B2(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_115),
.A2(n_169),
.B1(n_402),
.B2(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_130),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_123),
.B2(n_127),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g288 ( 
.A(n_127),
.Y(n_288)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_130),
.A2(n_210),
.B(n_212),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_130),
.A2(n_212),
.B(n_356),
.Y(n_355)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_133),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_134),
.Y(n_135)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_134),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_134),
.Y(n_378)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_139),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_144),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_145),
.B(n_146),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_147),
.A2(n_259),
.B(n_266),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_147),
.B(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_147),
.A2(n_266),
.B(n_459),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_513),
.B(n_518),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_485),
.B(n_510),
.Y(n_150)
);

OAI311xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_365),
.A3(n_461),
.B1(n_479),
.C1(n_480),
.Y(n_151)
);

AOI21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_315),
.B(n_364),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_293),
.B(n_314),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_247),
.B(n_292),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_215),
.B(n_246),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_178),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_157),
.B(n_178),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_170),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_158),
.A2(n_170),
.B1(n_171),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_162),
.A2(n_189),
.B(n_196),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_162),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_SL g344 ( 
.A1(n_162),
.A2(n_332),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_207),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_208),
.C(n_214),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_189),
.B(n_196),
.Y(n_179)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_182),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_189),
.A2(n_198),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_189),
.A2(n_371),
.B1(n_374),
.B2(n_376),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_189),
.A2(n_198),
.B(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_200),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_190),
.A2(n_276),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_190),
.A2(n_337),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_192),
.Y(n_312)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_195),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_225),
.B(n_234),
.Y(n_224)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_237),
.B(n_245),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_236),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_235),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_235),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_234),
.A2(n_275),
.B(n_282),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_243),
.Y(n_245)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_249),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_273),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_257),
.B2(n_258),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_257),
.C(n_273),
.Y(n_294)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_256),
.Y(n_384)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_286),
.A3(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_272),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_285),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_284),
.Y(n_375)
);

INVx4_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_295),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_300),
.B2(n_313),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_299),
.C(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_306),
.C(n_307),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_316),
.B(n_317),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_341),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_318)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_333),
.B2(n_334),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_321),
.B(n_333),
.Y(n_457)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.A3(n_324),
.B1(n_327),
.B2(n_332),
.Y(n_321)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_329),
.Y(n_328)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_338),
.B(n_340),
.C(n_341),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_351),
.B2(n_363),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_342),
.B(n_352),
.C(n_355),
.Y(n_470)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_353),
.Y(n_459)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_447),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_366),
.A2(n_447),
.B(n_481),
.C(n_484),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_419),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_367),
.B(n_419),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_399),
.C(n_406),
.Y(n_367)
);

FAx1_ASAP7_75t_SL g460 ( 
.A(n_368),
.B(n_399),
.CI(n_406),
.CON(n_460),
.SN(n_460)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_385),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_386),
.C(n_394),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_379),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_370),
.B(n_379),
.Y(n_453)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_380),
.Y(n_409)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_387),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx6_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_392),
.Y(n_426)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_404),
.B2(n_405),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_404),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_404),
.A2(n_405),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_404),
.A2(n_438),
.B(n_441),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_414),
.C(n_417),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_408),
.B(n_410),
.Y(n_469)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_414),
.A2(n_415),
.B1(n_417),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_417),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_420),
.B(n_423),
.C(n_436),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_436),
.B2(n_437),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_432),
.B(n_435),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_433),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_427),
.Y(n_496)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_435),
.B(n_488),
.CI(n_489),
.CON(n_487),
.SN(n_487)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_435),
.B(n_488),
.C(n_489),
.Y(n_509)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_443),
.Y(n_492)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_460),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_460),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_453),
.C(n_454),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_449),
.A2(n_450),
.B1(n_453),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.C(n_458),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_457),
.B(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_458),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_460),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_463),
.A2(n_482),
.B(n_483),
.Y(n_481)
);

NOR2x1_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_471),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_471),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.C(n_470),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_477),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_469),
.B1(n_470),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_470),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_475),
.B(n_476),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_499),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_498),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_498),
.Y(n_511)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_487),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_491),
.B1(n_493),
.B2(n_497),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_490),
.A2(n_491),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_501),
.C(n_505),
.Y(n_517)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_493),
.Y(n_497)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_499),
.A2(n_511),
.B(n_512),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_509),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_509),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_517),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_517),
.Y(n_518)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_521),
.Y(n_524)
);

INVx13_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);


endmodule