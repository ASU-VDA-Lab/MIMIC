module fake_jpeg_8149_n_98 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_16),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_32),
.B(n_26),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_26),
.B(n_39),
.C(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_55),
.B1(n_39),
.B2(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_27),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_64),
.B(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_45),
.A2(n_39),
.B1(n_14),
.B2(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_39),
.B1(n_56),
.B2(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_72),
.B1(n_65),
.B2(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_59),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_58),
.C(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_83),
.C(n_76),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_15),
.B(n_10),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_64),
.B1(n_54),
.B2(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_78),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_85),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_82),
.C(n_79),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_80),
.B(n_10),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_11),
.B(n_15),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_11),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_97),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_91),
.B1(n_92),
.B2(n_82),
.Y(n_97)
);


endmodule