module fake_jpeg_308_n_215 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_215);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g69 ( 
.A(n_15),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_53),
.Y(n_85)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_84),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_52),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_58),
.B1(n_64),
.B2(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_67),
.B1(n_75),
.B2(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_97),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_69),
.B1(n_67),
.B2(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_65),
.B1(n_82),
.B2(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_75),
.C(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_70),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_R g138 ( 
.A(n_105),
.B(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_111),
.A2(n_76),
.B1(n_65),
.B2(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_63),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.C(n_116),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_86),
.B1(n_90),
.B2(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_111),
.B1(n_110),
.B2(n_105),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_138),
.B1(n_65),
.B2(n_78),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_59),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_133),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_76),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_103),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_73),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_1),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_150),
.B1(n_158),
.B2(n_12),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_54),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_151),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_62),
.B1(n_99),
.B2(n_66),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_0),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_153),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_66),
.B(n_22),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_160),
.B(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_157),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_66),
.B(n_23),
.C(n_28),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_164),
.B1(n_13),
.B2(n_14),
.C(n_17),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_1),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_124),
.B1(n_130),
.B2(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_161),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_2),
.B(n_3),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_2),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_3),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_29),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_175),
.C(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_182),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_146),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_153),
.C(n_158),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_35),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g191 ( 
.A(n_183),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_193),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_179),
.C(n_178),
.Y(n_189)
);

XOR2x1_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_166),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_154),
.C(n_140),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_190),
.C(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_175),
.B(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.C(n_198),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_177),
.C(n_172),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_185),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_203),
.B1(n_39),
.B2(n_47),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_204),
.A2(n_36),
.B1(n_46),
.B2(n_45),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_204),
.A2(n_200),
.B1(n_194),
.B2(n_156),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_207),
.B(n_202),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_207),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_209),
.B(n_34),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_32),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_31),
.B(n_44),
.C(n_41),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_21),
.C(n_40),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_50),
.Y(n_215)
);


endmodule