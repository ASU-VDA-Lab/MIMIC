module fake_ariane_3029_n_769 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_769);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_769;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_423;
wire n_347;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_81),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_42),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_24),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_26),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_62),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_59),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_34),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_1),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_66),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_33),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_44),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_121),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_52),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_39),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_32),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_38),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_14),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_56),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_115),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_139),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_25),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_0),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_0),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_1),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_2),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_2),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_145),
.B(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_4),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

AND2x4_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_180),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_146),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_4),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_143),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_158),
.B(n_5),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_6),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_181),
.B1(n_184),
.B2(n_213),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_164),
.B1(n_192),
.B2(n_191),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_147),
.B1(n_192),
.B2(n_191),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_188),
.B1(n_193),
.B2(n_185),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_199),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_201),
.A2(n_188),
.B1(n_183),
.B2(n_176),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_194),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_155),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_156),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_215),
.A2(n_173),
.B1(n_162),
.B2(n_161),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_6),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_160),
.B1(n_159),
.B2(n_157),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_207),
.B(n_7),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g251 ( 
.A(n_208),
.B(n_8),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_253)
);

AOI22x1_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_220),
.Y(n_256)
);

AO22x2_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_16),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_202),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_259)
);

AO22x2_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_227),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_205),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_220),
.B(n_23),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_228),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_35),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_221),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_271)
);

OR2x6_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_43),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_227),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_197),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_227),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_233),
.B(n_55),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_200),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_229),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_230),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_230),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_230),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_230),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_212),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_237),
.B(n_212),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_216),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_212),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_242),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_212),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_212),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_258),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_252),
.B(n_195),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_217),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_278),
.A2(n_196),
.B(n_225),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_272),
.Y(n_315)
);

XOR2x2_ASAP7_75t_L g316 ( 
.A(n_234),
.B(n_224),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_217),
.Y(n_317)
);

NAND2x1p5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_217),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_249),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_196),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_247),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_218),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_260),
.B(n_218),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_241),
.B(n_218),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_264),
.B(n_229),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_254),
.B(n_200),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_254),
.B(n_200),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_272),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_240),
.B(n_200),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_265),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_284),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_297),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_283),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_196),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_224),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_210),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_206),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_206),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_206),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_321),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_288),
.B(n_214),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_206),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_320),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_289),
.B(n_196),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_286),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_298),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g376 ( 
.A(n_282),
.B(n_196),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_209),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_309),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_209),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_335),
.B(n_196),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_343),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_209),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_308),
.B(n_209),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_322),
.B(n_211),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_311),
.B(n_331),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_326),
.B(n_211),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_333),
.B(n_211),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_309),
.B(n_211),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_327),
.B(n_222),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_296),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_329),
.B(n_222),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_287),
.B(n_222),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_294),
.B(n_312),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_323),
.B(n_229),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_302),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_313),
.B(n_222),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_312),
.B(n_195),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_314),
.A2(n_226),
.B(n_223),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_324),
.B(n_223),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_315),
.B(n_57),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_L g407 ( 
.A1(n_335),
.A2(n_195),
.B(n_226),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_303),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_61),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_305),
.B(n_195),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_330),
.B(n_313),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_411),
.B(n_363),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_348),
.B(n_316),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_389),
.Y(n_414)
);

BUFx8_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

BUFx8_ASAP7_75t_SL g416 ( 
.A(n_406),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_336),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_345),
.B(n_351),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_337),
.Y(n_420)
);

NAND2x1p5_ASAP7_75t_L g421 ( 
.A(n_352),
.B(n_315),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_338),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_368),
.B(n_377),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_376),
.B(n_338),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_354),
.B(n_319),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_352),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_337),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_334),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_361),
.B(n_318),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_351),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_402),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_356),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_393),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_361),
.B(n_318),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_307),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_334),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_393),
.B(n_320),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_320),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_402),
.B(n_291),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_400),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_379),
.B(n_318),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_352),
.B(n_397),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_397),
.B(n_291),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_362),
.B(n_304),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_379),
.B(n_316),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_360),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_332),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_378),
.B(n_300),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_406),
.B(n_367),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_369),
.B(n_65),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_195),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_369),
.B(n_67),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_362),
.B(n_223),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_395),
.B(n_226),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_448),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_412),
.B(n_385),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_369),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

BUFx5_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_415),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

BUFx2_ASAP7_75t_R g480 ( 
.A(n_416),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_420),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_451),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_416),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_420),
.B(n_385),
.Y(n_485)
);

BUFx12f_ASAP7_75t_L g486 ( 
.A(n_415),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_392),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_415),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_451),
.A2(n_378),
.B1(n_406),
.B2(n_397),
.Y(n_489)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_431),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_413),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_417),
.A2(n_409),
.B1(n_376),
.B2(n_380),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_433),
.Y(n_494)
);

BUFx8_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_457),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_448),
.Y(n_499)
);

BUFx2_ASAP7_75t_SL g500 ( 
.A(n_423),
.Y(n_500)
);

BUFx8_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

BUFx2_ASAP7_75t_SL g502 ( 
.A(n_462),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_429),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_428),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_436),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_413),
.Y(n_507)
);

BUFx8_ASAP7_75t_L g508 ( 
.A(n_446),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_461),
.A2(n_406),
.B1(n_397),
.B2(n_409),
.Y(n_509)
);

CKINVDCx11_ASAP7_75t_R g510 ( 
.A(n_437),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_436),
.B(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_437),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_459),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

BUFx6f_ASAP7_75t_SL g516 ( 
.A(n_414),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_510),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_453),
.Y(n_518)
);

INVx4_ASAP7_75t_SL g519 ( 
.A(n_516),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_503),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_493),
.A2(n_430),
.B1(n_438),
.B2(n_445),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_486),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_481),
.B(n_434),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_492),
.A2(n_376),
.B1(n_453),
.B2(n_441),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_484),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_473),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_512),
.B(n_426),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_468),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_507),
.A2(n_441),
.B1(n_445),
.B2(n_405),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_469),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_425),
.B1(n_447),
.B2(n_449),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_496),
.A2(n_380),
.B1(n_465),
.B2(n_462),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_493),
.A2(n_495),
.B1(n_508),
.B2(n_490),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_495),
.A2(n_447),
.B1(n_449),
.B2(n_439),
.Y(n_535)
);

CKINVDCx11_ASAP7_75t_R g536 ( 
.A(n_484),
.Y(n_536)
);

BUFx4f_ASAP7_75t_L g537 ( 
.A(n_490),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_482),
.A2(n_424),
.B1(n_347),
.B2(n_349),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_515),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_487),
.B(n_414),
.Y(n_540)
);

BUFx4f_ASAP7_75t_SL g541 ( 
.A(n_483),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_480),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_506),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_471),
.A2(n_380),
.B1(n_465),
.B2(n_462),
.Y(n_544)
);

INVx6_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_470),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_471),
.B(n_444),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_497),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_508),
.A2(n_485),
.B1(n_447),
.B2(n_449),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_472),
.A2(n_424),
.B1(n_347),
.B2(n_349),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_489),
.A2(n_414),
.B1(n_439),
.B2(n_460),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_516),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_514),
.A2(n_439),
.B1(n_450),
.B2(n_392),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_500),
.A2(n_408),
.B1(n_421),
.B2(n_399),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_491),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_510),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_514),
.B(n_387),
.Y(n_559)
);

BUFx10_ASAP7_75t_L g560 ( 
.A(n_480),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_527),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_520),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_533),
.A2(n_471),
.B1(n_401),
.B2(n_476),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_556),
.A2(n_471),
.B1(n_502),
.B2(n_476),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_528),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_534),
.A2(n_509),
.B(n_488),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_537),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_546),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_538),
.A2(n_476),
.B1(n_494),
.B2(n_513),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_505),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_540),
.B(n_511),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_524),
.A2(n_511),
.B1(n_401),
.B2(n_398),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_550),
.A2(n_373),
.B(n_456),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_544),
.A2(n_551),
.B1(n_538),
.B2(n_550),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_529),
.A2(n_398),
.B1(n_476),
.B2(n_455),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_548),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_545),
.A2(n_476),
.B1(n_513),
.B2(n_494),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_521),
.A2(n_398),
.B1(n_476),
.B2(n_455),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_518),
.B(n_390),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_518),
.A2(n_477),
.B1(n_488),
.B2(n_455),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_537),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_543),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_554),
.A2(n_477),
.B(n_421),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_539),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_558),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_553),
.A2(n_346),
.B1(n_452),
.B2(n_432),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_557),
.B(n_387),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_531),
.A2(n_359),
.B1(n_371),
.B2(n_353),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_555),
.B(n_395),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_L g591 ( 
.A1(n_549),
.A2(n_382),
.B(n_408),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_530),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_530),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_541),
.A2(n_346),
.B1(n_452),
.B2(n_442),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_525),
.A2(n_421),
.B1(n_473),
.B2(n_395),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_545),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_535),
.A2(n_371),
.B1(n_370),
.B2(n_353),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_521),
.A2(n_358),
.B1(n_359),
.B2(n_370),
.Y(n_598)
);

INVx5_ASAP7_75t_SL g599 ( 
.A(n_532),
.Y(n_599)
);

INVx5_ASAP7_75t_SL g600 ( 
.A(n_532),
.Y(n_600)
);

AOI222xp33_ASAP7_75t_L g601 ( 
.A1(n_519),
.A2(n_386),
.B1(n_462),
.B2(n_465),
.C1(n_358),
.C2(n_407),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_517),
.A2(n_346),
.B1(n_432),
.B2(n_442),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_517),
.A2(n_465),
.B1(n_407),
.B2(n_374),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_526),
.B(n_469),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

OAI222xp33_ASAP7_75t_L g606 ( 
.A1(n_552),
.A2(n_455),
.B1(n_374),
.B2(n_384),
.C1(n_458),
.C2(n_443),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_519),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_536),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_522),
.A2(n_465),
.B1(n_384),
.B2(n_383),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_574),
.A2(n_465),
.B1(n_391),
.B2(n_383),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_598),
.A2(n_383),
.B1(n_388),
.B2(n_391),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_598),
.A2(n_522),
.B1(n_542),
.B2(n_547),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_573),
.A2(n_394),
.B1(n_388),
.B2(n_391),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_561),
.B(n_526),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_597),
.A2(n_522),
.B1(n_547),
.B2(n_504),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_595),
.A2(n_504),
.B1(n_560),
.B2(n_444),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_597),
.A2(n_344),
.B1(n_479),
.B2(n_435),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_584),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_582),
.B(n_479),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_591),
.A2(n_458),
.B1(n_443),
.B2(n_464),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_603),
.A2(n_404),
.B1(n_499),
.B2(n_475),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_603),
.A2(n_499),
.B1(n_475),
.B2(n_498),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g623 ( 
.A1(n_579),
.A2(n_560),
.B1(n_498),
.B2(n_469),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_605),
.A2(n_607),
.B1(n_571),
.B2(n_602),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_562),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_572),
.A2(n_464),
.B1(n_466),
.B2(n_394),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_587),
.B(n_469),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g629 ( 
.A1(n_566),
.A2(n_386),
.B1(n_396),
.B2(n_394),
.C(n_388),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_588),
.A2(n_601),
.B1(n_578),
.B2(n_580),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_568),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_576),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_592),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_588),
.A2(n_365),
.B1(n_366),
.B2(n_375),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_575),
.A2(n_467),
.B1(n_366),
.B2(n_375),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_570),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_594),
.A2(n_498),
.B1(n_467),
.B2(n_410),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_381),
.B1(n_463),
.B2(n_403),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_569),
.A2(n_381),
.B1(n_463),
.B2(n_498),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_563),
.A2(n_381),
.B1(n_454),
.B2(n_350),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_599),
.A2(n_350),
.B1(n_422),
.B2(n_427),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_590),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_583),
.A2(n_350),
.B(n_372),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_609),
.A2(n_454),
.B1(n_427),
.B2(n_422),
.Y(n_644)
);

OA21x2_ASAP7_75t_L g645 ( 
.A1(n_563),
.A2(n_350),
.B(n_381),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_636),
.B(n_592),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_614),
.B(n_593),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_618),
.B(n_626),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_631),
.B(n_596),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_633),
.B(n_567),
.Y(n_650)
);

NAND4xp25_ASAP7_75t_L g651 ( 
.A(n_619),
.B(n_585),
.C(n_581),
.D(n_609),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_SL g652 ( 
.A(n_610),
.B(n_608),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_645),
.B(n_564),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_610),
.A2(n_600),
.B(n_599),
.Y(n_654)
);

NAND3xp33_ASAP7_75t_L g655 ( 
.A(n_624),
.B(n_604),
.C(n_577),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_628),
.B(n_589),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_642),
.B(n_589),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_625),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_599),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_645),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_645),
.B(n_600),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_613),
.B(n_600),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_630),
.B(n_638),
.Y(n_664)
);

OAI211xp5_ASAP7_75t_L g665 ( 
.A1(n_630),
.A2(n_629),
.B(n_623),
.C(n_637),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_612),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_615),
.B(n_586),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_611),
.B(n_68),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_616),
.B(n_639),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_643),
.B(n_606),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_69),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_622),
.A2(n_381),
.B1(n_454),
.B2(n_427),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_621),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_SL g674 ( 
.A(n_650),
.B(n_617),
.C(n_644),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_646),
.B(n_620),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_664),
.A2(n_670),
.B1(n_669),
.B2(n_652),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_664),
.A2(n_635),
.B1(n_627),
.B2(n_634),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_648),
.B(n_640),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_666),
.B(n_641),
.C(n_634),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_651),
.B(n_422),
.Y(n_680)
);

AOI211xp5_ASAP7_75t_L g681 ( 
.A1(n_665),
.A2(n_652),
.B(n_669),
.C(n_654),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_649),
.B(n_70),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g683 ( 
.A(n_661),
.Y(n_683)
);

OAI211xp5_ASAP7_75t_L g684 ( 
.A1(n_673),
.A2(n_226),
.B(n_223),
.C(n_422),
.Y(n_684)
);

NAND4xp75_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_71),
.C(n_72),
.D(n_73),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_659),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_673),
.A2(n_454),
.B(n_226),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_653),
.A2(n_381),
.B1(n_422),
.B2(n_223),
.Y(n_688)
);

NOR3xp33_ASAP7_75t_L g689 ( 
.A(n_660),
.B(n_74),
.C(n_75),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_648),
.Y(n_690)
);

XOR2x2_ASAP7_75t_L g691 ( 
.A(n_681),
.B(n_655),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_686),
.Y(n_692)
);

NAND4xp75_ASAP7_75t_L g693 ( 
.A(n_674),
.B(n_662),
.C(n_653),
.D(n_663),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_690),
.B(n_656),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_690),
.B(n_647),
.Y(n_695)
);

INVxp67_ASAP7_75t_SL g696 ( 
.A(n_683),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_686),
.Y(n_697)
);

NAND2x1_ASAP7_75t_SL g698 ( 
.A(n_688),
.B(n_672),
.Y(n_698)
);

NAND4xp75_ASAP7_75t_SL g699 ( 
.A(n_682),
.B(n_667),
.C(n_671),
.D(n_668),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_676),
.B(n_658),
.C(n_657),
.Y(n_700)
);

NAND4xp75_ASAP7_75t_L g701 ( 
.A(n_675),
.B(n_659),
.C(n_78),
.D(n_79),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_691),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_694),
.B(n_696),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_692),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_695),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_691),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_705),
.Y(n_707)
);

OA22x2_ASAP7_75t_L g708 ( 
.A1(n_702),
.A2(n_696),
.B1(n_697),
.B2(n_692),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_706),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_703),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_707),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

OAI322xp33_ASAP7_75t_L g713 ( 
.A1(n_709),
.A2(n_700),
.A3(n_704),
.B1(n_679),
.B2(n_680),
.C1(n_694),
.C2(n_699),
.Y(n_713)
);

XOR2x2_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_693),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_712),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_711),
.Y(n_716)
);

OAI31xp33_ASAP7_75t_L g717 ( 
.A1(n_714),
.A2(n_710),
.A3(n_704),
.B(n_689),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

OAI211xp5_ASAP7_75t_L g719 ( 
.A1(n_717),
.A2(n_715),
.B(n_716),
.C(n_713),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_715),
.Y(n_720)
);

AND4x1_ASAP7_75t_L g721 ( 
.A(n_717),
.B(n_687),
.C(n_678),
.D(n_677),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_719),
.B(n_678),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_718),
.A2(n_701),
.B1(n_685),
.B2(n_684),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_720),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_721),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_719),
.A2(n_698),
.B1(n_685),
.B2(n_82),
.C(n_83),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_718),
.B(n_77),
.Y(n_727)
);

NOR2x1_ASAP7_75t_L g728 ( 
.A(n_718),
.B(n_80),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_726),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_724),
.B(n_88),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_728),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_727),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_725),
.B(n_140),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_723),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_722),
.B(n_89),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_731),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_732),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_SL g739 ( 
.A(n_734),
.B(n_90),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_735),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_733),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_729),
.Y(n_742)
);

NAND4xp25_ASAP7_75t_L g743 ( 
.A(n_731),
.B(n_91),
.C(n_92),
.D(n_93),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_731),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_736),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_736),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_740),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_737),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_738),
.Y(n_749)
);

INVxp33_ASAP7_75t_SL g750 ( 
.A(n_741),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_739),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_742),
.B(n_103),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_751),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_749),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_745),
.Y(n_755)
);

OAI22x1_ASAP7_75t_L g756 ( 
.A1(n_748),
.A2(n_743),
.B1(n_744),
.B2(n_107),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_746),
.Y(n_757)
);

AO22x1_ASAP7_75t_L g758 ( 
.A1(n_750),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_754),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_753),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_755),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_760),
.A2(n_757),
.B1(n_756),
.B2(n_752),
.Y(n_762)
);

NOR4xp25_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_752),
.C(n_758),
.D(n_747),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_761),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_762),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_765),
.A2(n_763),
.B1(n_764),
.B2(n_122),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_766),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_767),
.A2(n_119),
.B1(n_120),
.B2(n_124),
.C(n_125),
.Y(n_768)
);

AOI211xp5_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_126),
.B(n_127),
.C(n_128),
.Y(n_769)
);


endmodule