module real_jpeg_20034_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_335, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_335;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_0),
.A2(n_28),
.B1(n_32),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_71),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_71),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_68),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_28),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_2),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_270)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_4),
.A2(n_31),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_4),
.A2(n_31),
.B1(n_52),
.B2(n_53),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_5),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_99),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_99),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_5),
.A2(n_28),
.B1(n_32),
.B2(n_99),
.Y(n_260)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_7),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_93),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_93),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_93),
.Y(n_291)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_22),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_49),
.B(n_52),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_108),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_86),
.B1(n_89),
.B2(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_9),
.B(n_63),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_9),
.A2(n_25),
.B(n_198),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_10),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_105),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_105),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_105),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_11),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_110),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_110),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_110),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_13),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_103),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_103),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_103),
.Y(n_183)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_59),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_14),
.A2(n_25),
.A3(n_48),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_SL g48 ( 
.A(n_17),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_30),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B(n_28),
.C(n_29),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_22),
.A2(n_27),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_22),
.A2(n_27),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_25),
.Y(n_122)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_24),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_24),
.A2(n_29),
.B1(n_107),
.B2(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_24),
.B(n_108),
.Y(n_194)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_28),
.B(n_108),
.CON(n_107),
.SN(n_107)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_34),
.B(n_41),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_76),
.B(n_333),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_72),
.C(n_74),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_42),
.A2(n_43),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_55),
.C(n_64),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_44),
.A2(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_44),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_44),
.A2(n_55),
.B1(n_303),
.B2(n_316),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B(n_54),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_45),
.A2(n_51),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_51),
.B1(n_92),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_45),
.A2(n_51),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_45),
.A2(n_51),
.B1(n_163),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_45),
.A2(n_51),
.B1(n_183),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_45),
.A2(n_51),
.B1(n_98),
.B2(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_45),
.A2(n_51),
.B1(n_94),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_45),
.A2(n_51),
.B1(n_237),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_45),
.A2(n_51),
.B1(n_54),
.B2(n_270),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_47),
.B(n_59),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_48),
.A2(n_50),
.B(n_108),
.C(n_159),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_51),
.B(n_108),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_53),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_55),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_62),
.B(n_63),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_63),
.B1(n_135),
.B2(n_137),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_57),
.A2(n_63),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_61),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_58),
.A2(n_61),
.B1(n_104),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_58),
.A2(n_61),
.B1(n_136),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_58),
.A2(n_61),
.B1(n_118),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_58),
.A2(n_61),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_64),
.A2(n_65),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_70),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_69),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_66),
.A2(n_69),
.B1(n_116),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_66),
.A2(n_69),
.B1(n_244),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_74),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_326),
.B(n_332),
.Y(n_76)
);

OAI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_295),
.A3(n_318),
.B1(n_324),
.B2(n_325),
.C(n_335),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_274),
.B(n_294),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_250),
.B(n_273),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_142),
.B(n_226),
.C(n_249),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_127),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_82),
.B(n_127),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_111),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_95),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_84),
.B(n_95),
.C(n_111),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_85),
.B(n_91),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_88),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_86),
.A2(n_87),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_86),
.A2(n_125),
.B1(n_152),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_86),
.A2(n_89),
.B1(n_155),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_86),
.A2(n_125),
.B1(n_141),
.B2(n_185),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_86),
.A2(n_90),
.B1(n_125),
.B2(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_86),
.A2(n_125),
.B(n_235),
.Y(n_268)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_89),
.B(n_108),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_106),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_120),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_113),
.B(n_119),
.C(n_120),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_123),
.Y(n_131)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.C(n_132),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_128),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_139),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_134),
.B(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_225),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_220),
.B(n_224),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_206),
.B(n_219),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_187),
.B(n_205),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_175),
.B(n_186),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_164),
.B(n_174),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B(n_173),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_182),
.C(n_184),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_195),
.B1(n_203),
.B2(n_204),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_190),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_216),
.C(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_227),
.B(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_248),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_238),
.B2(n_239),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_239),
.C(n_248),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_242),
.C(n_247),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_247),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_272),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_265),
.B2(n_266),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_266),
.C(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_258),
.C(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_260),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_268),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_286),
.B(n_289),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_276),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_292),
.B2(n_293),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_285),
.C(n_293),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_284),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_297),
.C(n_308),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_284),
.A2(n_297),
.B1(n_298),
.B2(n_323),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_284),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_291),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_310),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_310),
.Y(n_325)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_304),
.B1(n_306),
.B2(n_307),
.Y(n_298)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_304),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_304),
.A2(n_307),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_304),
.B(n_312),
.C(n_317),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_308),
.A2(n_309),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_317),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_319),
.B(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_329),
.Y(n_331)
);


endmodule