module fake_netlist_1_3823_n_500 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_500);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_500;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_53), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_60), .Y(n_74) );
INVxp33_ASAP7_75t_L g75 ( .A(n_18), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_57), .Y(n_76) );
INVxp33_ASAP7_75t_SL g77 ( .A(n_7), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_59), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_35), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_54), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_24), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_30), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_4), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_6), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_0), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_20), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_3), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_62), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_14), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_44), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_16), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_67), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_71), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_63), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_23), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_19), .Y(n_102) );
INVxp33_ASAP7_75t_SL g103 ( .A(n_70), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_69), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_32), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_31), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_42), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_13), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_105), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_105), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_76), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_75), .B(n_0), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_96), .B(n_1), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_101), .B(n_1), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_98), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_79), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_74), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_94), .B(n_2), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_96), .Y(n_128) );
NAND2xp33_ASAP7_75t_L g129 ( .A(n_92), .B(n_36), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_84), .B(n_2), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
INVx5_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
INVx2_ASAP7_75t_SL g135 ( .A(n_110), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_122), .B(n_88), .Y(n_137) );
INVx4_ASAP7_75t_SL g138 ( .A(n_116), .Y(n_138) );
CKINVDCx8_ASAP7_75t_R g139 ( .A(n_125), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_121), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_122), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_110), .B(n_81), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_116), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_124), .B(n_88), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_111), .B(n_82), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
BUFx10_ASAP7_75t_L g156 ( .A(n_111), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_139), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_137), .B(n_128), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_156), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_135), .B(n_118), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_135), .B(n_118), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_150), .A2(n_130), .B1(n_115), .B2(n_126), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_150), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_138), .B(n_115), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_133), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_138), .B(n_130), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_150), .A2(n_119), .B1(n_89), .B2(n_90), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_135), .B(n_120), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_156), .B(n_120), .Y(n_175) );
OR2x6_ASAP7_75t_L g176 ( .A(n_150), .B(n_128), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_156), .B(n_103), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_139), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_156), .B(n_107), .Y(n_181) );
NAND3xp33_ASAP7_75t_L g182 ( .A(n_146), .B(n_129), .C(n_132), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_133), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_156), .B(n_120), .Y(n_186) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_137), .B(n_109), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_138), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
BUFx12f_ASAP7_75t_L g191 ( .A(n_176), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
INVx4_ASAP7_75t_L g193 ( .A(n_176), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_165), .B(n_152), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_175), .A2(n_146), .B(n_151), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_189), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_176), .B(n_152), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_175), .B(n_152), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_176), .B(n_138), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_189), .Y(n_201) );
BUFx12f_ASAP7_75t_L g202 ( .A(n_176), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_186), .B(n_146), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_186), .A2(n_146), .B(n_151), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_189), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_187), .A2(n_151), .B1(n_146), .B2(n_138), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_167), .B(n_151), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_164), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_159), .B(n_137), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_162), .A2(n_154), .B1(n_149), .B2(n_132), .Y(n_218) );
OAI22xp33_ASAP7_75t_L g219 ( .A1(n_171), .A2(n_149), .B1(n_154), .B2(n_89), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_162), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_170), .B(n_157), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_201), .Y(n_223) );
NAND2x1_ASAP7_75t_L g224 ( .A(n_205), .B(n_183), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_192), .B(n_189), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_221), .Y(n_226) );
OAI221xp5_ASAP7_75t_L g227 ( .A1(n_216), .A2(n_139), .B1(n_174), .B2(n_161), .C(n_158), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_198), .A2(n_187), .B1(n_170), .B2(n_167), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_221), .A2(n_163), .B1(n_171), .B2(n_172), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_201), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_197), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_197), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_195), .A2(n_163), .B(n_160), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_195), .A2(n_182), .B(n_172), .C(n_170), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_204), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_204), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_198), .B(n_167), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_207), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_192), .A2(n_170), .B1(n_160), .B2(n_182), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_192), .B(n_183), .Y(n_240) );
AOI222xp33_ASAP7_75t_L g241 ( .A1(n_216), .A2(n_161), .B1(n_174), .B2(n_77), .C1(n_93), .C2(n_179), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_191), .Y(n_242) );
INVx6_ASAP7_75t_L g243 ( .A(n_191), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_199), .B(n_177), .Y(n_245) );
OR2x6_ASAP7_75t_L g246 ( .A(n_191), .B(n_188), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_202), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_199), .B(n_157), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_226), .B(n_198), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_226), .B(n_194), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_241), .A2(n_202), .B1(n_192), .B2(n_193), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_229), .A2(n_193), .B1(n_202), .B2(n_219), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_237), .B(n_193), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_227), .A2(n_193), .B1(n_219), .B2(n_194), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_218), .B1(n_200), .B2(n_212), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_242), .A2(n_218), .B1(n_106), .B2(n_200), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_237), .B(n_222), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_228), .A2(n_212), .B1(n_215), .B2(n_207), .C(n_213), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g259 ( .A(n_234), .B(n_131), .C(n_127), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_245), .A2(n_215), .B1(n_213), .B2(n_114), .C(n_123), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g261 ( .A1(n_242), .A2(n_208), .B1(n_209), .B2(n_117), .C(n_114), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_243), .A2(n_200), .B1(n_222), .B2(n_214), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_235), .A2(n_123), .B1(n_117), .B2(n_91), .C(n_95), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_232), .B(n_222), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_200), .B1(n_205), .B2(n_211), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_246), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_243), .A2(n_200), .B1(n_222), .B2(n_214), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_247), .Y(n_269) );
AOI22xp33_ASAP7_75t_SL g270 ( .A1(n_243), .A2(n_211), .B1(n_205), .B2(n_222), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_252), .B(n_246), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_252), .A2(n_246), .B1(n_247), .B2(n_238), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_251), .A2(n_232), .B1(n_236), .B2(n_238), .C(n_104), .Y(n_273) );
AOI211xp5_ASAP7_75t_SL g274 ( .A1(n_256), .A2(n_239), .B(n_236), .C(n_87), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g275 ( .A1(n_255), .A2(n_95), .B1(n_91), .B2(n_102), .C(n_104), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_249), .B(n_246), .Y(n_276) );
OAI211xp5_ASAP7_75t_L g277 ( .A1(n_264), .A2(n_90), .B(n_102), .C(n_113), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_263), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_254), .A2(n_132), .B1(n_240), .B2(n_131), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_263), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_131), .B1(n_127), .B2(n_217), .C(n_157), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_249), .Y(n_282) );
NOR2xp67_ASAP7_75t_L g283 ( .A(n_269), .B(n_205), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_258), .A2(n_131), .B1(n_127), .B2(n_217), .C(n_157), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_269), .B(n_248), .Y(n_286) );
AO21x1_ASAP7_75t_L g287 ( .A1(n_250), .A2(n_225), .B(n_233), .Y(n_287) );
BUFx2_ASAP7_75t_L g288 ( .A(n_267), .Y(n_288) );
NAND4xp25_ASAP7_75t_L g289 ( .A(n_260), .B(n_86), .C(n_82), .D(n_108), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_257), .Y(n_290) );
OAI31xp33_ASAP7_75t_L g291 ( .A1(n_266), .A2(n_86), .A3(n_108), .B(n_100), .Y(n_291) );
OA222x2_ASAP7_75t_L g292 ( .A1(n_250), .A2(n_223), .B1(n_230), .B2(n_85), .C1(n_99), .C2(n_83), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_282), .B(n_267), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_278), .Y(n_295) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_288), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_287), .A2(n_259), .B(n_223), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_290), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_253), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_273), .A2(n_253), .B1(n_268), .B2(n_262), .Y(n_300) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_275), .A2(n_270), .B1(n_261), .B2(n_259), .C(n_83), .Y(n_301) );
NOR3xp33_ASAP7_75t_L g302 ( .A(n_289), .B(n_85), .C(n_99), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_285), .B(n_257), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_271), .A2(n_240), .B1(n_230), .B2(n_224), .Y(n_304) );
OAI21xp33_ASAP7_75t_SL g305 ( .A1(n_271), .A2(n_100), .B(n_97), .Y(n_305) );
OAI33xp33_ASAP7_75t_L g306 ( .A1(n_272), .A2(n_147), .A3(n_142), .B1(n_143), .B2(n_144), .B3(n_140), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_274), .A2(n_224), .B1(n_127), .B2(n_131), .C(n_214), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_291), .A2(n_127), .B1(n_131), .B2(n_214), .C(n_220), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
OA332x1_ASAP7_75t_L g310 ( .A1(n_292), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .C1(n_8), .C2(n_9), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_286), .B(n_127), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_276), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_279), .A2(n_209), .B(n_240), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_276), .B(n_5), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_277), .A2(n_155), .B1(n_142), .B2(n_147), .C(n_206), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_287), .A2(n_144), .B(n_136), .Y(n_316) );
OAI21xp33_ASAP7_75t_L g317 ( .A1(n_279), .A2(n_147), .B(n_142), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_283), .B(n_244), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_281), .B(n_155), .C(n_140), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_284), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_299), .B(n_9), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx3_ASAP7_75t_SL g324 ( .A(n_318), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_312), .B(n_10), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_314), .B(n_10), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_293), .B(n_11), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_299), .B(n_11), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_296), .B(n_12), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_304), .A2(n_136), .B(n_140), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_316), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_318), .B(n_244), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_297), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_303), .B(n_12), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_14), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_305), .B(n_244), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_318), .B(n_15), .Y(n_344) );
AOI321xp33_ASAP7_75t_L g345 ( .A1(n_310), .A2(n_307), .A3(n_302), .B1(n_300), .B2(n_301), .C(n_308), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_306), .A2(n_244), .B(n_210), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_313), .B(n_15), .Y(n_349) );
INVx6_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_317), .B(n_16), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_315), .B(n_17), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_319), .B(n_17), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_314), .B(n_18), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_298), .B(n_19), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_299), .B(n_20), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_299), .B(n_21), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_295), .Y(n_359) );
AOI21xp33_ASAP7_75t_SL g360 ( .A1(n_310), .A2(n_22), .B(n_26), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_295), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_325), .B(n_22), .Y(n_362) );
AO22x1_ASAP7_75t_L g363 ( .A1(n_348), .A2(n_244), .B1(n_211), .B2(n_210), .Y(n_363) );
XNOR2xp5_ASAP7_75t_L g364 ( .A(n_322), .B(n_220), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_347), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_323), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_341), .B(n_143), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_361), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_322), .B(n_27), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_341), .B(n_140), .Y(n_370) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_324), .A2(n_28), .B(n_29), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_331), .B(n_34), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_360), .A2(n_136), .B(n_211), .C(n_148), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_350), .B(n_37), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_342), .B(n_136), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_321), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_342), .B(n_148), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_321), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_361), .Y(n_379) );
AOI22x1_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_203), .B1(n_201), .B2(n_141), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_356), .B(n_141), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_359), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
NAND4xp25_ASAP7_75t_SL g384 ( .A(n_360), .B(n_208), .C(n_190), .D(n_188), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_325), .B(n_38), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_340), .B(n_141), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_358), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_340), .B(n_141), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_358), .B(n_40), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_324), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
XNOR2xp5_ASAP7_75t_L g392 ( .A(n_344), .B(n_220), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_324), .B(n_133), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_133), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_350), .A2(n_203), .B1(n_206), .B2(n_196), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_350), .B(n_41), .Y(n_396) );
OAI31xp33_ASAP7_75t_L g397 ( .A1(n_349), .A2(n_196), .A3(n_206), .B(n_190), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_332), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g399 ( .A1(n_326), .A2(n_349), .A3(n_327), .B1(n_354), .B2(n_339), .C1(n_344), .C2(n_355), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_350), .B(n_155), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_328), .B(n_155), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_348), .B(n_201), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_387), .B(n_357), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_366), .Y(n_404) );
NAND2xp33_ASAP7_75t_SL g405 ( .A(n_390), .B(n_348), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_391), .B(n_329), .Y(n_406) );
NOR2x1_ASAP7_75t_L g407 ( .A(n_373), .B(n_348), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_376), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
NAND4xp25_ASAP7_75t_SL g410 ( .A(n_399), .B(n_328), .C(n_330), .D(n_353), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_374), .B(n_345), .C(n_330), .D(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_382), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_383), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_365), .B(n_368), .Y(n_414) );
CKINVDCx14_ASAP7_75t_R g415 ( .A(n_364), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g416 ( .A1(n_398), .A2(n_353), .B(n_351), .C(n_343), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_400), .B(n_351), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_379), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_365), .B(n_338), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_374), .A2(n_338), .B1(n_337), .B2(n_334), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_390), .B(n_337), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_386), .B(n_335), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
OA22x2_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_333), .B1(n_335), .B2(n_334), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_362), .Y(n_426) );
XNOR2xp5_ASAP7_75t_L g427 ( .A(n_392), .B(n_336), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_393), .Y(n_428) );
XNOR2x1_ASAP7_75t_L g429 ( .A(n_380), .B(n_333), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_371), .A2(n_346), .B(n_196), .C(n_155), .Y(n_430) );
NOR2x1p5_ASAP7_75t_L g431 ( .A(n_362), .B(n_201), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_388), .B(n_45), .Y(n_432) );
OAI32xp33_ASAP7_75t_L g433 ( .A1(n_396), .A2(n_153), .A3(n_48), .B1(n_49), .B2(n_50), .Y(n_433) );
XNOR2x1_ASAP7_75t_L g434 ( .A(n_369), .B(n_46), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_388), .B(n_51), .Y(n_435) );
AOI32xp33_ASAP7_75t_L g436 ( .A1(n_396), .A2(n_153), .A3(n_55), .B1(n_56), .B2(n_58), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_394), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_385), .B(n_52), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_395), .A2(n_153), .B(n_181), .C(n_184), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_381), .B(n_61), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_367), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_370), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_384), .A2(n_153), .B1(n_134), .B2(n_185), .C(n_168), .Y(n_443) );
AOI22x1_ASAP7_75t_L g444 ( .A1(n_385), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_375), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_363), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_372), .A2(n_134), .B1(n_185), .B2(n_178), .C(n_169), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_385), .B(n_68), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_377), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_401), .Y(n_450) );
AOI321xp33_ASAP7_75t_L g451 ( .A1(n_389), .A2(n_72), .A3(n_184), .B1(n_168), .B2(n_169), .C(n_178), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_397), .A2(n_134), .B1(n_184), .B2(n_178), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_387), .A2(n_134), .B1(n_169), .B2(n_180), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_366), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_387), .Y(n_455) );
NOR2xp67_ASAP7_75t_L g456 ( .A(n_390), .B(n_134), .Y(n_456) );
XOR2x2_ASAP7_75t_L g457 ( .A(n_364), .B(n_134), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g458 ( .A1(n_373), .A2(n_180), .B(n_134), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_387), .A2(n_134), .B1(n_180), .B2(n_350), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_387), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_379), .B(n_365), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_414), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_410), .A2(n_456), .B(n_446), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_414), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_455), .B(n_460), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_460), .Y(n_466) );
AOI211xp5_ASAP7_75t_L g467 ( .A1(n_410), .A2(n_411), .B(n_416), .C(n_459), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_418), .A2(n_415), .B1(n_406), .B2(n_403), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_431), .A2(n_407), .B1(n_426), .B2(n_424), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_461), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_405), .A2(n_436), .B(n_426), .C(n_424), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_428), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_453), .A2(n_421), .B(n_448), .C(n_450), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_461), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_451), .B(n_443), .C(n_452), .D(n_438), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_428), .A2(n_422), .B1(n_409), .B2(n_412), .C(n_404), .Y(n_476) );
AND3x2_ASAP7_75t_L g477 ( .A(n_437), .B(n_434), .C(n_417), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_472), .B(n_423), .Y(n_478) );
OAI211xp5_ASAP7_75t_L g479 ( .A1(n_471), .A2(n_444), .B(n_430), .C(n_458), .Y(n_479) );
NAND4xp75_ASAP7_75t_L g480 ( .A(n_463), .B(n_435), .C(n_432), .D(n_440), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_467), .A2(n_433), .B(n_430), .C(n_432), .Y(n_481) );
AOI21xp33_ASAP7_75t_SL g482 ( .A1(n_469), .A2(n_429), .B(n_425), .Y(n_482) );
XNOR2xp5_ASAP7_75t_L g483 ( .A(n_477), .B(n_427), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_468), .A2(n_435), .B(n_422), .C(n_441), .Y(n_484) );
OAI322xp33_ASAP7_75t_L g485 ( .A1(n_472), .A2(n_419), .A3(n_420), .B1(n_408), .B2(n_413), .C1(n_454), .C2(n_425), .Y(n_485) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_473), .A2(n_449), .B(n_445), .C(n_442), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_482), .B(n_466), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_481), .B(n_465), .C(n_475), .D(n_476), .Y(n_488) );
XOR2xp5_ASAP7_75t_L g489 ( .A(n_483), .B(n_457), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_486), .B(n_439), .C(n_447), .D(n_474), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_478), .B(n_470), .Y(n_491) );
NAND3xp33_ASAP7_75t_SL g492 ( .A(n_489), .B(n_479), .C(n_484), .Y(n_492) );
OR4x2_ASAP7_75t_L g493 ( .A(n_487), .B(n_480), .C(n_485), .D(n_479), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_491), .Y(n_494) );
XOR2xp5_ASAP7_75t_L g495 ( .A(n_492), .B(n_488), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_494), .B(n_490), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_496), .B(n_492), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_497), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g499 ( .A1(n_498), .A2(n_493), .B1(n_495), .B2(n_464), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_499), .A2(n_462), .B(n_457), .Y(n_500) );
endmodule