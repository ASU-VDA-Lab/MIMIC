module fake_ariane_2813_n_427 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_427);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_427;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_261;
wire n_220;
wire n_370;
wire n_189;
wire n_286;
wire n_424;
wire n_387;
wire n_406;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_410;
wire n_379;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_285;
wire n_186;
wire n_202;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_152;
wire n_405;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_401;
wire n_267;
wire n_335;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_398;
wire n_210;
wire n_200;
wire n_253;
wire n_166;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_369;
wire n_224;
wire n_420;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_303;
wire n_168;
wire n_206;
wire n_352;
wire n_365;
wire n_238;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_390;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_413;
wire n_392;
wire n_376;
wire n_221;
wire n_321;
wire n_361;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_371;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_284;
wire n_249;
wire n_355;
wire n_212;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_409;
wire n_171;
wire n_384;
wire n_182;
wire n_316;
wire n_196;
wire n_407;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_298;
wire n_415;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_378;
wire n_150;
wire n_375;
wire n_324;
wire n_337;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_358;
wire n_263;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_191;
wire n_382;
wire n_211;
wire n_408;
wire n_322;
wire n_251;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_31),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_30),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_55),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_33),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_114),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_39),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_38),
.B(n_65),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_11),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_93),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_17),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g177 ( 
.A(n_19),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_5),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_62),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_27),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_101),
.B(n_97),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_71),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_22),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_56),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_68),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_106),
.B(n_34),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_L g203 ( 
.A(n_72),
.B(n_63),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_42),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_126),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_53),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_133),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_46),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_25),
.B(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_85),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_47),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g221 ( 
.A(n_52),
.B(n_115),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_20),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_48),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_24),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_70),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_3),
.Y(n_234)
);

INVxp33_ASAP7_75t_SL g235 ( 
.A(n_80),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_98),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_77),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_122),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_127),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_107),
.B(n_79),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_105),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_69),
.B(n_81),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_L g247 ( 
.A(n_49),
.B(n_15),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_23),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_41),
.B(n_10),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_28),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_110),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_61),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_0),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_9),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_50),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_89),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_148),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_180),
.B(n_2),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_183),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_153),
.B(n_18),
.Y(n_264)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_192),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_151),
.B(n_21),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_149),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_150),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_182),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_152),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_156),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_154),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_26),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

OR2x6_ASAP7_75t_L g278 ( 
.A(n_203),
.B(n_29),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_160),
.B(n_44),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_161),
.B(n_45),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_58),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_190),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_164),
.B(n_66),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_158),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_168),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_193),
.B(n_73),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_74),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_163),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_169),
.B(n_75),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_173),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_206),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_181),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_184),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_186),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_187),
.B(n_188),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_88),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_177),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_299)
);

BUFx4f_ASAP7_75t_L g300 ( 
.A(n_189),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_155),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_194),
.B(n_102),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_197),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_200),
.B(n_257),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_235),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_308)
);

NOR2x1p5_ASAP7_75t_L g309 ( 
.A(n_167),
.B(n_116),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_208),
.B(n_120),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_209),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_262),
.B(n_159),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_210),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_261),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_211),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_172),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_297),
.A2(n_246),
.B(n_234),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_300),
.B(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_303),
.B(n_256),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_217),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_289),
.B(n_254),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_260),
.A2(n_218),
.B(n_249),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_252),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_290),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_195),
.B(n_232),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_179),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_239),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_214),
.C(n_207),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_178),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_215),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_280),
.A2(n_284),
.B(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_229),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_286),
.A2(n_199),
.B(n_174),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_237),
.B(n_233),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_269),
.B(n_251),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_295),
.A2(n_248),
.B(n_227),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_213),
.C(n_226),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_279),
.A2(n_220),
.B(n_223),
.C(n_225),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_266),
.A2(n_247),
.B(n_221),
.Y(n_342)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_204),
.B(n_201),
.C(n_243),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_242),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_240),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

OR2x6_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_293),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_309),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_301),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_317),
.A2(n_276),
.B(n_275),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_281),
.B(n_288),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_338),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_334),
.A2(n_308),
.B(n_299),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_342),
.Y(n_354)
);

OR2x6_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_278),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_311),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_343),
.B(n_171),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_258),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_332),
.B(n_331),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_304),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_292),
.B(n_185),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_323),
.A2(n_294),
.B(n_170),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_266),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_267),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_331),
.B(n_285),
.Y(n_367)
);

CKINVDCx8_ASAP7_75t_R g368 ( 
.A(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_360),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_312),
.Y(n_373)
);

HB1xp67_ASAP7_75t_SL g374 ( 
.A(n_368),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_346),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_347),
.Y(n_377)
);

INVx5_ASAP7_75t_SL g378 ( 
.A(n_367),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g379 ( 
.A1(n_363),
.A2(n_341),
.B(n_336),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_354),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_370),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_320),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_352),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_348),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_350),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_355),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_373),
.B(n_365),
.Y(n_396)
);

AOI221xp5_ASAP7_75t_L g397 ( 
.A1(n_371),
.A2(n_339),
.B1(n_351),
.B2(n_271),
.C(n_327),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_386),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_355),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_271),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_230),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_392),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_378),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_391),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_378),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_401),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_407),
.B(n_394),
.Y(n_410)
);

NOR2x1_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_395),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_399),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_396),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_329),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_413),
.A2(n_374),
.B1(n_405),
.B2(n_402),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_219),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_202),
.Y(n_418)
);

OA22x2_ASAP7_75t_L g419 ( 
.A1(n_416),
.A2(n_414),
.B1(n_411),
.B2(n_212),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_417),
.B(n_415),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_419),
.A2(n_418),
.B1(n_238),
.B2(n_236),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_421),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_420),
.C(n_397),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_196),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_166),
.B(n_379),
.Y(n_425)
);

OA22x2_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_176),
.B1(n_224),
.B2(n_222),
.Y(n_426)
);

OAI221xp5_ASAP7_75t_R g427 ( 
.A1(n_426),
.A2(n_424),
.B1(n_137),
.B2(n_138),
.C(n_142),
.Y(n_427)
);


endmodule