module fake_jpeg_1918_n_665 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_665);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_665;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_653;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_60),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_19),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_75),
.Y(n_131)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_64),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_69),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_70),
.Y(n_197)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_102),
.Y(n_152)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_74),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_19),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_24),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g183 ( 
.A(n_76),
.Y(n_183)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_24),
.B(n_18),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g138 ( 
.A(n_87),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_88),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_89),
.Y(n_212)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_92),
.Y(n_215)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_93),
.Y(n_222)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_18),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_57),
.B(n_18),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_106),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_26),
.Y(n_97)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_52),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_30),
.B(n_17),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_40),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_117),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_57),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_33),
.B(n_51),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_121),
.Y(n_162)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_33),
.B(n_0),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_130),
.Y(n_181)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_41),
.Y(n_127)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_127),
.Y(n_202)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_39),
.B(n_0),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_64),
.A2(n_56),
.B1(n_54),
.B2(n_34),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_136),
.A2(n_34),
.B1(n_56),
.B2(n_47),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_145),
.B(n_173),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_147),
.B(n_151),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_166),
.B(n_178),
.Y(n_274)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_49),
.C(n_35),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_38),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_39),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_180),
.B(n_182),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_43),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_97),
.B(n_43),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_191),
.B(n_204),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_88),
.A2(n_28),
.B1(n_54),
.B2(n_48),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_200),
.B1(n_224),
.B2(n_34),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_114),
.B(n_43),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_203),
.Y(n_230)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_89),
.A2(n_28),
.B1(n_54),
.B2(n_48),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_63),
.B(n_51),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_116),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_74),
.B(n_50),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_127),
.B(n_50),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_84),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_68),
.B(n_49),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_36),
.Y(n_245)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_104),
.Y(n_221)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_92),
.A2(n_22),
.B1(n_48),
.B2(n_47),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_69),
.B(n_35),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_227),
.Y(n_270)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_99),
.Y(n_226)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_70),
.B(n_36),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_181),
.A2(n_85),
.B1(n_83),
.B2(n_109),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_228),
.A2(n_261),
.B1(n_295),
.B2(n_136),
.Y(n_346)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_229),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_231),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_234),
.A2(n_235),
.B1(n_263),
.B2(n_276),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_192),
.A2(n_165),
.B1(n_155),
.B2(n_157),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_236),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_237),
.B(n_283),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_238),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_239),
.Y(n_361)
);

CKINVDCx9p33_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

INVx8_ASAP7_75t_L g351 ( 
.A(n_240),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_131),
.B(n_22),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_265),
.C(n_150),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_245),
.B(n_249),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_247),
.B(n_269),
.Y(n_338)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_248),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_162),
.B(n_38),
.Y(n_249)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_251),
.Y(n_340)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_144),
.Y(n_256)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_256),
.Y(n_356)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_164),
.Y(n_258)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_152),
.Y(n_259)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_149),
.Y(n_260)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_181),
.A2(n_105),
.B1(n_56),
.B2(n_47),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_145),
.B(n_28),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_262),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_168),
.A2(n_23),
.B1(n_22),
.B2(n_29),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g265 ( 
.A(n_195),
.B(n_23),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_183),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_271),
.Y(n_369)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_214),
.Y(n_273)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_133),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_275),
.B(n_278),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_188),
.A2(n_23),
.B1(n_29),
.B2(n_3),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_205),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_277),
.B(n_279),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_162),
.B(n_1),
.Y(n_278)
);

OR2x2_ASAP7_75t_SL g279 ( 
.A(n_154),
.B(n_169),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_281),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_154),
.B(n_1),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_182),
.B(n_1),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_284),
.Y(n_365)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_139),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_173),
.B(n_2),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_288),
.Y(n_313)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_286),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_207),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_146),
.B(n_2),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_289),
.Y(n_324)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_176),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_177),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_291),
.Y(n_347)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_141),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_292),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_197),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_299),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_148),
.A2(n_29),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_159),
.B(n_2),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_296),
.B(n_7),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_225),
.B(n_2),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_298),
.A2(n_305),
.B1(n_4),
.B2(n_6),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_197),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_140),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_161),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_189),
.Y(n_312)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_187),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_306),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_150),
.B(n_4),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_186),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_142),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_212),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_339),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_230),
.A2(n_226),
.B1(n_224),
.B2(n_193),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_314),
.A2(n_321),
.B1(n_327),
.B2(n_330),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_316),
.A2(n_7),
.B(n_8),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_270),
.A2(n_184),
.B1(n_215),
.B2(n_213),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_244),
.A2(n_215),
.B1(n_213),
.B2(n_212),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_283),
.A2(n_200),
.B1(n_170),
.B2(n_211),
.Y(n_330)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

AO22x1_ASAP7_75t_L g339 ( 
.A1(n_262),
.A2(n_179),
.B1(n_202),
.B2(n_222),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_255),
.B(n_265),
.C(n_279),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_355),
.C(n_362),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_346),
.B(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_265),
.B(n_211),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_350),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_171),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_250),
.B(n_156),
.C(n_198),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_209),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_360),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_274),
.B(n_201),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_156),
.C(n_201),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g363 ( 
.A1(n_234),
.A2(n_185),
.B1(n_206),
.B2(n_156),
.Y(n_363)
);

AO22x2_ASAP7_75t_L g364 ( 
.A1(n_234),
.A2(n_158),
.B1(n_175),
.B2(n_163),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_366),
.B(n_371),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_247),
.A2(n_175),
.B1(n_163),
.B2(n_158),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_233),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_342),
.A2(n_235),
.B1(n_286),
.B2(n_263),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_385),
.B1(n_413),
.B2(n_339),
.Y(n_444)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_381),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_238),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_342),
.A2(n_302),
.B1(n_276),
.B2(n_258),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_232),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_401),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_388),
.Y(n_430)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_291),
.B1(n_289),
.B2(n_252),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_390),
.A2(n_318),
.B1(n_324),
.B2(n_347),
.Y(n_426)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_348),
.A2(n_241),
.B1(n_246),
.B2(n_257),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_393),
.A2(n_394),
.B1(n_398),
.B2(n_340),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_357),
.A2(n_257),
.B1(n_293),
.B2(n_294),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_320),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_400),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_350),
.A2(n_293),
.B1(n_299),
.B2(n_256),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_399),
.A2(n_409),
.B1(n_414),
.B2(n_352),
.Y(n_442)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_273),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_402),
.B(n_407),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_329),
.B(n_240),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_404),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_349),
.B(n_272),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_313),
.B(n_268),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_406),
.B(n_408),
.Y(n_433)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_353),
.B(n_231),
.Y(n_408)
);

CKINVDCx12_ASAP7_75t_R g409 ( 
.A(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_264),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_412),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_313),
.B(n_292),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_415),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_333),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_332),
.A2(n_310),
.B1(n_251),
.B2(n_267),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g414 ( 
.A1(n_315),
.A2(n_253),
.B1(n_243),
.B2(n_295),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_371),
.B(n_243),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_312),
.A2(n_364),
.B(n_363),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_363),
.B(n_364),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_326),
.B(n_354),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_417),
.B(n_319),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_366),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_333),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_319),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_316),
.C(n_341),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_437),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_423),
.A2(n_427),
.B(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_359),
.B(n_339),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_383),
.A2(n_375),
.B(n_416),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_449),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_405),
.B(n_331),
.C(n_362),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_375),
.A2(n_364),
.B(n_363),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_438),
.A2(n_367),
.B(n_380),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_386),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_396),
.A2(n_321),
.B1(n_327),
.B2(n_334),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_440),
.A2(n_444),
.B1(n_452),
.B2(n_396),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_SL g476 ( 
.A1(n_442),
.A2(n_451),
.B(n_458),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_338),
.C(n_369),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_445),
.B(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_446),
.B(n_410),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_375),
.B(n_412),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_453),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_378),
.A2(n_370),
.B1(n_343),
.B2(n_335),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_396),
.A2(n_318),
.B1(n_368),
.B2(n_317),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_343),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_379),
.B(n_325),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_455),
.B(n_340),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_400),
.B(n_317),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_391),
.A2(n_337),
.B(n_345),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_376),
.B(n_337),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_387),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_462),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_463),
.B(n_425),
.Y(n_514)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_453),
.Y(n_464)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_449),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_481),
.Y(n_498)
);

OR2x4_ASAP7_75t_L g466 ( 
.A(n_432),
.B(n_373),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_466),
.A2(n_490),
.B(n_452),
.Y(n_513)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_424),
.Y(n_467)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_467),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_468),
.B(n_478),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_444),
.A2(n_372),
.B1(n_389),
.B2(n_376),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_469),
.A2(n_482),
.B1(n_484),
.B2(n_486),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_455),
.Y(n_470)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_479),
.C(n_483),
.Y(n_517)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_424),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_472),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_413),
.B1(n_372),
.B2(n_385),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_473),
.A2(n_480),
.B1(n_435),
.B2(n_431),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_456),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_428),
.B(n_393),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_429),
.A2(n_391),
.B1(n_384),
.B2(n_398),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_428),
.A2(n_394),
.B1(n_407),
.B2(n_377),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_450),
.Y(n_483)
);

OAI22x1_ASAP7_75t_SL g484 ( 
.A1(n_429),
.A2(n_403),
.B1(n_392),
.B2(n_381),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_402),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_489),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_423),
.A2(n_340),
.B1(n_311),
.B2(n_356),
.Y(n_486)
);

INVx13_ASAP7_75t_L g487 ( 
.A(n_447),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_487),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_445),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_493),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g492 ( 
.A(n_425),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_492),
.Y(n_519)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_457),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_441),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_494),
.B(n_495),
.Y(n_521)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_438),
.A2(n_311),
.B1(n_356),
.B2(n_388),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_496),
.A2(n_422),
.B1(n_443),
.B2(n_448),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_437),
.C(n_459),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_504),
.C(n_474),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_466),
.A2(n_458),
.B(n_427),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_500),
.A2(n_515),
.B(n_461),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_480),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_502),
.A2(n_461),
.B1(n_482),
.B2(n_486),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_460),
.B(n_431),
.C(n_420),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_433),
.Y(n_507)
);

INVxp33_ASAP7_75t_SL g538 ( 
.A(n_507),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_479),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_508),
.B(n_509),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_469),
.B(n_433),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_481),
.B(n_446),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_510),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_420),
.Y(n_512)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_512),
.A2(n_514),
.B(n_518),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_513),
.A2(n_488),
.B(n_490),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_478),
.A2(n_435),
.B1(n_439),
.B2(n_422),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_395),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_491),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_479),
.Y(n_537)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_522),
.Y(n_546)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_488),
.A2(n_443),
.B(n_430),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_523),
.A2(n_529),
.B1(n_467),
.B2(n_472),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_468),
.A2(n_430),
.B1(n_399),
.B2(n_388),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_526),
.A2(n_531),
.B1(n_484),
.B2(n_496),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_471),
.B(n_399),
.Y(n_527)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_464),
.B(n_434),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_528),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_473),
.A2(n_367),
.B1(n_239),
.B2(n_323),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_323),
.Y(n_530)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_530),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_478),
.A2(n_7),
.B1(n_12),
.B2(n_13),
.Y(n_531)
);

XNOR2x1_ASAP7_75t_L g570 ( 
.A(n_533),
.B(n_523),
.Y(n_570)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_498),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_535),
.B(n_560),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_536),
.A2(n_559),
.B1(n_531),
.B2(n_503),
.Y(n_581)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_537),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_544),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_497),
.B(n_474),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_530),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_542),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_545),
.A2(n_549),
.B1(n_562),
.B2(n_563),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_495),
.Y(n_547)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_547),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_494),
.Y(n_548)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_548),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_519),
.B(n_476),
.Y(n_551)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_551),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_519),
.B(n_462),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_553),
.B(n_554),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_511),
.B(n_462),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_511),
.B(n_462),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_555),
.B(n_561),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_500),
.A2(n_465),
.B(n_487),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_556),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_504),
.B(n_12),
.C(n_13),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_558),
.B(n_499),
.C(n_525),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_515),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_559)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_513),
.A2(n_12),
.B(n_13),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_521),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_502),
.A2(n_14),
.B1(n_524),
.B2(n_516),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_521),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_562),
.A2(n_516),
.B1(n_498),
.B2(n_524),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_564),
.A2(n_573),
.B1(n_559),
.B2(n_552),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_557),
.A2(n_514),
.B1(n_499),
.B2(n_506),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_569),
.B(n_571),
.Y(n_599)
);

XNOR2x1_ASAP7_75t_L g603 ( 
.A(n_570),
.B(n_574),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_540),
.B(n_501),
.C(n_508),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_572),
.B(n_576),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_546),
.A2(n_524),
.B1(n_523),
.B2(n_517),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g574 ( 
.A(n_541),
.B(n_544),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_538),
.A2(n_529),
.B1(n_522),
.B2(n_523),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_577),
.B(n_578),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_527),
.C(n_526),
.Y(n_578)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_523),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_586),
.B(n_587),
.C(n_554),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_542),
.B(n_523),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_583),
.A2(n_533),
.B(n_537),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_588),
.A2(n_593),
.B(n_597),
.Y(n_621)
);

INVx13_ASAP7_75t_L g589 ( 
.A(n_585),
.Y(n_589)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_589),
.Y(n_616)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_583),
.Y(n_591)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_591),
.Y(n_619)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_566),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_592),
.B(n_594),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_584),
.A2(n_543),
.B(n_563),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_579),
.A2(n_561),
.B1(n_546),
.B2(n_545),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_596),
.Y(n_622)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_581),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_543),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_568),
.A2(n_549),
.B1(n_536),
.B2(n_550),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_601),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_601),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_575),
.A2(n_550),
.B1(n_552),
.B2(n_555),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_605),
.A2(n_596),
.B1(n_590),
.B2(n_591),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_580),
.B(n_539),
.C(n_547),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_606),
.B(n_607),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_565),
.A2(n_539),
.B(n_553),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_534),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_611),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_609),
.B(n_615),
.Y(n_633)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_610),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_607),
.B(n_534),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_599),
.B(n_582),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_614),
.B(n_617),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_SL g615 ( 
.A(n_603),
.B(n_580),
.C(n_572),
.Y(n_615)
);

XOR2x1_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_603),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_604),
.B(n_578),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_593),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_602),
.B(n_574),
.C(n_576),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_623),
.B(n_624),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_605),
.A2(n_565),
.B1(n_564),
.B2(n_573),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_621),
.A2(n_619),
.B1(n_597),
.B2(n_592),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_634),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_616),
.B(n_590),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_631),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_595),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_594),
.Y(n_632)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_632),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_609),
.B(n_571),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_613),
.B(n_598),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_635),
.B(n_636),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_613),
.B(n_600),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_637),
.B(n_624),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_622),
.B(n_503),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_638),
.A2(n_548),
.B(n_558),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_625),
.A2(n_623),
.B(n_612),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_640),
.A2(n_648),
.B(n_633),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_625),
.A2(n_627),
.B(n_621),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_641),
.B(n_646),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_628),
.B(n_627),
.C(n_633),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_642),
.B(n_647),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_637),
.A2(n_610),
.B(n_617),
.Y(n_648)
);

INVx11_ASAP7_75t_L g649 ( 
.A(n_643),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_649),
.B(n_652),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_645),
.B(n_630),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_644),
.B(n_630),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_653),
.B(n_639),
.Y(n_656)
);

INVxp33_ASAP7_75t_L g657 ( 
.A(n_654),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_656),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_654),
.B(n_639),
.C(n_586),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_658),
.B(n_651),
.C(n_650),
.Y(n_660)
);

AOI31xp33_ASAP7_75t_L g661 ( 
.A1(n_660),
.A2(n_655),
.A3(n_649),
.B(n_657),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_661),
.B(n_659),
.C(n_651),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_662),
.Y(n_663)
);

AOI322xp5_ASAP7_75t_L g664 ( 
.A1(n_663),
.A2(n_589),
.A3(n_525),
.B1(n_505),
.B2(n_570),
.C1(n_560),
.C2(n_587),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_664),
.B(n_505),
.Y(n_665)
);


endmodule