module fake_jpeg_30078_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_SL g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_33),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_84),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_77),
.Y(n_95)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_60),
.B1(n_53),
.B2(n_69),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_77),
.Y(n_122)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_65),
.B1(n_66),
.B2(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_62),
.B1(n_56),
.B2(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_68),
.C(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_108),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_61),
.B1(n_56),
.B2(n_67),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_114),
.B1(n_117),
.B2(n_102),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_19),
.B(n_40),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_79),
.B1(n_75),
.B2(n_63),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_54),
.C(n_55),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_65),
.B1(n_74),
.B2(n_73),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_122),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_59),
.B1(n_76),
.B2(n_57),
.Y(n_121)
);

OA21x2_ASAP7_75t_R g146 ( 
.A1(n_121),
.A2(n_4),
.B(n_5),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_76),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_123),
.A2(n_94),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_128),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_139),
.Y(n_163)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_135),
.B1(n_138),
.B2(n_7),
.Y(n_156)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_1),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_45),
.B1(n_38),
.B2(n_37),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_1),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_146),
.B1(n_10),
.B2(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_36),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_7),
.Y(n_158)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_35),
.B(n_34),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_31),
.B(n_30),
.Y(n_149)
);

NOR2x1p5_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_138),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_29),
.C(n_26),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_151),
.C(n_157),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_24),
.C(n_8),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_131),
.C(n_142),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_14),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_162),
.B1(n_164),
.B2(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_135),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_167),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_152),
.B1(n_153),
.B2(n_148),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_165),
.B1(n_157),
.B2(n_170),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_176),
.B(n_173),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_175),
.B(n_150),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_172),
.B(n_149),
.C(n_151),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_149),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_154),
.A3(n_161),
.B1(n_132),
.B2(n_143),
.C1(n_134),
.C2(n_17),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_130),
.B(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_130),
.C(n_17),
.Y(n_186)
);


endmodule