module fake_jpeg_21165_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_30),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_15),
.B1(n_25),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_15),
.B1(n_25),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_31),
.B1(n_22),
.B2(n_40),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_15),
.B1(n_25),
.B2(n_41),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_76),
.B1(n_54),
.B2(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_36),
.B1(n_41),
.B2(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_61),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_35),
.CON(n_59),
.SN(n_59)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_62),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_33),
.B1(n_39),
.B2(n_29),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_24),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_38),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_51),
.B1(n_44),
.B2(n_37),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_38),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_77),
.A3(n_59),
.B1(n_70),
.B2(n_66),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_34),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_34),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_26),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_21),
.B1(n_54),
.B2(n_18),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_98),
.B1(n_91),
.B2(n_72),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_78),
.B1(n_63),
.B2(n_72),
.Y(n_110)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_54),
.C(n_32),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_27),
.C(n_19),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_17),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_23),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_62),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_32),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_28),
.B1(n_84),
.B2(n_3),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_113),
.B(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_112),
.B1(n_83),
.B2(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_72),
.B1(n_79),
.B2(n_32),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_23),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_116),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_55),
.B1(n_67),
.B2(n_30),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_30),
.B(n_18),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_12),
.B(n_11),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_11),
.C(n_10),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_93),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_19),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_23),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_103),
.C(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_28),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_124),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_115),
.C(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_83),
.B1(n_86),
.B2(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_130),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_27),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_133),
.A2(n_137),
.B(n_119),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_107),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_113),
.B1(n_110),
.B2(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_142),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_99),
.B1(n_101),
.B2(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_99),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_159),
.B1(n_133),
.B2(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_126),
.C(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_116),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_162),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_170),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_129),
.B1(n_136),
.B2(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_150),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_131),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_150),
.B1(n_158),
.B2(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_168),
.B1(n_166),
.B2(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_177),
.B(n_180),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_137),
.B(n_132),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_178),
.A2(n_168),
.B(n_143),
.Y(n_181)
);

OAI21x1_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_144),
.B(n_128),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_178),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_104),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_105),
.B(n_2),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_170),
.C(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_1),
.Y(n_192)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_162),
.A3(n_154),
.B1(n_153),
.B2(n_105),
.C(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_173),
.B(n_2),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_192),
.B(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_186),
.B1(n_183),
.B2(n_5),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_194),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_4),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_8),
.B(n_5),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_195),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_199),
.B(n_195),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_6),
.Y(n_203)
);


endmodule