module fake_netlist_5_479_n_1275 (n_137, n_294, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_286, n_122, n_282, n_10, n_24, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_9, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1275);

input n_137;
input n_294;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_9;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1275;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_1270;
wire n_582;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_833;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1136;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_318;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_903;
wire n_740;
wire n_384;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_226),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_241),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_227),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_155),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_125),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_74),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_149),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_152),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_202),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_188),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_29),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_209),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_163),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_162),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_94),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_128),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_295),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_232),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_234),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_302),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_59),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_316),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_238),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_81),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_160),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_233),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_190),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_236),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_240),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_97),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_75),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_161),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_55),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_104),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_48),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_140),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_294),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_182),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_15),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_74),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_144),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_113),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_138),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_245),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_166),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_62),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_158),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_181),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_82),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_210),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_230),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_109),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_246),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_105),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_257),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_39),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_231),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_169),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_110),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_243),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_203),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_267),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_21),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_103),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_95),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_300),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_206),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_168),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_252),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_298),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_86),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_280),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_59),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_221),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_65),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_239),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_291),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_13),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_146),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_165),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_145),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_235),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_180),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_137),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_301),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_79),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_119),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_34),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_199),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_164),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_178),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_256),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_127),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_200),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_132),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_237),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_36),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_157),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_141),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_34),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_136),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_314),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_150),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_223),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_36),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_112),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_64),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_224),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_194),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_249),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_11),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_53),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_80),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_131),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_45),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_277),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_217),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_49),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_290),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_62),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_185),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_273),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_156),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_253),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_9),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_28),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_75),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_215),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_117),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_311),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_310),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_254),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_29),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_222),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_153),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_102),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_216),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_9),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_244),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_54),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_14),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_25),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_115),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_195),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_139),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_134),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_130),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_24),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_214),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_90),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_196),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_315),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_284),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_250),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_24),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_7),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_307),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_65),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_80),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_308),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_1),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_133),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_292),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_56),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_122),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_64),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_58),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_304),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_204),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_92),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_309),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_78),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_108),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_259),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_14),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_7),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_47),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_143),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_71),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_258),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_148),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_312),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_255),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_364),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_336),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_356),
.B(n_0),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_364),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_363),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_336),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_352),
.B(n_426),
.Y(n_518)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_336),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_495),
.B(n_0),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_1),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_336),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_366),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_352),
.B(n_2),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_366),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_447),
.B(n_2),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_394),
.Y(n_529)
);

BUFx8_ASAP7_75t_SL g530 ( 
.A(n_454),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_394),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_355),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_378),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_380),
.B(n_445),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_355),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_374),
.B(n_3),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_390),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_363),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_456),
.B(n_3),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_361),
.B(n_4),
.Y(n_540)
);

BUFx8_ASAP7_75t_SL g541 ( 
.A(n_507),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_390),
.B(n_5),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_322),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_5),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_393),
.B(n_6),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_414),
.B(n_6),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_509),
.B(n_8),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_475),
.B(n_10),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_355),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_355),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_415),
.B(n_10),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_342),
.B(n_11),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_322),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_388),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_342),
.B(n_12),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_365),
.B(n_12),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_322),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_365),
.B(n_13),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_317),
.Y(n_560)
);

CKINVDCx11_ASAP7_75t_R g561 ( 
.A(n_448),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_427),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_415),
.B(n_468),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_423),
.B(n_15),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_423),
.B(n_16),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_355),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_468),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_355),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_474),
.B(n_16),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_427),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_427),
.B(n_17),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_359),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_437),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_492),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_388),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_328),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_460),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_462),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_462),
.B(n_17),
.Y(n_584)
);

NOR2x1_ASAP7_75t_L g585 ( 
.A(n_351),
.B(n_18),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_371),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_477),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_376),
.Y(n_588)
);

INVx5_ASAP7_75t_L g589 ( 
.A(n_477),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_481),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_320),
.B(n_18),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_384),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_373),
.B(n_19),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_392),
.B(n_19),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_345),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_324),
.B(n_20),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_331),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_333),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_505),
.B(n_20),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_481),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_357),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_435),
.B(n_21),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_443),
.B(n_446),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_339),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_340),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_469),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_318),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_470),
.Y(n_608)
);

INVx5_ASAP7_75t_L g609 ( 
.A(n_382),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_570),
.A2(n_329),
.B1(n_341),
.B2(n_332),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_518),
.A2(n_399),
.B1(n_401),
.B2(n_389),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_534),
.B(n_419),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_537),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_542),
.A2(n_500),
.B1(n_338),
.B2(n_327),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_554),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_544),
.A2(n_406),
.B1(n_411),
.B2(n_396),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_344),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_537),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_528),
.A2(n_413),
.B1(n_424),
.B2(n_404),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_319),
.Y(n_621)
);

AO22x2_ASAP7_75t_L g622 ( 
.A1(n_542),
.A2(n_347),
.B1(n_354),
.B2(n_346),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_560),
.B(n_362),
.Y(n_623)
);

BUFx6f_ASAP7_75t_SL g624 ( 
.A(n_523),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g625 ( 
.A1(n_514),
.A2(n_433),
.B1(n_440),
.B2(n_439),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_537),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_547),
.A2(n_375),
.B1(n_377),
.B2(n_367),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_536),
.A2(n_453),
.B1(n_455),
.B2(n_441),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_595),
.B(n_321),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_579),
.B(n_323),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_591),
.A2(n_420),
.B1(n_466),
.B2(n_461),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_538),
.B(n_379),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_607),
.B(n_386),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_593),
.A2(n_483),
.B1(n_484),
.B2(n_476),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_527),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_512),
.A2(n_487),
.B1(n_489),
.B2(n_486),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_581),
.A2(n_503),
.B1(n_504),
.B2(n_494),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_566),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_579),
.B(n_325),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_594),
.A2(n_330),
.B1(n_334),
.B2(n_326),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_584),
.A2(n_337),
.B1(n_343),
.B2(n_335),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_602),
.A2(n_395),
.B1(n_398),
.B2(n_391),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_539),
.A2(n_349),
.B1(n_350),
.B2(n_348),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_548),
.A2(n_358),
.B1(n_360),
.B2(n_353),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_520),
.A2(n_408),
.B1(n_409),
.B2(n_407),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_520),
.A2(n_429),
.B1(n_430),
.B2(n_416),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_568),
.B(n_22),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_516),
.A2(n_515),
.B1(n_590),
.B2(n_583),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_547),
.A2(n_442),
.B1(n_449),
.B2(n_434),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_579),
.B(n_368),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_533),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_573),
.A2(n_370),
.B1(n_372),
.B2(n_369),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_555),
.A2(n_383),
.B1(n_385),
.B2(n_381),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_551),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_607),
.B(n_457),
.Y(n_656)
);

AO22x2_ASAP7_75t_L g657 ( 
.A1(n_553),
.A2(n_478),
.B1(n_479),
.B2(n_465),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_589),
.B(n_387),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_582),
.A2(n_400),
.B1(n_402),
.B2(n_397),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_602),
.A2(n_485),
.B1(n_499),
.B2(n_482),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_521),
.A2(n_510),
.B1(n_511),
.B2(n_501),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_553),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_551),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_540),
.B(n_403),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_589),
.B(n_600),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g668 ( 
.A(n_587),
.B(n_23),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_524),
.A2(n_410),
.B1(n_412),
.B2(n_405),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_589),
.B(n_417),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_545),
.B(n_418),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_551),
.Y(n_672)
);

AND2x2_ASAP7_75t_SL g673 ( 
.A(n_552),
.B(n_26),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_600),
.B(n_421),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_571),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_600),
.B(n_422),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_556),
.A2(n_428),
.B1(n_431),
.B2(n_425),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_557),
.A2(n_436),
.B1(n_438),
.B2(n_432),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_559),
.A2(n_450),
.B1(n_451),
.B2(n_444),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_603),
.B(n_26),
.Y(n_680)
);

OAI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_521),
.A2(n_458),
.B1(n_459),
.B2(n_452),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_564),
.A2(n_467),
.B1(n_471),
.B2(n_463),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_546),
.A2(n_473),
.B1(n_480),
.B2(n_472),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_561),
.A2(n_490),
.B1(n_491),
.B2(n_488),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_572),
.B(n_493),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_SL g686 ( 
.A1(n_565),
.A2(n_497),
.B1(n_498),
.B2(n_496),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_596),
.A2(n_506),
.B1(n_508),
.B2(n_502),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_599),
.A2(n_30),
.B1(n_27),
.B2(n_28),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_614),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_619),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_655),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_611),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_639),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_617),
.B(n_649),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_639),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_610),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_616),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_665),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_613),
.B(n_601),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_621),
.B(n_601),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_667),
.B(n_609),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_666),
.A2(n_549),
.B(n_532),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_629),
.B(n_609),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_656),
.B(n_585),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_665),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_631),
.B(n_586),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_640),
.B(n_585),
.Y(n_710)
);

INVxp33_ASAP7_75t_L g711 ( 
.A(n_625),
.Y(n_711)
);

XOR2xp5_ASAP7_75t_L g712 ( 
.A(n_653),
.B(n_684),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_658),
.Y(n_713)
);

XNOR2x2_ASAP7_75t_L g714 ( 
.A(n_664),
.B(n_599),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_675),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_659),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_672),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_672),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_623),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_634),
.B(n_609),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_648),
.Y(n_722)
);

XNOR2xp5_ASAP7_75t_SL g723 ( 
.A(n_668),
.B(n_541),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_685),
.Y(n_724)
);

XOR2xp5_ASAP7_75t_L g725 ( 
.A(n_612),
.B(n_83),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_673),
.B(n_603),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_622),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_660),
.B(n_571),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_622),
.Y(n_729)
);

BUFx8_ASAP7_75t_L g730 ( 
.A(n_652),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_636),
.B(n_574),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_632),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_641),
.B(n_513),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_627),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_627),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_650),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_651),
.B(n_608),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_650),
.Y(n_738)
);

XNOR2xp5_ASAP7_75t_L g739 ( 
.A(n_681),
.B(n_27),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_635),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_657),
.Y(n_741)
);

INVxp33_ASAP7_75t_L g742 ( 
.A(n_637),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_671),
.B(n_535),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_657),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_674),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_643),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_676),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_662),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_664),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_680),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_638),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_642),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_615),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_680),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_677),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_615),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_688),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_SL g758 ( 
.A(n_628),
.B(n_530),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_654),
.B(n_606),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_670),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_678),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_668),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_679),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_SL g764 ( 
.A(n_669),
.B(n_576),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_661),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_646),
.B(n_567),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_644),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_645),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_663),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_687),
.B(n_513),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_620),
.B(n_597),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_745),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_695),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_697),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_719),
.B(n_720),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_737),
.B(n_549),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_713),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_726),
.B(n_550),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_743),
.B(n_683),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_726),
.B(n_550),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_742),
.B(n_686),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_701),
.B(n_569),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_731),
.B(n_569),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_700),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_743),
.B(n_576),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_716),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_757),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_773),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_698),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_759),
.B(n_575),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_699),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_770),
.B(n_578),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_740),
.B(n_633),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_771),
.B(n_578),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_706),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_727),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_747),
.B(n_576),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_707),
.B(n_577),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_757),
.B(n_709),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_709),
.Y(n_802)
);

BUFx12f_ASAP7_75t_L g803 ( 
.A(n_730),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_715),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_741),
.B(n_84),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_707),
.B(n_577),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_710),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_742),
.B(n_633),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_R g809 ( 
.A(n_729),
.B(n_577),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_690),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_691),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_705),
.B(n_597),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_L g813 ( 
.A1(n_704),
.A2(n_519),
.B(n_513),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_763),
.B(n_597),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_689),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_734),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_744),
.B(n_85),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_704),
.B(n_598),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_735),
.B(n_736),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_708),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_692),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_722),
.B(n_598),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_760),
.B(n_87),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_767),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_710),
.Y(n_826)
);

NAND2x1p5_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_580),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_707),
.B(n_580),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_769),
.B(n_598),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_693),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_755),
.B(n_88),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_750),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_761),
.B(n_604),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_766),
.B(n_604),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_710),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_732),
.B(n_604),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_724),
.Y(n_837)
);

AND2x2_ASAP7_75t_SL g838 ( 
.A(n_749),
.B(n_605),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_740),
.B(n_605),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_710),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_765),
.B(n_605),
.Y(n_841)
);

AND2x4_ASAP7_75t_L g842 ( 
.A(n_733),
.B(n_89),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_710),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_756),
.B(n_580),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_746),
.B(n_588),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_717),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_707),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_754),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_707),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_772),
.B(n_91),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_748),
.B(n_588),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_702),
.B(n_588),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_702),
.B(n_592),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_728),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_753),
.B(n_592),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_753),
.B(n_517),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_764),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_718),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_721),
.B(n_519),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_728),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_703),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_714),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_739),
.Y(n_863)
);

OR2x2_ASAP7_75t_SL g864 ( 
.A(n_696),
.B(n_30),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_751),
.B(n_517),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_712),
.A2(n_529),
.B(n_517),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_822),
.B(n_751),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_777),
.B(n_711),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_789),
.B(n_790),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_775),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_775),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_822),
.B(n_758),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_774),
.B(n_846),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_845),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_774),
.B(n_768),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_801),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_779),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_789),
.B(n_839),
.Y(n_878)
);

CKINVDCx8_ASAP7_75t_R g879 ( 
.A(n_815),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_825),
.B(n_758),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_818),
.B(n_752),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_776),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_839),
.B(n_762),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_774),
.B(n_529),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_779),
.Y(n_885)
);

BUFx8_ASAP7_75t_L g886 ( 
.A(n_803),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_774),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_785),
.B(n_762),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_774),
.B(n_694),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_836),
.B(n_519),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_835),
.B(n_529),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_776),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_803),
.B(n_723),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_793),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_785),
.B(n_725),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_807),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_798),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_SL g898 ( 
.A(n_849),
.B(n_730),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_855),
.B(n_31),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_788),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_855),
.B(n_31),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_802),
.B(n_786),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_788),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_807),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_825),
.B(n_531),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_797),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_786),
.B(n_531),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_845),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_815),
.Y(n_909)
);

OR2x6_ASAP7_75t_L g910 ( 
.A(n_820),
.B(n_531),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_836),
.B(n_522),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_802),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_807),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_807),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_793),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_865),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_820),
.B(n_32),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_846),
.B(n_807),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_793),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_849),
.B(n_522),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_805),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_826),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_791),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_831),
.B(n_32),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_831),
.B(n_33),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_791),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_780),
.B(n_558),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_780),
.B(n_558),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_792),
.B(n_33),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_778),
.B(n_35),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_782),
.B(n_93),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_883),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_882),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_888),
.B(n_836),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_897),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_879),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_870),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_892),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_868),
.B(n_862),
.Y(n_940)
);

BUFx4f_ASAP7_75t_SL g941 ( 
.A(n_886),
.Y(n_941)
);

NAND2x1p5_ASAP7_75t_L g942 ( 
.A(n_921),
.B(n_849),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_887),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_867),
.B(n_782),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_889),
.Y(n_945)
);

INVx6_ASAP7_75t_SL g946 ( 
.A(n_893),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_867),
.B(n_778),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_871),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_876),
.B(n_781),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_889),
.Y(n_950)
);

NAND2x1p5_ASAP7_75t_L g951 ( 
.A(n_921),
.B(n_826),
.Y(n_951)
);

BUFx2_ASAP7_75t_SL g952 ( 
.A(n_873),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_887),
.Y(n_953)
);

BUFx5_ASAP7_75t_L g954 ( 
.A(n_894),
.Y(n_954)
);

INVx3_ASAP7_75t_SL g955 ( 
.A(n_909),
.Y(n_955)
);

INVx4_ASAP7_75t_L g956 ( 
.A(n_887),
.Y(n_956)
);

BUFx4f_ASAP7_75t_SL g957 ( 
.A(n_886),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_892),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_878),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_930),
.Y(n_960)
);

BUFx6f_ASAP7_75t_SL g961 ( 
.A(n_893),
.Y(n_961)
);

CKINVDCx14_ASAP7_75t_R g962 ( 
.A(n_895),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_896),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_875),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_873),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_896),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_875),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_896),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_923),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_907),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_904),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_874),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_907),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_904),
.Y(n_974)
);

BUFx2_ASAP7_75t_SL g975 ( 
.A(n_908),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_899),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_926),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_904),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_910),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_913),
.Y(n_980)
);

INVx6_ASAP7_75t_L g981 ( 
.A(n_910),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_877),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_917),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_885),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_916),
.B(n_784),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_913),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_913),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_944),
.A2(n_862),
.B1(n_925),
.B2(n_924),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_934),
.Y(n_989)
);

CKINVDCx11_ASAP7_75t_R g990 ( 
.A(n_955),
.Y(n_990)
);

CKINVDCx8_ASAP7_75t_R g991 ( 
.A(n_975),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_939),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_944),
.B(n_947),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_958),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_969),
.Y(n_995)
);

BUFx4_ASAP7_75t_SL g996 ( 
.A(n_937),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_960),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_940),
.B(n_881),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_977),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_950),
.B(n_819),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_943),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_959),
.Y(n_1002)
);

BUFx8_ASAP7_75t_SL g1003 ( 
.A(n_961),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_947),
.A2(n_925),
.B1(n_924),
.B2(n_872),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_955),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_936),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_982),
.Y(n_1007)
);

BUFx12f_ASAP7_75t_L g1008 ( 
.A(n_945),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_SL g1009 ( 
.A1(n_940),
.A2(n_808),
.B1(n_783),
.B2(n_863),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_941),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_961),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_935),
.A2(n_880),
.B1(n_872),
.B2(n_831),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_971),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_984),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_967),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_938),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_948),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_943),
.Y(n_1018)
);

BUFx12f_ASAP7_75t_L g1019 ( 
.A(n_933),
.Y(n_1019)
);

BUFx8_ASAP7_75t_L g1020 ( 
.A(n_964),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_985),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_949),
.A2(n_869),
.B(n_851),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_985),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_972),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_983),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_971),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_943),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_972),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_949),
.B(n_851),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_976),
.A2(n_962),
.B1(n_831),
.B2(n_857),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_941),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_981),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_976),
.A2(n_932),
.B1(n_914),
.B2(n_929),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_959),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_SL g1035 ( 
.A1(n_962),
.A2(n_863),
.B1(n_898),
.B2(n_858),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_957),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_978),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_965),
.A2(n_857),
.B1(n_824),
.B2(n_931),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_965),
.A2(n_824),
.B1(n_805),
.B2(n_817),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_963),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_978),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_988),
.A2(n_898),
.B1(n_864),
.B2(n_932),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_R g1043 ( 
.A(n_990),
.B(n_981),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_1026),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_1003),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1030),
.A2(n_795),
.B1(n_858),
.B2(n_890),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1009),
.A2(n_911),
.B1(n_901),
.B2(n_902),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_998),
.A2(n_824),
.B1(n_833),
.B2(n_829),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1004),
.A2(n_841),
.B1(n_834),
.B2(n_842),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_SL g1050 ( 
.A1(n_1035),
.A2(n_988),
.B(n_1004),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1012),
.A2(n_841),
.B1(n_842),
.B2(n_850),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_1039),
.A2(n_838),
.B1(n_914),
.B2(n_860),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1029),
.B(n_814),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1038),
.A2(n_838),
.B1(n_860),
.B2(n_952),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_1022),
.A2(n_814),
.B(n_823),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1022),
.A2(n_794),
.B1(n_796),
.B2(n_823),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_989),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1002),
.B(n_865),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_1034),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_1006),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1033),
.B(n_853),
.C(n_852),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1017),
.Y(n_1062)
);

AOI222xp33_ASAP7_75t_L g1063 ( 
.A1(n_1021),
.A2(n_864),
.B1(n_794),
.B2(n_796),
.C1(n_844),
.C2(n_856),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_SL g1064 ( 
.A1(n_991),
.A2(n_957),
.B1(n_1036),
.B2(n_1005),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_992),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_993),
.A2(n_850),
.B1(n_817),
.B2(n_805),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1023),
.B(n_856),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1024),
.B(n_844),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1008),
.A2(n_817),
.B1(n_805),
.B2(n_835),
.Y(n_1069)
);

OAI222xp33_ASAP7_75t_L g1070 ( 
.A1(n_994),
.A2(n_905),
.B1(n_928),
.B2(n_927),
.C1(n_894),
.C2(n_919),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_1028),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_1026),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1019),
.A2(n_843),
.B1(n_840),
.B2(n_799),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1000),
.A2(n_843),
.B1(n_840),
.B2(n_852),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_995),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_999),
.A2(n_838),
.B1(n_866),
.B2(n_813),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1000),
.A2(n_853),
.B1(n_812),
.B2(n_912),
.Y(n_1077)
);

OAI222xp33_ASAP7_75t_L g1078 ( 
.A1(n_1007),
.A2(n_905),
.B1(n_927),
.B2(n_928),
.C1(n_919),
.C2(n_915),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1014),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1016),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1037),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1015),
.B(n_819),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_SL g1083 ( 
.A1(n_1011),
.A2(n_866),
.B1(n_847),
.B2(n_826),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1041),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1040),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_SL g1086 ( 
.A(n_1020),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1032),
.A2(n_979),
.B1(n_970),
.B2(n_854),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_997),
.A2(n_903),
.B1(n_906),
.B2(n_900),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1025),
.A2(n_854),
.B1(n_973),
.B2(n_918),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1013),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_1013),
.B(n_956),
.Y(n_1091)
);

AOI211xp5_ASAP7_75t_L g1092 ( 
.A1(n_1010),
.A2(n_848),
.B(n_832),
.C(n_861),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1001),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_1001),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1031),
.A2(n_854),
.B1(n_827),
.B2(n_816),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1050),
.A2(n_830),
.B1(n_810),
.B2(n_821),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1058),
.B(n_1018),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1053),
.B(n_1063),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_SL g1099 ( 
.A1(n_1061),
.A2(n_828),
.B1(n_800),
.B2(n_806),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1047),
.A2(n_954),
.B1(n_971),
.B2(n_920),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1095),
.A2(n_1046),
.B1(n_1054),
.B2(n_1052),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1049),
.A2(n_811),
.B1(n_821),
.B2(n_810),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1055),
.A2(n_1048),
.B1(n_1056),
.B2(n_1051),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1067),
.B(n_787),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1059),
.A2(n_920),
.B1(n_946),
.B2(n_915),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1086),
.A2(n_1064),
.B1(n_1089),
.B2(n_1060),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1066),
.A2(n_804),
.B1(n_954),
.B2(n_1027),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_1092),
.A2(n_1073),
.B1(n_1069),
.B2(n_1059),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1076),
.A2(n_954),
.B1(n_1027),
.B2(n_891),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1074),
.A2(n_827),
.B1(n_951),
.B2(n_942),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1076),
.A2(n_1027),
.B1(n_891),
.B2(n_884),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1083),
.A2(n_1082),
.B(n_1087),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1077),
.A2(n_891),
.B1(n_859),
.B2(n_956),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1057),
.Y(n_1114)
);

OAI222xp33_ASAP7_75t_L g1115 ( 
.A1(n_1083),
.A2(n_951),
.B1(n_942),
.B2(n_974),
.C1(n_987),
.C2(n_986),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1071),
.A2(n_971),
.B1(n_922),
.B2(n_980),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1070),
.A2(n_922),
.B(n_974),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1068),
.B(n_1062),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1085),
.A2(n_1080),
.B1(n_1065),
.B2(n_1090),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1081),
.B(n_953),
.Y(n_1120)
);

NAND3xp33_ASAP7_75t_L g1121 ( 
.A(n_1071),
.B(n_966),
.C(n_963),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1079),
.B(n_819),
.Y(n_1122)
);

OAI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1075),
.A2(n_922),
.B1(n_968),
.B2(n_996),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_1044),
.A2(n_968),
.B1(n_809),
.B2(n_525),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1093),
.B(n_1084),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1088),
.A2(n_525),
.B1(n_526),
.B2(n_522),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1094),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1088),
.Y(n_1128)
);

OAI222xp33_ASAP7_75t_L g1129 ( 
.A1(n_1091),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_1129)
);

AOI222xp33_ASAP7_75t_L g1130 ( 
.A1(n_1043),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.C1(n_43),
.C2(n_44),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1072),
.A2(n_1045),
.B1(n_1078),
.B2(n_1070),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1042),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1042),
.A2(n_50),
.B1(n_46),
.B2(n_49),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1057),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1042),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1042),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_1042),
.B(n_57),
.C(n_58),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1042),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1042),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1042),
.A2(n_66),
.B(n_67),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1042),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1114),
.B(n_71),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1130),
.A2(n_72),
.B(n_73),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1132),
.A2(n_1135),
.B1(n_1136),
.B2(n_1133),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1118),
.B(n_72),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1134),
.B(n_73),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1125),
.B(n_76),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1097),
.B(n_77),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1128),
.B(n_77),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1123),
.B(n_1108),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1132),
.A2(n_1135),
.B1(n_1136),
.B2(n_1133),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1119),
.B(n_78),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1109),
.B(n_79),
.Y(n_1153)
);

OAI221xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1139),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_100),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_1117),
.A2(n_101),
.B(n_106),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1098),
.B(n_107),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1106),
.B(n_111),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1140),
.A2(n_1137),
.B1(n_1139),
.B2(n_1141),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1120),
.B(n_114),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1101),
.B(n_116),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1131),
.B(n_118),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1123),
.B(n_120),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1111),
.A2(n_121),
.B(n_123),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1104),
.B(n_124),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1105),
.B(n_126),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1127),
.B(n_129),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1103),
.B(n_1138),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1100),
.B(n_135),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1122),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1099),
.B(n_142),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1112),
.A2(n_147),
.B(n_151),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1105),
.B(n_154),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1096),
.B(n_159),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1143),
.B(n_1102),
.C(n_1121),
.Y(n_1174)
);

NAND4xp75_ASAP7_75t_L g1175 ( 
.A(n_1171),
.B(n_1129),
.C(n_1115),
.D(n_1124),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1169),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_L g1177 ( 
.A(n_1150),
.B(n_1113),
.C(n_1107),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1169),
.B(n_1116),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1154),
.B(n_1126),
.C(n_1110),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1158),
.B(n_167),
.C(n_170),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1169),
.B(n_171),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1142),
.Y(n_1182)
);

NAND4xp75_ASAP7_75t_L g1183 ( 
.A(n_1171),
.B(n_172),
.C(n_173),
.D(n_174),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1144),
.A2(n_175),
.B(n_176),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1148),
.B(n_177),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1151),
.B(n_179),
.C(n_183),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1156),
.B(n_184),
.C(n_186),
.Y(n_1187)
);

AO21x2_ASAP7_75t_L g1188 ( 
.A1(n_1172),
.A2(n_187),
.B(n_189),
.Y(n_1188)
);

NAND3xp33_ASAP7_75t_L g1189 ( 
.A(n_1160),
.B(n_191),
.C(n_192),
.Y(n_1189)
);

NAND4xp75_ASAP7_75t_L g1190 ( 
.A(n_1171),
.B(n_193),
.C(n_197),
.D(n_198),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1142),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1145),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_L g1193 ( 
.A(n_1160),
.B(n_201),
.C(n_205),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1146),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1148),
.B(n_207),
.Y(n_1195)
);

AND2x4_ASAP7_75t_SL g1196 ( 
.A(n_1159),
.B(n_208),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1147),
.B(n_211),
.Y(n_1197)
);

NAND3xp33_ASAP7_75t_L g1198 ( 
.A(n_1167),
.B(n_212),
.C(n_213),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1182),
.B(n_1147),
.Y(n_1199)
);

NAND4xp75_ASAP7_75t_L g1200 ( 
.A(n_1184),
.B(n_1171),
.C(n_1157),
.D(n_1165),
.Y(n_1200)
);

NAND4xp75_ASAP7_75t_L g1201 ( 
.A(n_1178),
.B(n_1162),
.C(n_1152),
.D(n_1170),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1176),
.Y(n_1202)
);

NAND4xp75_ASAP7_75t_L g1203 ( 
.A(n_1197),
.B(n_1152),
.C(n_1170),
.D(n_1161),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1191),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1194),
.B(n_1146),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1192),
.B(n_1149),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1185),
.B(n_1149),
.Y(n_1207)
);

NAND4xp75_ASAP7_75t_L g1208 ( 
.A(n_1175),
.B(n_1153),
.C(n_1163),
.D(n_1155),
.Y(n_1208)
);

AO22x2_ASAP7_75t_L g1209 ( 
.A1(n_1183),
.A2(n_1168),
.B1(n_1173),
.B2(n_1164),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_1190),
.Y(n_1210)
);

XOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1195),
.B(n_1159),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1188),
.B(n_1181),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1188),
.B(n_1155),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1174),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1196),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1198),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1193),
.B(n_1155),
.Y(n_1217)
);

XOR2x2_ASAP7_75t_L g1218 ( 
.A(n_1203),
.B(n_1189),
.Y(n_1218)
);

CKINVDCx16_ASAP7_75t_R g1219 ( 
.A(n_1206),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1212),
.Y(n_1220)
);

XNOR2x1_ASAP7_75t_L g1221 ( 
.A(n_1211),
.B(n_1177),
.Y(n_1221)
);

XOR2x2_ASAP7_75t_L g1222 ( 
.A(n_1201),
.B(n_1180),
.Y(n_1222)
);

INVxp67_ASAP7_75t_SL g1223 ( 
.A(n_1214),
.Y(n_1223)
);

NOR2x1_ASAP7_75t_L g1224 ( 
.A(n_1208),
.B(n_1217),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1202),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1202),
.Y(n_1226)
);

XNOR2x2_ASAP7_75t_L g1227 ( 
.A(n_1200),
.B(n_1209),
.Y(n_1227)
);

XOR2x2_ASAP7_75t_L g1228 ( 
.A(n_1207),
.B(n_1186),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1204),
.Y(n_1229)
);

OA22x2_ASAP7_75t_L g1230 ( 
.A1(n_1227),
.A2(n_1216),
.B1(n_1215),
.B2(n_1217),
.Y(n_1230)
);

AO22x2_ASAP7_75t_L g1231 ( 
.A1(n_1223),
.A2(n_1213),
.B1(n_1198),
.B2(n_1199),
.Y(n_1231)
);

AOI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1223),
.A2(n_1216),
.B1(n_1209),
.B2(n_1222),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_SL g1233 ( 
.A(n_1220),
.Y(n_1233)
);

XNOR2xp5_ASAP7_75t_L g1234 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1234)
);

OAI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1224),
.A2(n_1210),
.B1(n_1205),
.B2(n_1215),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1219),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1229),
.A2(n_1210),
.B1(n_1209),
.B2(n_1179),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1225),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1228),
.Y(n_1239)
);

XOR2x2_ASAP7_75t_L g1240 ( 
.A(n_1226),
.B(n_1187),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1236),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1233),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1238),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1237),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_1242),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1244),
.A2(n_1232),
.B1(n_1234),
.B2(n_1230),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1241),
.A2(n_1239),
.B1(n_1231),
.B2(n_1235),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1243),
.A2(n_1231),
.B1(n_1210),
.B2(n_1240),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1243),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1246),
.A2(n_1247),
.B1(n_1248),
.B2(n_1245),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1249),
.Y(n_1251)
);

NOR2x1_ASAP7_75t_L g1252 ( 
.A(n_1251),
.B(n_1166),
.Y(n_1252)
);

OA22x2_ASAP7_75t_L g1253 ( 
.A1(n_1250),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1253),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1252),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1255),
.Y(n_1256)
);

AOI211xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1254),
.A2(n_225),
.B(n_228),
.C(n_229),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1254),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1256),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1258),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1257),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1260),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1261),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_1263)
);

AO22x2_ASAP7_75t_L g1264 ( 
.A1(n_1259),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1262),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1264),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1263),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1266),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1265),
.A2(n_275),
.B(n_276),
.C(n_278),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1269),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_1268),
.B1(n_1270),
.B2(n_279),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1272),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1273),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.C(n_286),
.Y(n_1274)
);

AOI211xp5_ASAP7_75t_L g1275 ( 
.A1(n_1274),
.A2(n_287),
.B(n_288),
.C(n_289),
.Y(n_1275)
);


endmodule