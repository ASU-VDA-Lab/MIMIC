module fake_jpeg_28146_n_314 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_13),
.B1(n_14),
.B2(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_42),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_29),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_35),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_16),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_68),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_14),
.B1(n_17),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_69),
.B1(n_47),
.B2(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_26),
.C(n_27),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_27),
.C(n_61),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_47),
.B1(n_69),
.B2(n_40),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_26),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_77),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_36),
.B1(n_31),
.B2(n_32),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_82),
.B1(n_47),
.B2(n_65),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_26),
.B(n_32),
.C(n_28),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_100),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_68),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_110),
.B1(n_62),
.B2(n_31),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_30),
.C(n_34),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_58),
.Y(n_107)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_53),
.B1(n_17),
.B2(n_28),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_75),
.B(n_77),
.Y(n_125)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_27),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_70),
.B1(n_79),
.B2(n_83),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_115),
.B1(n_127),
.B2(n_132),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_82),
.B1(n_73),
.B2(n_77),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_74),
.B(n_82),
.C(n_71),
.Y(n_118)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_137),
.B(n_144),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_51),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_77),
.B1(n_87),
.B2(n_36),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_94),
.B(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_20),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_103),
.B(n_98),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_136),
.B(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_133),
.B1(n_97),
.B2(n_109),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_87),
.B1(n_62),
.B2(n_31),
.Y(n_132)
);

OAI22x1_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_25),
.B1(n_38),
.B2(n_30),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_51),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_81),
.B(n_64),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_57),
.A3(n_67),
.B1(n_66),
.B2(n_15),
.Y(n_137)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_22),
.B(n_18),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_141),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_15),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_143),
.C(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_86),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_108),
.B(n_51),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_153),
.B1(n_166),
.B2(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_92),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_72),
.B1(n_112),
.B2(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_108),
.Y(n_155)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_157),
.B(n_162),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_127),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_108),
.Y(n_159)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_67),
.B1(n_112),
.B2(n_57),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_174),
.B1(n_176),
.B2(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_92),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_169),
.B(n_171),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_46),
.B1(n_43),
.B2(n_67),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_92),
.C(n_34),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_170),
.C(n_140),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_93),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_34),
.C(n_51),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_117),
.A2(n_115),
.B1(n_137),
.B2(n_125),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_18),
.B(n_24),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_138),
.B(n_24),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_22),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_114),
.A2(n_43),
.B1(n_46),
.B2(n_18),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_169),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_123),
.C(n_136),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_185),
.C(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_134),
.C(n_135),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_190),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_134),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_203),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_166),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_132),
.B1(n_138),
.B2(n_139),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_196),
.B1(n_178),
.B2(n_147),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_144),
.C(n_131),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_170),
.C(n_164),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_43),
.B1(n_19),
.B2(n_24),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_145),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_10),
.C(n_11),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_175),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_10),
.B(n_11),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_202),
.A2(n_190),
.B(n_188),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_148),
.B(n_15),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_34),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_148),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_191),
.A2(n_172),
.B1(n_165),
.B2(n_162),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_227),
.B1(n_228),
.B2(n_202),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_152),
.B(n_164),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_222),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_180),
.B1(n_207),
.B2(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_230),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_161),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_157),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_174),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_45),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_192),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_243),
.B1(n_210),
.B2(n_209),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_185),
.C(n_186),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_241),
.C(n_222),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_194),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_181),
.C(n_183),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_206),
.B1(n_180),
.B2(n_203),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_218),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_224),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_25),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_237),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_216),
.B1(n_226),
.B2(n_217),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_265),
.B1(n_253),
.B2(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_252),
.C(n_262),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_205),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_232),
.A2(n_228),
.B1(n_223),
.B2(n_215),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_196),
.B1(n_227),
.B2(n_213),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_242),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_256),
.Y(n_270)
);

AO22x1_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_234),
.B1(n_243),
.B2(n_238),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_213),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_240),
.B(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_268),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_276),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_15),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_277),
.C(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_233),
.B1(n_23),
.B2(n_25),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_15),
.B1(n_16),
.B2(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_233),
.C(n_51),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_7),
.Y(n_280)
);

OR2x6_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_25),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g297 ( 
.A1(n_279),
.A2(n_5),
.A3(n_10),
.B1(n_8),
.B2(n_3),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_282),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_7),
.B(n_9),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_290),
.B(n_0),
.Y(n_292)
);

AOI31xp67_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_7),
.A3(n_9),
.B(n_11),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_287),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_0),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_15),
.C(n_6),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_278),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_15),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_5),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_292),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_269),
.C(n_6),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_298),
.B(n_4),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_299),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_300),
.B1(n_5),
.B2(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_4),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_290),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_293),
.A2(n_4),
.B(n_5),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_302),
.Y(n_307)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_304),
.C(n_298),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_305),
.A3(n_306),
.B1(n_291),
.B2(n_11),
.C1(n_2),
.C2(n_0),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_307),
.B(n_305),
.C(n_2),
.D(n_1),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_1),
.B(n_2),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_1),
.B(n_2),
.Y(n_314)
);


endmodule