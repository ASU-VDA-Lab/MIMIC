module fake_jpeg_10566_n_176 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_53),
.B1(n_52),
.B2(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_55),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_25),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_24),
.B1(n_28),
.B2(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_63),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_42),
.B1(n_14),
.B2(n_17),
.Y(n_78)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_78),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_53),
.B1(n_46),
.B2(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_79),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_39),
.B(n_51),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_38),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_62),
.C(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_41),
.C(n_50),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_106),
.C(n_84),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_102),
.B1(n_82),
.B2(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_13),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_41),
.C(n_44),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_117),
.Y(n_127)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_79),
.C(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_74),
.B1(n_78),
.B2(n_77),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_116),
.B1(n_100),
.B2(n_17),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_86),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_89),
.B1(n_82),
.B2(n_28),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22x1_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_90),
.B1(n_103),
.B2(n_96),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_95),
.B(n_98),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_41),
.C(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_41),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_120),
.A2(n_95),
.B1(n_102),
.B2(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_128),
.B1(n_27),
.B2(n_17),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_129),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_126),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_21),
.B(n_23),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_65),
.C(n_44),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_108),
.B1(n_111),
.B2(n_113),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_144),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_107),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

AO21x1_ASAP7_75t_SL g138 ( 
.A1(n_128),
.A2(n_115),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_131),
.B1(n_123),
.B2(n_130),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_145),
.B1(n_131),
.B2(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_85),
.B1(n_27),
.B2(n_58),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_150),
.B(n_154),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_127),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_153),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_139),
.B1(n_145),
.B2(n_126),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_156),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_139),
.B1(n_9),
.B2(n_10),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_12),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_8),
.A3(n_27),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_146),
.B(n_150),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_162),
.A2(n_156),
.B(n_155),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_165),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_160),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_165)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_157),
.B(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_168),
.B(n_163),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_3),
.B(n_5),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_174),
.B(n_23),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_58),
.B1(n_7),
.B2(n_6),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_23),
.Y(n_176)
);


endmodule