module fake_jpeg_13940_n_73 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx12_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_45)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_43),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_45),
.B1(n_2),
.B2(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_7),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_50),
.B1(n_23),
.B2(n_18),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_44),
.B1(n_39),
.B2(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_9),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_60),
.Y(n_66)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_10),
.CON(n_60),
.SN(n_60)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_22),
.B2(n_19),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_62),
.C(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_67),
.C(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_65),
.CI(n_20),
.CON(n_72),
.SN(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_16),
.Y(n_73)
);


endmodule