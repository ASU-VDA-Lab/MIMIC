module real_jpeg_21624_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_21),
.B1(n_22),
.B2(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_0),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_0),
.A2(n_1),
.B1(n_30),
.B2(n_79),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_24),
.B(n_35),
.C(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_1),
.A2(n_5),
.B1(n_35),
.B2(n_79),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_2),
.A2(n_26),
.B(n_31),
.Y(n_25)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_40),
.B(n_45),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_22),
.B(n_23),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_8),
.B(n_29),
.Y(n_104)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_20),
.B(n_79),
.C(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_7),
.B(n_79),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_53)
);

BUFx3_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_96),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_94),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_66),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_49),
.C(n_56),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_14),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_37),
.B2(n_38),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_25),
.B2(n_36),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_36),
.C(n_38),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_19),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_40),
.Y(n_42)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_22),
.A2(n_35),
.B(n_41),
.C(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_25),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_25),
.B(n_101),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_27),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_28),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_32),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_33),
.B(n_35),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_35),
.A2(n_45),
.B(n_52),
.C(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_35),
.B(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_35),
.B(n_43),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_36),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_39),
.B(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_49),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_49),
.B(n_73),
.C(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_49),
.A2(n_56),
.B1(n_57),
.B2(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_50),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_72),
.A2(n_73),
.B1(n_121),
.B2(n_125),
.Y(n_120)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2x1_ASAP7_75t_R g114 ( 
.A(n_73),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_115),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_93),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_92),
.B1(n_105),
.B2(n_109),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_105),
.C(n_130),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_133),
.B(n_137),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_127),
.B(n_132),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_118),
.B(n_126),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_110),
.B(n_117),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_105),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B(n_116),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);


endmodule