module fake_jpeg_25044_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_13),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_12),
.Y(n_49)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_17),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_23),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_17),
.B1(n_11),
.B2(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_25),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_50),
.B(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_49),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_18),
.B(n_14),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_28),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_1),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_28),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_25),
.C(n_26),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.C(n_25),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_50),
.B1(n_40),
.B2(n_52),
.C(n_41),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_74),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_46),
.B1(n_48),
.B2(n_45),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_72),
.B1(n_66),
.B2(n_75),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_58),
.C(n_60),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_43),
.C(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_76),
.B(n_66),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_61),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_62),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_1),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_85),
.A2(n_71),
.B(n_19),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_75),
.B1(n_59),
.B2(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_89),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_55),
.B(n_54),
.C(n_49),
.D(n_63),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_77),
.C(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_88),
.C(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_84),
.C(n_87),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_97),
.B(n_93),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_10),
.B(n_8),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_10),
.B(n_8),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_102),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);


endmodule