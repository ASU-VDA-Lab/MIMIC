module fake_jpeg_23855_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_18),
.B(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_21),
.Y(n_85)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_60),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_67),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_39),
.C(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_20),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_26),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_27),
.B1(n_19),
.B2(n_26),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_45),
.B1(n_40),
.B2(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_44),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_28),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_96),
.B1(n_50),
.B2(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_59),
.B(n_43),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_95),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_45),
.B1(n_38),
.B2(n_40),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_55),
.B(n_63),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_103),
.C(n_113),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_48),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_76),
.Y(n_132)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_72),
.B(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_122),
.B1(n_76),
.B2(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_116),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_50),
.B1(n_19),
.B2(n_49),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_68),
.C(n_46),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_1),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_92),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_50),
.B1(n_46),
.B2(n_52),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_89),
.C(n_71),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_128),
.Y(n_159)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_140),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_139),
.Y(n_170)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_135),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_96),
.B1(n_38),
.B2(n_40),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_137),
.B1(n_106),
.B2(n_110),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_25),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_74),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_25),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_147),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_101),
.B(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_115),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_81),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_78),
.C(n_70),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_113),
.C(n_103),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_154),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_167),
.B(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_122),
.C(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_109),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_71),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_172),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_115),
.B(n_106),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_133),
.Y(n_169)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_126),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_78),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_130),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_136),
.B1(n_148),
.B2(n_134),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_173),
.B1(n_91),
.B2(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_192),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_141),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_126),
.B1(n_139),
.B2(n_125),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_172),
.B1(n_154),
.B2(n_161),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_164),
.C(n_171),
.Y(n_212)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_201),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_70),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_165),
.B(n_160),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_155),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_169),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_202),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_158),
.B(n_124),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_203),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_211),
.B1(n_228),
.B2(n_200),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_168),
.B(n_151),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_227),
.C(n_198),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_215),
.B1(n_222),
.B2(n_200),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_166),
.B1(n_175),
.B2(n_119),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_32),
.B(n_18),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_226),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_119),
.B1(n_104),
.B2(n_105),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_178),
.B(n_184),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_105),
.C(n_94),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_180),
.B1(n_187),
.B2(n_185),
.Y(n_228)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_179),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_244),
.B1(n_216),
.B2(n_220),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_240),
.C(n_241),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_192),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_242),
.B1(n_246),
.B2(n_248),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_218),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_183),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_239),
.Y(n_272)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_212),
.C(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_247),
.C(n_216),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_191),
.C(n_181),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_202),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_229),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_234),
.B1(n_235),
.B2(n_242),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_199),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_44),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_267),
.C(n_268),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_217),
.B(n_205),
.C(n_213),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_244),
.B1(n_238),
.B2(n_230),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_206),
.B1(n_225),
.B2(n_219),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_263),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_94),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_31),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_271),
.B1(n_239),
.B2(n_33),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_54),
.C(n_83),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_54),
.C(n_83),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_88),
.C(n_44),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_31),
.C(n_33),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_88),
.B1(n_32),
.B2(n_17),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_285),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_28),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_1),
.B(n_2),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_282),
.B1(n_288),
.B2(n_255),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_259),
.A2(n_45),
.B1(n_40),
.B2(n_33),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_28),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_28),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_31),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_268),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_262),
.B(n_4),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_5),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_266),
.C(n_267),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_298),
.C(n_299),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_269),
.C(n_259),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_282),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_289),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_45),
.C(n_31),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_304),
.A2(n_29),
.B(n_22),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_308),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_275),
.B(n_287),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_311),
.B(n_313),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_303),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_293),
.B(n_5),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_315),
.Y(n_318)
);

AO221x1_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_29),
.B1(n_22),
.B2(n_8),
.C(n_9),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_295),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_300),
.C(n_302),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_6),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_7),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_322),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_321),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_297),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_312),
.B(n_305),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_29),
.C(n_22),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_11),
.C(n_12),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_327),
.B(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_319),
.C(n_318),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_11),
.C(n_13),
.Y(n_330)
);

INVx11_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_332),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_335),
.C(n_331),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_333),
.B(n_326),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_339),
.Y(n_340)
);

BUFx24_ASAP7_75t_SL g341 ( 
.A(n_340),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_13),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_14),
.C(n_326),
.Y(n_343)
);


endmodule