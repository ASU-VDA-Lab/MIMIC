module fake_netlist_5_1744_n_5454 (n_137, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_637, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_645, n_539, n_175, n_538, n_262, n_238, n_639, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_5454);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_639;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_5454;

wire n_924;
wire n_977;
wire n_2417;
wire n_2756;
wire n_2253;
wire n_4706;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_671;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_1107;
wire n_668;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_3188;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_2091;
wire n_1517;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_2032;
wire n_1566;
wire n_2587;
wire n_5406;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_882;
wire n_3156;
wire n_696;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_3653;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_2100;
wire n_5236;
wire n_3487;
wire n_3310;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_870;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_4790;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_727;
wire n_5210;
wire n_4967;
wire n_957;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_3200;
wire n_1664;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_4452;
wire n_4348;
wire n_5430;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_802;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_690;
wire n_4521;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_5322;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_5418;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_1661;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_1726;
wire n_3035;
wire n_5194;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_1109;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_687;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_5394;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5428;
wire n_3391;
wire n_4259;
wire n_2709;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_685;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2552;
wire n_2157;
wire n_1012;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_3114;
wire n_3125;
wire n_4981;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_695;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_1074;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_5401;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_666;
wire n_1433;
wire n_3152;
wire n_2256;
wire n_5106;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_667;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_951;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_4330;
wire n_3695;
wire n_2482;
wire n_2677;
wire n_3832;
wire n_3987;
wire n_902;
wire n_5352;
wire n_4991;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_5410;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_3638;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_4485;
wire n_4626;
wire n_1097;
wire n_1036;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_3089;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_663;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_858;
wire n_2985;
wire n_691;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_705;
wire n_3775;
wire n_4133;
wire n_678;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_677;
wire n_2723;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_906;
wire n_919;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_662;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5034;
wire n_1708;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_967;
wire n_2731;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_1283;
wire n_762;
wire n_5325;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_2646;
wire n_1605;
wire n_5173;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_984;
wire n_694;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4668;
wire n_4953;
wire n_3898;
wire n_849;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1998;
wire n_1019;
wire n_4686;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_1174;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_665;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_2003;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_5312;
wire n_985;
wire n_3404;
wire n_3217;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_676;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_672;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_898;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_5214;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2742;
wire n_2183;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_4171;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_3497;
wire n_1601;
wire n_5409;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_4636;
wire n_4584;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_3413;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_927;
wire n_2689;
wire n_3259;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_3261;
wire n_2200;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_688;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_864;
wire n_5420;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_947;
wire n_3710;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_897;
wire n_5280;
wire n_1428;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_680;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4912;
wire n_4813;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_857;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_2808;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_4491;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_689;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5216;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_765;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_701;
wire n_1023;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_842;
wire n_5434;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_5090;
wire n_1616;
wire n_4476;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_749;
wire n_5359;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_1506;
wire n_2867;
wire n_990;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_726;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1777;
wire n_1335;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1991;
wire n_2224;
wire n_1543;
wire n_732;
wire n_4743;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_5423;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_684;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_664;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_905;
wire n_5077;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_5314;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_682;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_4839;
wire n_5222;
wire n_1028;
wire n_4016;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_2027;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_1089;
wire n_5217;
wire n_1004;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_5396;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_2374;
wire n_1545;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_2761;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_976;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4472;
wire n_4462;
wire n_3433;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_2450;
wire n_3447;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_913;
wire n_3833;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_5426;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_1593;
wire n_3767;
wire n_2299;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5439;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_700;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_1366;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_3105;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_692;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_1188;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_5384;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_2619;
wire n_2444;
wire n_1110;
wire n_3123;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_866;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_693;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_679;
wire n_710;
wire n_3090;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_737;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_1225;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_2570;
wire n_1086;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_699;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_2823;
wire n_1076;
wire n_1408;
wire n_1761;
wire n_730;
wire n_5270;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_1032;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_14),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_365),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_170),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_461),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_660),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_201),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_572),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_134),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_419),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_437),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_55),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_186),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_10),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_50),
.Y(n_676)
);

CKINVDCx14_ASAP7_75t_R g677 ( 
.A(n_298),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_220),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_635),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_288),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_369),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_95),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_277),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_576),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_61),
.Y(n_685)
);

INVx4_ASAP7_75t_R g686 ( 
.A(n_511),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_185),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_403),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_646),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_219),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_81),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_19),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_317),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_227),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_350),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_135),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_105),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_268),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_389),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_247),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_410),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_594),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_99),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_23),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_260),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_25),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_506),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_17),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_161),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_395),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_415),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_293),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_137),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_286),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_497),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_442),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_467),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_583),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_283),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_189),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_554),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_91),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_615),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_304),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_224),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_561),
.Y(n_726)
);

BUFx10_ASAP7_75t_L g727 ( 
.A(n_547),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_463),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_327),
.Y(n_729)
);

INVxp33_ASAP7_75t_SL g730 ( 
.A(n_69),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_178),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_40),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_246),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_243),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_268),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_189),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_33),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_58),
.Y(n_738)
);

INVxp33_ASAP7_75t_R g739 ( 
.A(n_448),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_543),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_469),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_414),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_159),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_110),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_293),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_600),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_631),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_346),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_291),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_491),
.Y(n_750)
);

CKINVDCx14_ASAP7_75t_R g751 ( 
.A(n_249),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_36),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_632),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_137),
.Y(n_754)
);

INVxp67_ASAP7_75t_SL g755 ( 
.A(n_310),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_295),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_214),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_150),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_113),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_169),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_474),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_645),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_589),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_319),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_208),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_546),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_380),
.Y(n_767)
);

BUFx5_ASAP7_75t_L g768 ( 
.A(n_580),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_558),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_430),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_389),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_8),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_208),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_608),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_150),
.Y(n_775)
);

BUFx5_ASAP7_75t_L g776 ( 
.A(n_508),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_644),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_421),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_536),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_443),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_148),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_192),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_590),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_641),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_545),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_12),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_596),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_255),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_289),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_178),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_62),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_177),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_480),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_387),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_446),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_346),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_575),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_190),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_361),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_204),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_657),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_48),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_271),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_193),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_326),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_121),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_36),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_643),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_8),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_351),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_454),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_409),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_521),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_458),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_164),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_168),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_76),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_499),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_153),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_324),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_294),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_475),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_168),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_177),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_442),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_441),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_514),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_171),
.Y(n_828)
);

BUFx2_ASAP7_75t_R g829 ( 
.A(n_55),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_100),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_404),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_303),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_148),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_46),
.Y(n_834)
);

INVx1_ASAP7_75t_SL g835 ( 
.A(n_227),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_14),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_473),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_489),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_610),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_328),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_577),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_437),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_422),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_618),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_559),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_59),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_602),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_337),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_226),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_20),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_123),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_423),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_218),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_585),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_288),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_76),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_111),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_185),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_90),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_494),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_395),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_340),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_405),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_510),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_57),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_329),
.Y(n_866)
);

CKINVDCx14_ASAP7_75t_R g867 ( 
.A(n_119),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_599),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_478),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_298),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_257),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_13),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_250),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_249),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_254),
.Y(n_875)
);

CKINVDCx14_ASAP7_75t_R g876 ( 
.A(n_43),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_626),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_505),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_638),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_402),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_568),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_66),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_147),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_515),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_100),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_378),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_350),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_446),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_186),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_648),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_516),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_212),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_0),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_345),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_422),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_101),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_98),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_128),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_147),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_375),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_107),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_354),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_57),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_18),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_17),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_351),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_99),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_454),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_317),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_75),
.Y(n_910)
);

CKINVDCx14_ASAP7_75t_R g911 ( 
.A(n_465),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_352),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_407),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_5),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_108),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_11),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_281),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_604),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_280),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_358),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_344),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_209),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_544),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_367),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_485),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_556),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_477),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_513),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_560),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_340),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_232),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_138),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_367),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_176),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_650),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_654),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_309),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_541),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_258),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_83),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_241),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_54),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_292),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_37),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_214),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_518),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_301),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_58),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_564),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_134),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_539),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_282),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_31),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_218),
.Y(n_954)
);

CKINVDCx14_ASAP7_75t_R g955 ( 
.A(n_411),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_484),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_25),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_192),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_254),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_628),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_633),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_224),
.Y(n_962)
);

INVxp33_ASAP7_75t_L g963 ( 
.A(n_616),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_102),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_490),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_394),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_507),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_647),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_530),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_199),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_61),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_381),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_157),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_203),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_470),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_320),
.Y(n_976)
);

BUFx10_ASAP7_75t_L g977 ( 
.A(n_634),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_203),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_551),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_40),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_584),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_343),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_656),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_295),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_623),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_108),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_37),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_239),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_67),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_448),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_376),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_294),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_221),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_234),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_393),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_270),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_324),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_661),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_548),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_242),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_592),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_533),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_377),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_128),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_630),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_300),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_376),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_261),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_269),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_419),
.Y(n_1010)
);

BUFx2_ASAP7_75t_SL g1011 ( 
.A(n_571),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_144),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_342),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_443),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_603),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_436),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_321),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_562),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_11),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_420),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_252),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_614),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_496),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_391),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_323),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_282),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_459),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_659),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_582),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_244),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_79),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_127),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_210),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_375),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_26),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_269),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_451),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_239),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_88),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_15),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_204),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_362),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_382),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_609),
.Y(n_1044)
);

BUFx5_ASAP7_75t_L g1045 ( 
.A(n_410),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_233),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_323),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_161),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_458),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_597),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_38),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_481),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_574),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_512),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_336),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_49),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_49),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_290),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_86),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_651),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_310),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_620),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_302),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_427),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_257),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_217),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_283),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_135),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_260),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_105),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_371),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_483),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_35),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_194),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_273),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_605),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_453),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_456),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_549),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_466),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_215),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_64),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_343),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_397),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_465),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_428),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_495),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_476),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_39),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_451),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_611),
.Y(n_1091)
);

BUFx10_ASAP7_75t_L g1092 ( 
.A(n_424),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_217),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_470),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_175),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_42),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_542),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_237),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_82),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_405),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_207),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_69),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_333),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_285),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_251),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_306),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_540),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_624),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_355),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_223),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_527),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_4),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_487),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_359),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_118),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_103),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_595),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_374),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_364),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_432),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_5),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_4),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_407),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_152),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_353),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_325),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_115),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_235),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_334),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_348),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_416),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_336),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_180),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_297),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_408),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_438),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_612),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_87),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_409),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_467),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_393),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_92),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_235),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_50),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_52),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_464),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_685),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_851),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_851),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_851),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_851),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_851),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_851),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_851),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_851),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_677),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_851),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_995),
.B(n_0),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_669),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_733),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1045),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1045),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1045),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_733),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1045),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_881),
.B(n_1),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1045),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1045),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1045),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1045),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1045),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_689),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_662),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_689),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_718),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_718),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_685),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_723),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_723),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_862),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1146),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_747),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_751),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_867),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_747),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_813),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_665),
.Y(n_1188)
);

INVxp33_ASAP7_75t_SL g1189 ( 
.A(n_811),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_671),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_753),
.Y(n_1191)
);

INVxp33_ASAP7_75t_SL g1192 ( 
.A(n_930),
.Y(n_1192)
);

INVxp33_ASAP7_75t_SL g1193 ( 
.A(n_862),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_871),
.Y(n_1194)
);

INVxp33_ASAP7_75t_L g1195 ( 
.A(n_871),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_753),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_774),
.Y(n_1197)
);

INVx4_ASAP7_75t_R g1198 ( 
.A(n_938),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_876),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_774),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_777),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_881),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_777),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_793),
.Y(n_1204)
);

INVxp33_ASAP7_75t_SL g1205 ( 
.A(n_1035),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_793),
.Y(n_1206)
);

INVxp33_ASAP7_75t_SL g1207 ( 
.A(n_1035),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_818),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_818),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_911),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_827),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_827),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_844),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_844),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_682),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_685),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_847),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_847),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_860),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_676),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_860),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_955),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_864),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_864),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_891),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_685),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_891),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_929),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_903),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_903),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_929),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1075),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1075),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1122),
.Y(n_1234)
);

INVxp33_ASAP7_75t_SL g1235 ( 
.A(n_663),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_946),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_946),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_682),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_949),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1122),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_949),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_690),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_951),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_951),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_705),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_968),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_968),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_664),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1146),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_979),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_979),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_760),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_998),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_685),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_668),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_998),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_743),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_672),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1001),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1001),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_846),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_690),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1002),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_743),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_727),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_667),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1002),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1028),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1028),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1054),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1054),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1111),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1111),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_917),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1117),
.Y(n_1275)
);

CKINVDCx16_ASAP7_75t_R g1276 ( 
.A(n_673),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_727),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1117),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_724),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_691),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_724),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1072),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_724),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_883),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1146),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_883),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_915),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_915),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_948),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1146),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_932),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_948),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_980),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_743),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_980),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_743),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1126),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1126),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_667),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_743),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_796),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_796),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_973),
.Y(n_1303)
);

CKINVDCx16_ASAP7_75t_R g1304 ( 
.A(n_673),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_796),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_674),
.Y(n_1306)
);

INVxp33_ASAP7_75t_SL g1307 ( 
.A(n_675),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_987),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_796),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_667),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_796),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_997),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1014),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_815),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_667),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_815),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_815),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_678),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_815),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_673),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_815),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_842),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1069),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_842),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_842),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_681),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_842),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_683),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_727),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_842),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_889),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_1082),
.Y(n_1332)
);

XOR2x2_ASAP7_75t_L g1333 ( 
.A(n_739),
.B(n_730),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_687),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1089),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_889),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_889),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1119),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_889),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_889),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_688),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_916),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_916),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_692),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1146),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_916),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_916),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1131),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_694),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_916),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1021),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1021),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1021),
.Y(n_1353)
);

CKINVDCx16_ASAP7_75t_R g1354 ( 
.A(n_673),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_727),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_697),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1021),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_698),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1021),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1043),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_700),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_691),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_701),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_703),
.Y(n_1364)
);

INVxp33_ASAP7_75t_SL g1365 ( 
.A(n_708),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_977),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1043),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1043),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_695),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1043),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1043),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1103),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1103),
.Y(n_1373)
);

INVxp33_ASAP7_75t_L g1374 ( 
.A(n_695),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_977),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1103),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1103),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1103),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_699),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_699),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_706),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_706),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_768),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_717),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_717),
.Y(n_1385)
);

INVxp33_ASAP7_75t_L g1386 ( 
.A(n_737),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_737),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_711),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_742),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_768),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_742),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_754),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_754),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_767),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_963),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_767),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_770),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_770),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_772),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_667),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_772),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_709),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_775),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_775),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_778),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_778),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_789),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_789),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_790),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_790),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_794),
.Y(n_1411)
);

CKINVDCx16_ASAP7_75t_R g1412 ( 
.A(n_711),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_794),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_710),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_712),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_798),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_798),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_799),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_713),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_799),
.Y(n_1420)
);

BUFx6f_ASAP7_75t_L g1421 ( 
.A(n_1062),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_679),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_977),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_803),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_977),
.Y(n_1425)
);

CKINVDCx16_ASAP7_75t_R g1426 ( 
.A(n_711),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_768),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_679),
.Y(n_1428)
);

CKINVDCx16_ASAP7_75t_R g1429 ( 
.A(n_711),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_803),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_768),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_807),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_807),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1062),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_735),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_812),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_812),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_768),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1062),
.Y(n_1439)
);

INVxp33_ASAP7_75t_SL g1440 ( 
.A(n_716),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_814),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_814),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_823),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_823),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_830),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_719),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_830),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_833),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_720),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_833),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_722),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_728),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_768),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_840),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_840),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_768),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_848),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_750),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_848),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_849),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_849),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_729),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_852),
.Y(n_1463)
);

CKINVDCx16_ASAP7_75t_R g1464 ( 
.A(n_735),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_852),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1072),
.B(n_1),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_750),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_857),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_731),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_768),
.Y(n_1470)
);

CKINVDCx14_ASAP7_75t_R g1471 ( 
.A(n_666),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_857),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_865),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_865),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_885),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_776),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_761),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_761),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_885),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_887),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_784),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_887),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_732),
.Y(n_1483)
);

INVxp67_ASAP7_75t_SL g1484 ( 
.A(n_784),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_894),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_776),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_894),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_896),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_896),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_736),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_899),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_738),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_899),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_908),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_741),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_776),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_908),
.Y(n_1497)
);

INVxp33_ASAP7_75t_SL g1498 ( 
.A(n_744),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_910),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_910),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_912),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_912),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_921),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_921),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_924),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_924),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_745),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_941),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_941),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_959),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_959),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_748),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_981),
.B(n_2),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_693),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_749),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_993),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_993),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1009),
.Y(n_1518)
);

BUFx3_ASAP7_75t_L g1519 ( 
.A(n_981),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_752),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1009),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1079),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_776),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1024),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1024),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1025),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1025),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1027),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1079),
.B(n_2),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_756),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1027),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_758),
.Y(n_1532)
);

INVxp33_ASAP7_75t_SL g1533 ( 
.A(n_759),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1108),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1038),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_776),
.Y(n_1536)
);

INVxp33_ASAP7_75t_SL g1537 ( 
.A(n_764),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_704),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1038),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1040),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_776),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1040),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1041),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_765),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1041),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1062),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_771),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_773),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_776),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1047),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1047),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1049),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1108),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1049),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1062),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1059),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_781),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1059),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1068),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1068),
.Y(n_1560)
);

INVxp33_ASAP7_75t_SL g1561 ( 
.A(n_782),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1070),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_776),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1070),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1081),
.Y(n_1565)
);

INVx5_ASAP7_75t_L g1566 ( 
.A(n_1266),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1178),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1157),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1395),
.B(n_787),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1349),
.Y(n_1570)
);

BUFx8_ASAP7_75t_SL g1571 ( 
.A(n_1174),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1265),
.B(n_923),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1266),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1157),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1248),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1265),
.B(n_1277),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1174),
.Y(n_1577)
);

BUFx6f_ASAP7_75t_L g1578 ( 
.A(n_1266),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1216),
.Y(n_1579)
);

INVx5_ASAP7_75t_L g1580 ( 
.A(n_1266),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1328),
.B(n_735),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1266),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1178),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1299),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1419),
.B(n_735),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1512),
.B(n_1202),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1254),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1299),
.Y(n_1588)
);

INVx4_ASAP7_75t_L g1589 ( 
.A(n_1248),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_L g1590 ( 
.A(n_1277),
.B(n_1011),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1296),
.B(n_684),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1514),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1301),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1321),
.B(n_702),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1167),
.B(n_786),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1299),
.Y(n_1596)
);

INVx5_ASAP7_75t_L g1597 ( 
.A(n_1299),
.Y(n_1597)
);

BUFx12f_ASAP7_75t_L g1598 ( 
.A(n_1184),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1255),
.Y(n_1599)
);

INVx5_ASAP7_75t_L g1600 ( 
.A(n_1299),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1255),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1310),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1258),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1331),
.B(n_707),
.Y(n_1604)
);

BUFx12f_ASAP7_75t_L g1605 ( 
.A(n_1184),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1182),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1310),
.Y(n_1607)
);

BUFx8_ASAP7_75t_L g1608 ( 
.A(n_1165),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1343),
.B(n_1422),
.Y(n_1609)
);

INVx6_ASAP7_75t_L g1610 ( 
.A(n_1294),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1329),
.B(n_890),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1428),
.B(n_715),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1147),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1310),
.Y(n_1614)
);

BUFx12f_ASAP7_75t_L g1615 ( 
.A(n_1185),
.Y(n_1615)
);

INVx5_ASAP7_75t_L g1616 ( 
.A(n_1310),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1310),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1315),
.Y(n_1618)
);

BUFx8_ASAP7_75t_SL g1619 ( 
.A(n_1188),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1329),
.B(n_983),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1182),
.Y(n_1621)
);

INVx5_ASAP7_75t_L g1622 ( 
.A(n_1315),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_SL g1623 ( 
.A(n_1466),
.B(n_786),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1300),
.Y(n_1624)
);

INVx5_ASAP7_75t_L g1625 ( 
.A(n_1315),
.Y(n_1625)
);

INVx4_ASAP7_75t_L g1626 ( 
.A(n_1258),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1282),
.B(n_670),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1478),
.B(n_721),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1294),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1282),
.B(n_670),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1355),
.B(n_821),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1315),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1481),
.B(n_1484),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1226),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1538),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1294),
.Y(n_1636)
);

BUFx8_ASAP7_75t_SL g1637 ( 
.A(n_1188),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1355),
.B(n_786),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1306),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1240),
.Y(n_1640)
);

AND2x6_ASAP7_75t_L g1641 ( 
.A(n_1152),
.B(n_680),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1315),
.Y(n_1642)
);

INVx5_ASAP7_75t_L g1643 ( 
.A(n_1400),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1366),
.B(n_786),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1302),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1400),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1366),
.B(n_1092),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1400),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1148),
.Y(n_1649)
);

INVx5_ASAP7_75t_L g1650 ( 
.A(n_1400),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1229),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1160),
.B(n_821),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1400),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1421),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1421),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1185),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1421),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1147),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1187),
.B(n_855),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1226),
.Y(n_1660)
);

INVx5_ASAP7_75t_L g1661 ( 
.A(n_1421),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1189),
.B(n_855),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1305),
.Y(n_1663)
);

INVx5_ASAP7_75t_L g1664 ( 
.A(n_1421),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1229),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1434),
.Y(n_1666)
);

INVx5_ASAP7_75t_L g1667 ( 
.A(n_1434),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1199),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1189),
.B(n_874),
.Y(n_1669)
);

BUFx12f_ASAP7_75t_L g1670 ( 
.A(n_1199),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1306),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1148),
.B(n_726),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1309),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1434),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1349),
.Y(n_1675)
);

BUFx12f_ASAP7_75t_L g1676 ( 
.A(n_1210),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1314),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1148),
.B(n_740),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1375),
.B(n_1092),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1161),
.B(n_714),
.Y(n_1680)
);

BUFx12f_ASAP7_75t_L g1681 ( 
.A(n_1210),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1439),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1192),
.B(n_874),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1249),
.Y(n_1684)
);

CKINVDCx11_ASAP7_75t_R g1685 ( 
.A(n_1190),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1326),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1439),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1249),
.Y(n_1688)
);

AND2x6_ASAP7_75t_L g1689 ( 
.A(n_1152),
.B(n_680),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1375),
.B(n_1423),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1316),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1423),
.B(n_892),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1192),
.B(n_892),
.Y(n_1693)
);

BUFx12f_ASAP7_75t_L g1694 ( 
.A(n_1222),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1546),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1317),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1546),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1546),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1425),
.B(n_1092),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1257),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1326),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1425),
.B(n_696),
.Y(n_1702)
);

AND2x6_ASAP7_75t_L g1703 ( 
.A(n_1154),
.B(n_696),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1222),
.B(n_1092),
.Y(n_1704)
);

INVx3_ASAP7_75t_L g1705 ( 
.A(n_1546),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1319),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1320),
.B(n_725),
.Y(n_1707)
);

BUFx8_ASAP7_75t_SL g1708 ( 
.A(n_1190),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1230),
.Y(n_1709)
);

AND2x6_ASAP7_75t_L g1710 ( 
.A(n_1154),
.B(n_1149),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1320),
.B(n_725),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1546),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1555),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1322),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1235),
.B(n_1037),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1318),
.B(n_755),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1324),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1555),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1318),
.B(n_746),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1356),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1235),
.B(n_1057),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1414),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1284),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1307),
.B(n_1093),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1555),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1555),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1307),
.B(n_788),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1257),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1264),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1555),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1264),
.Y(n_1731)
);

INVx3_ASAP7_75t_L g1732 ( 
.A(n_1285),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1365),
.B(n_791),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1327),
.B(n_1330),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1285),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1290),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1414),
.B(n_802),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1336),
.B(n_763),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1365),
.B(n_792),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1290),
.Y(n_1740)
);

BUFx12f_ASAP7_75t_L g1741 ( 
.A(n_1230),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1311),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1232),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1311),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1337),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1339),
.B(n_1340),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1440),
.B(n_795),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1547),
.B(n_802),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1325),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1547),
.B(n_1279),
.Y(n_1750)
);

INVx5_ASAP7_75t_L g1751 ( 
.A(n_1325),
.Y(n_1751)
);

INVx5_ASAP7_75t_L g1752 ( 
.A(n_1345),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1342),
.B(n_769),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1334),
.B(n_779),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1346),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1440),
.B(n_800),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1356),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1281),
.B(n_843),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1159),
.B(n_1134),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1283),
.B(n_843),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1345),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1286),
.B(n_895),
.Y(n_1763)
);

INVx5_ASAP7_75t_L g1764 ( 
.A(n_1347),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1352),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1498),
.B(n_804),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1347),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1353),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1287),
.B(n_895),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1498),
.B(n_809),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1357),
.B(n_783),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_SL g1772 ( 
.A(n_1193),
.B(n_829),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1359),
.B(n_785),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1360),
.B(n_797),
.Y(n_1774)
);

BUFx8_ASAP7_75t_SL g1775 ( 
.A(n_1220),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1370),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1334),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1367),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1288),
.B(n_920),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1358),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1368),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1370),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1371),
.B(n_801),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1372),
.B(n_808),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1533),
.B(n_816),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_1373),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1289),
.B(n_920),
.Y(n_1787)
);

INVx5_ASAP7_75t_L g1788 ( 
.A(n_1458),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1458),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1193),
.B(n_734),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1376),
.B(n_822),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1377),
.Y(n_1792)
);

CKINVDCx6p67_ASAP7_75t_R g1793 ( 
.A(n_1276),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1378),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1467),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1467),
.Y(n_1796)
);

BUFx8_ASAP7_75t_SL g1797 ( 
.A(n_1220),
.Y(n_1797)
);

AND2x4_ASAP7_75t_L g1798 ( 
.A(n_1292),
.B(n_982),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1150),
.Y(n_1799)
);

INVxp33_ASAP7_75t_SL g1800 ( 
.A(n_1232),
.Y(n_1800)
);

BUFx3_ASAP7_75t_L g1801 ( 
.A(n_1293),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1477),
.Y(n_1802)
);

BUFx12f_ASAP7_75t_L g1803 ( 
.A(n_1233),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1533),
.B(n_817),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1477),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1519),
.B(n_837),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1519),
.B(n_838),
.Y(n_1807)
);

AND2x6_ASAP7_75t_L g1808 ( 
.A(n_1151),
.B(n_982),
.Y(n_1808)
);

BUFx8_ASAP7_75t_SL g1809 ( 
.A(n_1252),
.Y(n_1809)
);

BUFx12f_ASAP7_75t_L g1810 ( 
.A(n_1233),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1173),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1537),
.B(n_1561),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1522),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1295),
.B(n_1031),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1537),
.B(n_819),
.Y(n_1815)
);

NAND2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1522),
.B(n_757),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1534),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1534),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1175),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1553),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1553),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1153),
.B(n_839),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1379),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1155),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1156),
.B(n_845),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1380),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1358),
.Y(n_1827)
);

BUFx12f_ASAP7_75t_L g1828 ( 
.A(n_1234),
.Y(n_1828)
);

BUFx6f_ASAP7_75t_L g1829 ( 
.A(n_1381),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1382),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1341),
.B(n_854),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1341),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1561),
.B(n_825),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_L g1834 ( 
.A(n_1384),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1158),
.B(n_868),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1344),
.Y(n_1836)
);

BUFx8_ASAP7_75t_SL g1837 ( 
.A(n_1252),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1297),
.Y(n_1838)
);

INVx5_ASAP7_75t_L g1839 ( 
.A(n_1383),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1205),
.B(n_826),
.Y(n_1840)
);

HB1xp67_ASAP7_75t_L g1841 ( 
.A(n_1234),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1298),
.B(n_1031),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1344),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1205),
.B(n_828),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1361),
.Y(n_1845)
);

AND2x4_ASAP7_75t_L g1846 ( 
.A(n_1165),
.B(n_1061),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1207),
.B(n_831),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1181),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1385),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1361),
.B(n_869),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1363),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1162),
.B(n_877),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1163),
.B(n_878),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1207),
.B(n_832),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1164),
.B(n_879),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1194),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1176),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1166),
.B(n_884),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1194),
.B(n_1061),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1387),
.Y(n_1860)
);

INVx5_ASAP7_75t_L g1861 ( 
.A(n_1383),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1389),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1364),
.B(n_918),
.Y(n_1863)
);

BUFx12f_ASAP7_75t_L g1864 ( 
.A(n_1364),
.Y(n_1864)
);

INVx2_ASAP7_75t_SL g1865 ( 
.A(n_1402),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1215),
.B(n_1078),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1168),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_SL g1868 ( 
.A(n_1304),
.B(n_780),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1169),
.B(n_1170),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1171),
.B(n_1172),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1402),
.B(n_925),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1177),
.Y(n_1872)
);

AND2x6_ASAP7_75t_L g1873 ( 
.A(n_1390),
.B(n_1078),
.Y(n_1873)
);

BUFx8_ASAP7_75t_SL g1874 ( 
.A(n_1274),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1391),
.Y(n_1875)
);

BUFx8_ASAP7_75t_L g1876 ( 
.A(n_1179),
.Y(n_1876)
);

AND2x6_ASAP7_75t_L g1877 ( 
.A(n_1427),
.B(n_1109),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1513),
.B(n_820),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1363),
.Y(n_1879)
);

NOR2x1_ASAP7_75t_L g1880 ( 
.A(n_1180),
.B(n_1011),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1392),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1393),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1394),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1415),
.B(n_926),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1183),
.Y(n_1885)
);

BUFx8_ASAP7_75t_SL g1886 ( 
.A(n_1274),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1238),
.B(n_1109),
.Y(n_1887)
);

BUFx8_ASAP7_75t_SL g1888 ( 
.A(n_1303),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1415),
.B(n_927),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1186),
.B(n_928),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1242),
.B(n_1114),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1191),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1449),
.B(n_935),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1529),
.B(n_836),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1196),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1396),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1449),
.B(n_936),
.Y(n_1897)
);

AND2x6_ASAP7_75t_L g1898 ( 
.A(n_1427),
.B(n_1114),
.Y(n_1898)
);

BUFx8_ASAP7_75t_L g1899 ( 
.A(n_1197),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1262),
.B(n_1120),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1452),
.B(n_850),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1452),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1397),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1469),
.B(n_960),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1398),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1469),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1490),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1200),
.B(n_956),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1201),
.B(n_961),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1490),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1492),
.B(n_965),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1492),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1567),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1583),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1592),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1606),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1795),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1569),
.B(n_1471),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1592),
.B(n_1203),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1795),
.Y(n_1920)
);

BUFx6f_ASAP7_75t_L g1921 ( 
.A(n_1573),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1621),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1869),
.A2(n_1206),
.B(n_1204),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1569),
.B(n_1471),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1591),
.B(n_1594),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1635),
.Y(n_1926)
);

INVx6_ASAP7_75t_L g1927 ( 
.A(n_1788),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1795),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1634),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1813),
.B(n_1208),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1796),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1660),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1796),
.Y(n_1933)
);

INVx6_ASAP7_75t_L g1934 ( 
.A(n_1788),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1796),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1635),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1707),
.B(n_1209),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1684),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1840),
.A2(n_1308),
.B1(n_1312),
.B2(n_1303),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1802),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1802),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1813),
.B(n_1211),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1869),
.A2(n_1213),
.B(n_1212),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1680),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1707),
.B(n_1214),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1802),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1711),
.B(n_1217),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1805),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1591),
.B(n_1218),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1805),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1688),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1594),
.B(n_1219),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1613),
.Y(n_1953)
);

INVxp67_ASAP7_75t_L g1954 ( 
.A(n_1901),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1805),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1573),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1817),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1700),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1901),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1840),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1611),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1822),
.A2(n_1438),
.B(n_1431),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1658),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1604),
.B(n_1221),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1817),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_1571),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1817),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1728),
.Y(n_1968)
);

AND2x6_ASAP7_75t_L g1969 ( 
.A(n_1590),
.B(n_1438),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1604),
.B(n_1223),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1711),
.B(n_1627),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1729),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1821),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1740),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1627),
.B(n_1224),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1821),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1821),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1811),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1573),
.Y(n_1979)
);

AND2x6_ASAP7_75t_L g1980 ( 
.A(n_1638),
.B(n_1453),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1578),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1640),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1611),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1819),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1857),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1609),
.B(n_1495),
.Y(n_1986)
);

OA21x2_ASAP7_75t_L g1987 ( 
.A1(n_1870),
.A2(n_1825),
.B(n_1822),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1872),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1824),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1742),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1824),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1617),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1818),
.B(n_1225),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1870),
.A2(n_1228),
.B(n_1227),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1744),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1578),
.Y(n_1996)
);

BUFx2_ASAP7_75t_L g1997 ( 
.A(n_1620),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1617),
.Y(n_1998)
);

INVx5_ASAP7_75t_L g1999 ( 
.A(n_1710),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1629),
.B(n_1231),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1629),
.B(n_1236),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1824),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1824),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1578),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1640),
.Y(n_2005)
);

INVx3_ASAP7_75t_L g2006 ( 
.A(n_1617),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1644),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1620),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1647),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_L g2010 ( 
.A(n_1641),
.B(n_776),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1885),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1617),
.Y(n_2012)
);

AND2x6_ASAP7_75t_L g2013 ( 
.A(n_1679),
.B(n_1453),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1844),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1584),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1892),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1895),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1630),
.B(n_1237),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1609),
.B(n_1495),
.Y(n_2019)
);

XNOR2xp5_ASAP7_75t_L g2020 ( 
.A(n_1577),
.B(n_1333),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1572),
.B(n_1520),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1723),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1801),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1838),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1649),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1572),
.B(n_1595),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1856),
.B(n_1245),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1584),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1649),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1595),
.B(n_1520),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1799),
.Y(n_2031)
);

INVx3_ASAP7_75t_L g2032 ( 
.A(n_1674),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1749),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1636),
.B(n_1239),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1630),
.B(n_1241),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1776),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1818),
.B(n_1243),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1571),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1867),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1579),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1636),
.B(n_1244),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_SL g2042 ( 
.A(n_1868),
.B(n_762),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1587),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1806),
.B(n_1246),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_1584),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1699),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1593),
.Y(n_2047)
);

BUFx3_ASAP7_75t_L g2048 ( 
.A(n_1820),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1823),
.Y(n_2049)
);

AND2x2_ASAP7_75t_SL g2050 ( 
.A(n_1790),
.B(n_1120),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1816),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1856),
.B(n_1261),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1823),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1820),
.B(n_1247),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1702),
.B(n_1250),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1588),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1823),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1794),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1806),
.B(n_1807),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1674),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1826),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1826),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1826),
.Y(n_2063)
);

BUFx8_ASAP7_75t_L g2064 ( 
.A(n_1570),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1731),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1588),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1731),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1816),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1702),
.B(n_1758),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1758),
.B(n_1251),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1829),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1829),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1731),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1829),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1735),
.Y(n_2075)
);

BUFx2_ASAP7_75t_L g2076 ( 
.A(n_1608),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1716),
.B(n_1253),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1588),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_1674),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_1651),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1735),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1761),
.B(n_1256),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_1735),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1830),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1830),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1602),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1762),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1830),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1807),
.B(n_1259),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1761),
.B(n_1260),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1576),
.B(n_1263),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1834),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1834),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1834),
.Y(n_2094)
);

BUFx2_ASAP7_75t_L g2095 ( 
.A(n_1608),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1849),
.Y(n_2096)
);

AND2x2_ASAP7_75t_SL g2097 ( 
.A(n_1790),
.B(n_1123),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1762),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1586),
.B(n_1267),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1762),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1623),
.B(n_1530),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1767),
.Y(n_2102)
);

HB1xp67_ASAP7_75t_L g2103 ( 
.A(n_1651),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1576),
.B(n_1268),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1849),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1849),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1825),
.B(n_1269),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1610),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_1844),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1767),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1767),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1860),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1602),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1860),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1835),
.B(n_1270),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1860),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1782),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1847),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1862),
.Y(n_2119)
);

AND2x6_ASAP7_75t_L g2120 ( 
.A(n_1878),
.B(n_1456),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1835),
.B(n_1271),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1782),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1862),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1862),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1602),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1875),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1607),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1852),
.B(n_1272),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1782),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1852),
.B(n_1853),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1853),
.B(n_1273),
.Y(n_2131)
);

AND2x2_ASAP7_75t_SL g2132 ( 
.A(n_1868),
.B(n_1878),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1631),
.B(n_1275),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1732),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1875),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1665),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1875),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1732),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1736),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1881),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1881),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1665),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1881),
.Y(n_2143)
);

BUFx8_ASAP7_75t_L g2144 ( 
.A(n_1675),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_1631),
.B(n_1278),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_1692),
.B(n_1362),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_1722),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1692),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1736),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1607),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1786),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1709),
.Y(n_2152)
);

HB1xp67_ASAP7_75t_L g2153 ( 
.A(n_1709),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1786),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1792),
.Y(n_2155)
);

NAND2xp33_ASAP7_75t_R g2156 ( 
.A(n_1599),
.B(n_1530),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1882),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1690),
.B(n_1399),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1792),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1624),
.Y(n_2160)
);

CKINVDCx8_ASAP7_75t_R g2161 ( 
.A(n_1720),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1645),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1663),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1882),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1882),
.Y(n_2165)
);

AND2x4_ASAP7_75t_L g2166 ( 
.A(n_1690),
.B(n_1401),
.Y(n_2166)
);

INVxp67_ASAP7_75t_L g2167 ( 
.A(n_1847),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_1607),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1763),
.B(n_1403),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1673),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1623),
.B(n_1532),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_1763),
.B(n_1404),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1652),
.B(n_1362),
.Y(n_2173)
);

XNOR2xp5_ASAP7_75t_L g2174 ( 
.A(n_1577),
.B(n_1333),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1883),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1614),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1677),
.Y(n_2177)
);

OAI22xp5_ASAP7_75t_SL g2178 ( 
.A1(n_1854),
.A2(n_1312),
.B1(n_1313),
.B2(n_1308),
.Y(n_2178)
);

OAI22xp5_ASAP7_75t_SL g2179 ( 
.A1(n_1854),
.A2(n_1323),
.B1(n_1332),
.B2(n_1313),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1883),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1883),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1896),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1896),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_1633),
.B(n_1612),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1896),
.Y(n_2185)
);

INVxp67_ASAP7_75t_L g2186 ( 
.A(n_1727),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1691),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1696),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1614),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_1652),
.B(n_1374),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1706),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1614),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1855),
.B(n_1532),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1855),
.B(n_1544),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1858),
.B(n_1612),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1714),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1717),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1769),
.B(n_1405),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1743),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1674),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1745),
.Y(n_2201)
);

CKINVDCx16_ASAP7_75t_R g2202 ( 
.A(n_1741),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1755),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1765),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1659),
.B(n_1374),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1768),
.Y(n_2206)
);

INVx5_ASAP7_75t_L g2207 ( 
.A(n_1710),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1778),
.Y(n_2208)
);

INVxp67_ASAP7_75t_L g2209 ( 
.A(n_1727),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1781),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1903),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1858),
.B(n_1544),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1618),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1618),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1618),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1905),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1632),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1632),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1659),
.B(n_1386),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1734),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1734),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1632),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1642),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1746),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1746),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1760),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1642),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1642),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1760),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1646),
.Y(n_2230)
);

NAND2xp33_ASAP7_75t_L g2231 ( 
.A(n_1641),
.B(n_1548),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1628),
.B(n_1548),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1646),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1705),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1646),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_1737),
.B(n_1386),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1648),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1705),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1712),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1648),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_1769),
.B(n_1406),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_1779),
.B(n_1407),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1648),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1712),
.Y(n_2244)
);

CKINVDCx11_ASAP7_75t_R g2245 ( 
.A(n_1685),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1710),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_1653),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1653),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1653),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1654),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1654),
.Y(n_2251)
);

NOR2x1_ASAP7_75t_L g2252 ( 
.A(n_1589),
.B(n_766),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1654),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_1779),
.B(n_1408),
.Y(n_2254)
);

BUFx6f_ASAP7_75t_L g2255 ( 
.A(n_1655),
.Y(n_2255)
);

INVx3_ASAP7_75t_L g2256 ( 
.A(n_1655),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1655),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1710),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_1657),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1710),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1657),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1657),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1641),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1666),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1666),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1641),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1628),
.B(n_967),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1641),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1666),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1682),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1689),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1682),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1787),
.B(n_1409),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1689),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1689),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_1682),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1687),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1689),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_1787),
.B(n_1410),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1689),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1737),
.B(n_1195),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1748),
.B(n_1195),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1703),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_1687),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1687),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1633),
.B(n_969),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1672),
.B(n_985),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1695),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1703),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1703),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1703),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_1798),
.B(n_1411),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1703),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1748),
.B(n_1413),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1873),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1695),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_1695),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1697),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1873),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1873),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_1750),
.B(n_1416),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1672),
.B(n_1005),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1678),
.B(n_1015),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1678),
.B(n_1018),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_1697),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1697),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_2048),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_1986),
.B(n_2019),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_2048),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2151),
.Y(n_2310)
);

CKINVDCx20_ASAP7_75t_R g2311 ( 
.A(n_1939),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1978),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2186),
.B(n_1800),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_2209),
.B(n_1639),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_1986),
.B(n_1910),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2184),
.B(n_1719),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2151),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2154),
.Y(n_2318)
);

INVx2_ASAP7_75t_SL g2319 ( 
.A(n_1915),
.Y(n_2319)
);

INVx2_ASAP7_75t_SL g2320 ( 
.A(n_1915),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1984),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_1985),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2154),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1988),
.Y(n_2324)
);

INVx5_ASAP7_75t_L g2325 ( 
.A(n_1999),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2019),
.B(n_2148),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2155),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2155),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2184),
.B(n_1894),
.Y(n_2329)
);

BUFx10_ASAP7_75t_L g2330 ( 
.A(n_2132),
.Y(n_2330)
);

BUFx10_ASAP7_75t_L g2331 ( 
.A(n_2132),
.Y(n_2331)
);

AND2x6_ASAP7_75t_L g2332 ( 
.A(n_2263),
.B(n_1581),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2159),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2159),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1913),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2148),
.B(n_1910),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1913),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1914),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_SL g2339 ( 
.A(n_2042),
.B(n_1864),
.Y(n_2339)
);

AOI21x1_ASAP7_75t_L g2340 ( 
.A1(n_2130),
.A2(n_1753),
.B(n_1738),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_1960),
.B(n_1671),
.Y(n_2341)
);

AOI21x1_ASAP7_75t_L g2342 ( 
.A1(n_1925),
.A2(n_1753),
.B(n_1738),
.Y(n_2342)
);

INVxp33_ASAP7_75t_L g2343 ( 
.A(n_1936),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2195),
.B(n_1894),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2014),
.B(n_1832),
.Y(n_2345)
);

INVx2_ASAP7_75t_SL g2346 ( 
.A(n_2236),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1914),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1916),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1916),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1922),
.Y(n_2350)
);

INVxp33_ASAP7_75t_SL g2351 ( 
.A(n_2178),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1922),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2109),
.B(n_1902),
.Y(n_2353)
);

INVx5_ASAP7_75t_L g2354 ( 
.A(n_1999),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2059),
.B(n_1754),
.Y(n_2355)
);

AO22x2_ASAP7_75t_L g2356 ( 
.A1(n_2101),
.A2(n_1704),
.B1(n_1722),
.B2(n_1846),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_1929),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1929),
.Y(n_2358)
);

INVxp67_ASAP7_75t_SL g2359 ( 
.A(n_1921),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_1932),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1932),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1938),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1938),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_1954),
.B(n_1589),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1951),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2220),
.B(n_1831),
.Y(n_2366)
);

OAI22xp33_ASAP7_75t_SL g2367 ( 
.A1(n_2026),
.A2(n_2171),
.B1(n_2101),
.B2(n_2030),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1951),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_1956),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2118),
.B(n_1626),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1958),
.Y(n_2371)
);

INVx2_ASAP7_75t_SL g2372 ( 
.A(n_2236),
.Y(n_2372)
);

AND3x2_ASAP7_75t_L g2373 ( 
.A(n_2076),
.B(n_1772),
.C(n_1757),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2221),
.B(n_1850),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_1944),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1958),
.Y(n_2376)
);

NAND2xp33_ASAP7_75t_SL g2377 ( 
.A(n_2026),
.B(n_841),
.Y(n_2377)
);

CKINVDCx6p67_ASAP7_75t_R g2378 ( 
.A(n_2245),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2245),
.Y(n_2379)
);

INVx4_ASAP7_75t_L g2380 ( 
.A(n_1999),
.Y(n_2380)
);

AO21x2_ASAP7_75t_L g2381 ( 
.A1(n_1962),
.A2(n_1773),
.B(n_1771),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1968),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1968),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1972),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_2167),
.B(n_1626),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1972),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_1959),
.B(n_2193),
.Y(n_2387)
);

CKINVDCx6p67_ASAP7_75t_R g2388 ( 
.A(n_2202),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2224),
.B(n_2225),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1974),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2173),
.B(n_1701),
.Y(n_2391)
);

INVx3_ASAP7_75t_L g2392 ( 
.A(n_2246),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1974),
.Y(n_2393)
);

NOR2x1p5_ASAP7_75t_L g2394 ( 
.A(n_2027),
.B(n_1793),
.Y(n_2394)
);

INVx4_ASAP7_75t_L g2395 ( 
.A(n_1999),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2226),
.B(n_1863),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2258),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1990),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1990),
.Y(n_2399)
);

OAI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2194),
.A2(n_2212),
.B1(n_2232),
.B2(n_1983),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_1961),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_1995),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2229),
.B(n_1871),
.Y(n_2403)
);

AND3x2_ASAP7_75t_L g2404 ( 
.A(n_2076),
.B(n_1772),
.C(n_1780),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2069),
.B(n_1750),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2120),
.B(n_1884),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1995),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2033),
.Y(n_2408)
);

AO21x2_ASAP7_75t_L g2409 ( 
.A1(n_1962),
.A2(n_1773),
.B(n_1771),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2120),
.B(n_1889),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_1956),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2033),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2120),
.B(n_1893),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2036),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_1918),
.B(n_1701),
.Y(n_2415)
);

BUFx3_ASAP7_75t_L g2416 ( 
.A(n_2108),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2036),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_1919),
.B(n_1585),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_2260),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2134),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_1919),
.B(n_1846),
.Y(n_2421)
);

INVx8_ASAP7_75t_L g2422 ( 
.A(n_1980),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2173),
.B(n_1777),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2134),
.Y(n_2424)
);

NOR2x1p5_ASAP7_75t_L g2425 ( 
.A(n_2027),
.B(n_1568),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2211),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2216),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1930),
.Y(n_2428)
);

INVx3_ASAP7_75t_L g2429 ( 
.A(n_2266),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2120),
.B(n_1904),
.Y(n_2430)
);

BUFx10_ASAP7_75t_L g2431 ( 
.A(n_2158),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1930),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2069),
.B(n_1859),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_1924),
.A2(n_1601),
.B1(n_1603),
.B2(n_1575),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1930),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2138),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2138),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_2190),
.B(n_1777),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1942),
.Y(n_2439)
);

INVx5_ASAP7_75t_L g2440 ( 
.A(n_1999),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2139),
.Y(n_2441)
);

INVx5_ASAP7_75t_L g2442 ( 
.A(n_2207),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2139),
.Y(n_2443)
);

INVx1_ASAP7_75t_SL g2444 ( 
.A(n_1944),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1966),
.Y(n_2445)
);

BUFx16f_ASAP7_75t_R g2446 ( 
.A(n_2064),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1942),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2149),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2120),
.B(n_1897),
.Y(n_2449)
);

AND2x6_ASAP7_75t_L g2450 ( 
.A(n_2268),
.B(n_1911),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2149),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_1923),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2190),
.B(n_1836),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1923),
.Y(n_2454)
);

NAND2xp33_ASAP7_75t_L g2455 ( 
.A(n_2120),
.B(n_1980),
.Y(n_2455)
);

AOI22xp33_ASAP7_75t_L g2456 ( 
.A1(n_2050),
.A2(n_1662),
.B1(n_1683),
.B2(n_1669),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1942),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2107),
.B(n_1774),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2115),
.B(n_1774),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_1926),
.B(n_1836),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_1923),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1943),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_1961),
.Y(n_2463)
);

CKINVDCx6p67_ASAP7_75t_R g2464 ( 
.A(n_2095),
.Y(n_2464)
);

AO21x2_ASAP7_75t_L g2465 ( 
.A1(n_2171),
.A2(n_1784),
.B(n_1783),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2121),
.B(n_1783),
.Y(n_2466)
);

INVx3_ASAP7_75t_L g2467 ( 
.A(n_2271),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2128),
.B(n_1784),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2131),
.B(n_1791),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1966),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_1943),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1943),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1993),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2146),
.B(n_1859),
.Y(n_2474)
);

AND3x2_ASAP7_75t_L g2475 ( 
.A(n_2095),
.B(n_1851),
.C(n_1827),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2205),
.B(n_1843),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1993),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2108),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_1993),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_1994),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2069),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2037),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_1983),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1994),
.Y(n_2484)
);

OAI22xp5_ASAP7_75t_L g2485 ( 
.A1(n_1971),
.A2(n_1845),
.B1(n_1865),
.B2(n_1686),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_1994),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2025),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_1949),
.B(n_1952),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_1956),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2205),
.B(n_1843),
.Y(n_2490)
);

INVx1_ASAP7_75t_SL g2491 ( 
.A(n_2052),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2058),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_1956),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2274),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2058),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2160),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1964),
.B(n_1791),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2219),
.B(n_1812),
.Y(n_2498)
);

BUFx3_ASAP7_75t_L g2499 ( 
.A(n_2158),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_2275),
.Y(n_2500)
);

BUFx3_ASAP7_75t_L g2501 ( 
.A(n_2158),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2160),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_1997),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2029),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2278),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2162),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2162),
.Y(n_2507)
);

INVx5_ASAP7_75t_L g2508 ( 
.A(n_2207),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2163),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2163),
.Y(n_2510)
);

AND3x2_ASAP7_75t_L g2511 ( 
.A(n_1997),
.B(n_2008),
.C(n_2051),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2170),
.Y(n_2512)
);

INVx6_ASAP7_75t_L g2513 ( 
.A(n_2207),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2219),
.B(n_1812),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2170),
.Y(n_2515)
);

INVx2_ASAP7_75t_SL g2516 ( 
.A(n_2008),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2146),
.B(n_1733),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_2030),
.B(n_1733),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2177),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2177),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_1971),
.B(n_1739),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2050),
.A2(n_1662),
.B1(n_1683),
.B2(n_1669),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2188),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2188),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1970),
.B(n_1890),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2097),
.B(n_1739),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2097),
.B(n_1747),
.Y(n_2527)
);

AO21x2_ASAP7_75t_L g2528 ( 
.A1(n_2287),
.A2(n_1908),
.B(n_1890),
.Y(n_2528)
);

INVx3_ASAP7_75t_L g2529 ( 
.A(n_2280),
.Y(n_2529)
);

AND3x2_ASAP7_75t_L g2530 ( 
.A(n_2068),
.B(n_1879),
.C(n_1841),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2191),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2191),
.Y(n_2532)
);

INVx4_ASAP7_75t_L g2533 ( 
.A(n_2207),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2197),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2197),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2201),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_2099),
.B(n_1747),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2077),
.B(n_1693),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_2099),
.B(n_1756),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2283),
.Y(n_2540)
);

AOI22xp5_ASAP7_75t_L g2541 ( 
.A1(n_2231),
.A2(n_1766),
.B1(n_1770),
.B2(n_1756),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2289),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2201),
.Y(n_2543)
);

NAND2xp33_ASAP7_75t_L g2544 ( 
.A(n_1980),
.B(n_1873),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2065),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2077),
.B(n_1975),
.Y(n_2546)
);

INVxp67_ASAP7_75t_SL g2547 ( 
.A(n_1921),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_L g2548 ( 
.A(n_1980),
.B(n_1873),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2044),
.B(n_1908),
.Y(n_2549)
);

INVx1_ASAP7_75t_SL g2550 ( 
.A(n_2052),
.Y(n_2550)
);

INVx4_ASAP7_75t_L g2551 ( 
.A(n_2207),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2089),
.B(n_2286),
.Y(n_2552)
);

AOI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2231),
.A2(n_1770),
.B1(n_1785),
.B2(n_1766),
.Y(n_2553)
);

NAND2xp33_ASAP7_75t_L g2554 ( 
.A(n_1980),
.B(n_1877),
.Y(n_2554)
);

INVx2_ASAP7_75t_SL g2555 ( 
.A(n_2091),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2091),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2065),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2067),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2091),
.B(n_1785),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2067),
.Y(n_2560)
);

INVx3_ASAP7_75t_L g2561 ( 
.A(n_2290),
.Y(n_2561)
);

BUFx3_ASAP7_75t_L g2562 ( 
.A(n_2166),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_1980),
.A2(n_1815),
.B1(n_1833),
.B2(n_1804),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2073),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2073),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2075),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_2104),
.B(n_1804),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2104),
.B(n_1815),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2075),
.Y(n_2569)
);

INVxp67_ASAP7_75t_SL g2570 ( 
.A(n_1921),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2081),
.Y(n_2571)
);

INVx2_ASAP7_75t_SL g2572 ( 
.A(n_2104),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2081),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2083),
.Y(n_2574)
);

INVx1_ASAP7_75t_SL g2575 ( 
.A(n_2147),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2166),
.B(n_1833),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2291),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2083),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2087),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2267),
.B(n_1909),
.Y(n_2580)
);

INVxp33_ASAP7_75t_L g2581 ( 
.A(n_1982),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_SL g2582 ( 
.A(n_2252),
.B(n_1906),
.Y(n_2582)
);

OAI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2007),
.A2(n_1721),
.B1(n_1724),
.B2(n_1715),
.Y(n_2583)
);

INVx2_ASAP7_75t_SL g2584 ( 
.A(n_2281),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2087),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2166),
.B(n_1715),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2098),
.Y(n_2587)
);

NOR2x1p5_ASAP7_75t_L g2588 ( 
.A(n_2038),
.B(n_1574),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2021),
.B(n_1907),
.Y(n_2589)
);

AOI22xp33_ASAP7_75t_L g2590 ( 
.A1(n_1987),
.A2(n_2013),
.B1(n_1945),
.B2(n_1947),
.Y(n_2590)
);

OR2x6_ASAP7_75t_L g2591 ( 
.A(n_2133),
.B(n_1803),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_1975),
.B(n_1693),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_L g2593 ( 
.A(n_1956),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2293),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2295),
.Y(n_2595)
);

BUFx10_ASAP7_75t_L g2596 ( 
.A(n_2038),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_1987),
.A2(n_1724),
.B1(n_1721),
.B2(n_1877),
.Y(n_2597)
);

BUFx6f_ASAP7_75t_L g2598 ( 
.A(n_1979),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2299),
.Y(n_2599)
);

OAI22xp33_ASAP7_75t_L g2600 ( 
.A1(n_2009),
.A2(n_1907),
.B1(n_1912),
.B2(n_1848),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2300),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2098),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2100),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2187),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2046),
.B(n_1912),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2196),
.Y(n_2606)
);

BUFx2_ASAP7_75t_L g2607 ( 
.A(n_2005),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2100),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2013),
.B(n_1987),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2011),
.Y(n_2610)
);

INVxp67_ASAP7_75t_SL g2611 ( 
.A(n_1921),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2102),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2203),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2016),
.Y(n_2614)
);

NAND2xp33_ASAP7_75t_SL g2615 ( 
.A(n_2018),
.B(n_999),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2102),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2281),
.B(n_1704),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2110),
.Y(n_2618)
);

NAND2xp33_ASAP7_75t_R g2619 ( 
.A(n_2147),
.B(n_1866),
.Y(n_2619)
);

BUFx3_ASAP7_75t_L g2620 ( 
.A(n_2017),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2204),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2110),
.Y(n_2622)
);

BUFx10_ASAP7_75t_L g2623 ( 
.A(n_1969),
.Y(n_2623)
);

NAND2xp33_ASAP7_75t_SL g2624 ( 
.A(n_2018),
.B(n_1023),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2035),
.B(n_1848),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_SL g2626 ( 
.A(n_2282),
.B(n_1354),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2206),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2013),
.B(n_1909),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2156),
.Y(n_2629)
);

NAND2xp33_ASAP7_75t_L g2630 ( 
.A(n_2013),
.B(n_1877),
.Y(n_2630)
);

INVx3_ASAP7_75t_L g2631 ( 
.A(n_2111),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2208),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2111),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2117),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2013),
.B(n_1880),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2210),
.Y(n_2636)
);

AOI22xp33_ASAP7_75t_L g2637 ( 
.A1(n_2013),
.A2(n_1877),
.B1(n_1898),
.B2(n_1808),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2282),
.B(n_1388),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2117),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2037),
.Y(n_2640)
);

BUFx4f_ASAP7_75t_L g2641 ( 
.A(n_1969),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2054),
.Y(n_2642)
);

BUFx2_ASAP7_75t_L g2643 ( 
.A(n_2080),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2122),
.Y(n_2644)
);

NAND2xp33_ASAP7_75t_SL g2645 ( 
.A(n_2035),
.B(n_2021),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2122),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2129),
.Y(n_2647)
);

NAND2xp33_ASAP7_75t_SL g2648 ( 
.A(n_2133),
.B(n_1446),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2129),
.Y(n_2649)
);

INVx8_ASAP7_75t_L g2650 ( 
.A(n_1969),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2054),
.Y(n_2651)
);

INVx2_ASAP7_75t_SL g2652 ( 
.A(n_2055),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2055),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2302),
.B(n_1788),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2303),
.B(n_1788),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2031),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2213),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2040),
.B(n_1446),
.Y(n_2658)
);

OR2x6_ASAP7_75t_L g2659 ( 
.A(n_2145),
.B(n_1810),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2039),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2043),
.B(n_1451),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2213),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2304),
.B(n_1789),
.Y(n_2663)
);

CKINVDCx6p67_ASAP7_75t_R g2664 ( 
.A(n_2103),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_2301),
.B(n_1412),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2214),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2047),
.B(n_1451),
.Y(n_2667)
);

NOR2x1p5_ASAP7_75t_L g2668 ( 
.A(n_2022),
.B(n_1598),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2301),
.B(n_1426),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2000),
.B(n_1789),
.Y(n_2670)
);

NAND2xp33_ASAP7_75t_L g2671 ( 
.A(n_1969),
.B(n_1877),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2214),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2215),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2234),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_1937),
.A2(n_1947),
.B1(n_1945),
.B2(n_2145),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2238),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_SL g2677 ( 
.A(n_1937),
.B(n_2070),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2001),
.B(n_1789),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2034),
.B(n_1789),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2215),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2218),
.Y(n_2681)
);

BUFx6f_ASAP7_75t_L g2682 ( 
.A(n_1979),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2041),
.B(n_1989),
.Y(n_2683)
);

BUFx6f_ASAP7_75t_L g2684 ( 
.A(n_1979),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2169),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2070),
.B(n_1429),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2070),
.B(n_1435),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_1991),
.B(n_1898),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2169),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2169),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2218),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2223),
.Y(n_2692)
);

INVx4_ASAP7_75t_L g2693 ( 
.A(n_1927),
.Y(n_2693)
);

BUFx2_ASAP7_75t_L g2694 ( 
.A(n_2136),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2223),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2294),
.B(n_1900),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2172),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2294),
.B(n_1900),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2172),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2230),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2023),
.B(n_1462),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2230),
.Y(n_2702)
);

AND3x2_ASAP7_75t_L g2703 ( 
.A(n_2142),
.B(n_1841),
.C(n_1743),
.Y(n_2703)
);

BUFx2_ASAP7_75t_L g2704 ( 
.A(n_2152),
.Y(n_2704)
);

BUFx3_ASAP7_75t_L g2705 ( 
.A(n_2024),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2235),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2239),
.A2(n_1483),
.B1(n_1507),
.B2(n_1462),
.Y(n_2707)
);

NOR2x1p5_ASAP7_75t_L g2708 ( 
.A(n_2172),
.B(n_1605),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2327),
.Y(n_2709)
);

AND2x4_ASAP7_75t_L g2710 ( 
.A(n_2433),
.B(n_2198),
.Y(n_2710)
);

CKINVDCx20_ASAP7_75t_R g2711 ( 
.A(n_2388),
.Y(n_2711)
);

XNOR2x2_ASAP7_75t_L g2712 ( 
.A(n_2308),
.B(n_2020),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_2388),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2609),
.A2(n_2010),
.B(n_2003),
.Y(n_2714)
);

INVx2_ASAP7_75t_SL g2715 ( 
.A(n_2319),
.Y(n_2715)
);

XOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2629),
.B(n_2020),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2420),
.Y(n_2717)
);

INVxp67_ASAP7_75t_L g2718 ( 
.A(n_2619),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2625),
.B(n_1291),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2327),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2328),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2328),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_SL g2723 ( 
.A(n_2518),
.B(n_2161),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2310),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2310),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2317),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2317),
.Y(n_2727)
);

CKINVDCx20_ASAP7_75t_R g2728 ( 
.A(n_2629),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2318),
.Y(n_2729)
);

INVx1_ASAP7_75t_SL g2730 ( 
.A(n_2375),
.Y(n_2730)
);

INVxp33_ASAP7_75t_L g2731 ( 
.A(n_2343),
.Y(n_2731)
);

CKINVDCx20_ASAP7_75t_R g2732 ( 
.A(n_2445),
.Y(n_2732)
);

XNOR2xp5_ASAP7_75t_L g2733 ( 
.A(n_2425),
.B(n_2174),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2318),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2625),
.B(n_1348),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2538),
.B(n_2153),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2329),
.B(n_1969),
.Y(n_2737)
);

XOR2xp5_ASAP7_75t_L g2738 ( 
.A(n_2445),
.B(n_2174),
.Y(n_2738)
);

XNOR2xp5_ASAP7_75t_L g2739 ( 
.A(n_2470),
.B(n_2179),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2323),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2433),
.B(n_2198),
.Y(n_2741)
);

NOR2xp67_ASAP7_75t_L g2742 ( 
.A(n_2460),
.B(n_1615),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2323),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2333),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2333),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2470),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2334),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2334),
.Y(n_2748)
);

XOR2xp5_ASAP7_75t_L g2749 ( 
.A(n_2379),
.B(n_1323),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2348),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2498),
.B(n_2199),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2348),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2358),
.Y(n_2753)
);

CKINVDCx16_ASAP7_75t_R g2754 ( 
.A(n_2339),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2378),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2538),
.B(n_1953),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2514),
.B(n_1963),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2358),
.Y(n_2758)
);

XOR2xp5_ASAP7_75t_L g2759 ( 
.A(n_2379),
.B(n_1332),
.Y(n_2759)
);

XOR2xp5_ASAP7_75t_L g2760 ( 
.A(n_2311),
.B(n_1335),
.Y(n_2760)
);

XNOR2xp5_ASAP7_75t_L g2761 ( 
.A(n_2708),
.B(n_1335),
.Y(n_2761)
);

XOR2xp5_ASAP7_75t_L g2762 ( 
.A(n_2311),
.B(n_1338),
.Y(n_2762)
);

NOR2xp33_ASAP7_75t_L g2763 ( 
.A(n_2387),
.B(n_1483),
.Y(n_2763)
);

INVx2_ASAP7_75t_SL g2764 ( 
.A(n_2319),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2344),
.B(n_1338),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2420),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2361),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2361),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2365),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2365),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2376),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2376),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_2378),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2546),
.B(n_2198),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2316),
.B(n_1507),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2382),
.Y(n_2776)
);

CKINVDCx14_ASAP7_75t_R g2777 ( 
.A(n_2596),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2382),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2384),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2488),
.B(n_1969),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2546),
.B(n_2241),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2424),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2384),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2386),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2592),
.B(n_2241),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2355),
.B(n_1515),
.Y(n_2786)
);

NAND2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2641),
.B(n_1917),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2386),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2424),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2592),
.B(n_2241),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2390),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2320),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2390),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2455),
.A2(n_2010),
.B(n_2002),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2393),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2393),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2407),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2407),
.Y(n_2798)
);

XOR2xp5_ASAP7_75t_L g2799 ( 
.A(n_2541),
.B(n_1515),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2491),
.B(n_1464),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_2320),
.Y(n_2801)
);

XOR2x2_ASAP7_75t_L g2802 ( 
.A(n_2351),
.B(n_1619),
.Y(n_2802)
);

INVxp33_ASAP7_75t_L g2803 ( 
.A(n_2581),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2412),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2550),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2307),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2418),
.B(n_2242),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2552),
.B(n_2082),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2389),
.B(n_1557),
.Y(n_2809)
);

CKINVDCx20_ASAP7_75t_R g2810 ( 
.A(n_2464),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2412),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2436),
.Y(n_2812)
);

XNOR2xp5_ASAP7_75t_L g2813 ( 
.A(n_2394),
.B(n_1557),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2418),
.B(n_2242),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2436),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2437),
.Y(n_2816)
);

INVx3_ASAP7_75t_R g2817 ( 
.A(n_2607),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2437),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2441),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2441),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2443),
.Y(n_2821)
);

XNOR2x2_ASAP7_75t_L g2822 ( 
.A(n_2589),
.B(n_739),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2443),
.Y(n_2823)
);

CKINVDCx20_ASAP7_75t_R g2824 ( 
.A(n_2464),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2448),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2448),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2451),
.Y(n_2827)
);

XNOR2x2_ASAP7_75t_L g2828 ( 
.A(n_2583),
.B(n_805),
.Y(n_2828)
);

AND2x6_ASAP7_75t_L g2829 ( 
.A(n_2452),
.B(n_2454),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2451),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2507),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2421),
.B(n_2242),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_2596),
.Y(n_2833)
);

AOI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2455),
.A2(n_2590),
.B(n_2410),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2507),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2509),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2509),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2515),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2515),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2523),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2523),
.Y(n_2841)
);

OR2x6_ASAP7_75t_L g2842 ( 
.A(n_2591),
.B(n_1828),
.Y(n_2842)
);

INVx4_ASAP7_75t_SL g2843 ( 
.A(n_2450),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2314),
.B(n_2161),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2524),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2341),
.B(n_1619),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2524),
.Y(n_2847)
);

INVxp33_ASAP7_75t_L g2848 ( 
.A(n_2607),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2421),
.B(n_2254),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2532),
.Y(n_2850)
);

INVx4_ASAP7_75t_SL g2851 ( 
.A(n_2450),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2532),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2474),
.B(n_2254),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2543),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2543),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2492),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2474),
.B(n_2254),
.Y(n_2857)
);

OAI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2452),
.A2(n_2090),
.B(n_2082),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2335),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2335),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2337),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2492),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2345),
.B(n_1637),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2406),
.A2(n_1861),
.B(n_1839),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2575),
.B(n_2273),
.Y(n_2865)
);

XOR2x2_ASAP7_75t_L g2866 ( 
.A(n_2351),
.B(n_1637),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2337),
.Y(n_2867)
);

INVxp33_ASAP7_75t_L g2868 ( 
.A(n_2643),
.Y(n_2868)
);

INVxp67_ASAP7_75t_SL g2869 ( 
.A(n_2369),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2353),
.B(n_1708),
.Y(n_2870)
);

AND2x2_ASAP7_75t_L g2871 ( 
.A(n_2463),
.B(n_2273),
.Y(n_2871)
);

INVxp67_ASAP7_75t_SL g2872 ( 
.A(n_2369),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_SL g2873 ( 
.A(n_2582),
.B(n_1656),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2366),
.B(n_1920),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2495),
.Y(n_2875)
);

INVxp33_ASAP7_75t_L g2876 ( 
.A(n_2643),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2525),
.B(n_2082),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2463),
.B(n_2292),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2495),
.Y(n_2879)
);

CKINVDCx5p33_ASAP7_75t_R g2880 ( 
.A(n_2596),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2483),
.B(n_2292),
.Y(n_2881)
);

XNOR2xp5_ASAP7_75t_L g2882 ( 
.A(n_2475),
.B(n_1708),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2591),
.Y(n_2883)
);

INVxp67_ASAP7_75t_SL g2884 ( 
.A(n_2369),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2338),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2496),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2496),
.Y(n_2887)
);

INVx4_ASAP7_75t_L g2888 ( 
.A(n_2307),
.Y(n_2888)
);

BUFx8_ASAP7_75t_L g2889 ( 
.A(n_2694),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2502),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2502),
.Y(n_2891)
);

INVx1_ASAP7_75t_SL g2892 ( 
.A(n_2444),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_2615),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2433),
.B(n_2273),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2506),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2374),
.B(n_1928),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2416),
.B(n_2279),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2307),
.Y(n_2898)
);

CKINVDCx16_ASAP7_75t_R g2899 ( 
.A(n_2591),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2396),
.B(n_1931),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2338),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2506),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_2307),
.Y(n_2903)
);

NOR2xp33_ASAP7_75t_SL g2904 ( 
.A(n_2641),
.B(n_1668),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2510),
.Y(n_2905)
);

INVx4_ASAP7_75t_SL g2906 ( 
.A(n_2450),
.Y(n_2906)
);

CKINVDCx20_ASAP7_75t_R g2907 ( 
.A(n_2615),
.Y(n_2907)
);

INVx2_ASAP7_75t_SL g2908 ( 
.A(n_2694),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2510),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2512),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2512),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2519),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2519),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2520),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2591),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2347),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2520),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2483),
.B(n_2516),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2531),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2516),
.B(n_2696),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2704),
.Y(n_2921)
);

INVxp33_ASAP7_75t_L g2922 ( 
.A(n_2704),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_SL g2923 ( 
.A(n_2659),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2531),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2534),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2534),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2347),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2416),
.B(n_2279),
.Y(n_2928)
);

NOR2x1_ASAP7_75t_L g2929 ( 
.A(n_2315),
.B(n_1933),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2403),
.B(n_1935),
.Y(n_2930)
);

CKINVDCx20_ASAP7_75t_R g2931 ( 
.A(n_2624),
.Y(n_2931)
);

XNOR2xp5_ASAP7_75t_L g2932 ( 
.A(n_2373),
.B(n_2404),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2535),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2659),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2535),
.Y(n_2935)
);

XOR2xp5_ASAP7_75t_L g2936 ( 
.A(n_2553),
.B(n_1775),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2536),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2549),
.B(n_2090),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2536),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2349),
.Y(n_2940)
);

INVxp33_ASAP7_75t_L g2941 ( 
.A(n_2701),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2349),
.Y(n_2942)
);

CKINVDCx5p33_ASAP7_75t_R g2943 ( 
.A(n_2659),
.Y(n_2943)
);

CKINVDCx20_ASAP7_75t_R g2944 ( 
.A(n_2624),
.Y(n_2944)
);

INVx4_ASAP7_75t_L g2945 ( 
.A(n_2307),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2350),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2350),
.Y(n_2947)
);

OAI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2454),
.A2(n_2090),
.B(n_2279),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2497),
.B(n_2292),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2352),
.Y(n_2950)
);

AND2x2_ASAP7_75t_L g2951 ( 
.A(n_2696),
.B(n_1866),
.Y(n_2951)
);

XOR2xp5_ASAP7_75t_L g2952 ( 
.A(n_2707),
.B(n_1775),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2352),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2401),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2458),
.B(n_1940),
.Y(n_2955)
);

XNOR2x2_ASAP7_75t_L g2956 ( 
.A(n_2356),
.B(n_806),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2357),
.Y(n_2957)
);

CKINVDCx20_ASAP7_75t_R g2958 ( 
.A(n_2648),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2478),
.B(n_1941),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2499),
.Y(n_2960)
);

OR2x6_ASAP7_75t_L g2961 ( 
.A(n_2659),
.B(n_1670),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2357),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2313),
.B(n_1946),
.Y(n_2963)
);

XOR2xp5_ASAP7_75t_L g2964 ( 
.A(n_2563),
.B(n_1797),
.Y(n_2964)
);

BUFx3_ASAP7_75t_L g2965 ( 
.A(n_2401),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2360),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2370),
.B(n_1797),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2360),
.Y(n_2968)
);

CKINVDCx16_ASAP7_75t_R g2969 ( 
.A(n_2648),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2362),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2459),
.B(n_1948),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2362),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2363),
.Y(n_2973)
);

BUFx3_ASAP7_75t_L g2974 ( 
.A(n_2503),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2521),
.B(n_1950),
.Y(n_2975)
);

BUFx8_ASAP7_75t_L g2976 ( 
.A(n_2503),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2698),
.B(n_1887),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2363),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2466),
.B(n_1955),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2368),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2698),
.B(n_1887),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2368),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2478),
.B(n_1957),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2371),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2499),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2371),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_2664),
.Y(n_2987)
);

NOR2xp67_ASAP7_75t_L g2988 ( 
.A(n_2658),
.B(n_1676),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2383),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2526),
.B(n_1965),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2346),
.B(n_1891),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2346),
.B(n_1891),
.Y(n_2992)
);

CKINVDCx20_ASAP7_75t_R g2993 ( 
.A(n_2664),
.Y(n_2993)
);

CKINVDCx20_ASAP7_75t_R g2994 ( 
.A(n_2377),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2383),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2527),
.B(n_1967),
.Y(n_2996)
);

CKINVDCx20_ASAP7_75t_R g2997 ( 
.A(n_2377),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2398),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2372),
.B(n_1759),
.Y(n_2999)
);

AND2x4_ASAP7_75t_L g3000 ( 
.A(n_2501),
.B(n_1973),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2398),
.Y(n_3001)
);

CKINVDCx20_ASAP7_75t_R g3002 ( 
.A(n_2645),
.Y(n_3002)
);

AND2x4_ASAP7_75t_L g3003 ( 
.A(n_2501),
.B(n_1976),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2399),
.Y(n_3004)
);

XOR2xp5_ASAP7_75t_L g3005 ( 
.A(n_2434),
.B(n_1809),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2399),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2402),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2402),
.Y(n_3008)
);

OR2x6_ASAP7_75t_L g3009 ( 
.A(n_2588),
.B(n_1681),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2372),
.B(n_1759),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2610),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2408),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2408),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2584),
.B(n_1694),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2414),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2414),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2413),
.A2(n_1861),
.B(n_1839),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2417),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2417),
.Y(n_3019)
);

XOR2xp5_ASAP7_75t_L g3020 ( 
.A(n_2485),
.B(n_2405),
.Y(n_3020)
);

INVxp33_ASAP7_75t_L g3021 ( 
.A(n_2626),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2577),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2577),
.Y(n_3023)
);

NOR2xp67_ASAP7_75t_L g3024 ( 
.A(n_2661),
.B(n_1977),
.Y(n_3024)
);

AND2x6_ASAP7_75t_L g3025 ( 
.A(n_2461),
.B(n_2235),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2545),
.Y(n_3026)
);

CKINVDCx20_ASAP7_75t_R g3027 ( 
.A(n_2645),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2595),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2595),
.Y(n_3029)
);

AND2x2_ASAP7_75t_L g3030 ( 
.A(n_2584),
.B(n_1798),
.Y(n_3030)
);

CKINVDCx20_ASAP7_75t_R g3031 ( 
.A(n_2517),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2562),
.B(n_2049),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2537),
.B(n_2053),
.Y(n_3033)
);

XOR2xp5_ASAP7_75t_L g3034 ( 
.A(n_2405),
.B(n_1809),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2405),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2599),
.Y(n_3036)
);

XOR2xp5_ASAP7_75t_L g3037 ( 
.A(n_2638),
.B(n_1837),
.Y(n_3037)
);

CKINVDCx14_ASAP7_75t_R g3038 ( 
.A(n_2667),
.Y(n_3038)
);

AOI21xp5_ASAP7_75t_L g3039 ( 
.A1(n_2430),
.A2(n_1861),
.B(n_1839),
.Y(n_3039)
);

CKINVDCx14_ASAP7_75t_R g3040 ( 
.A(n_2385),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2599),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2601),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2601),
.Y(n_3043)
);

CKINVDCx5p33_ASAP7_75t_R g3044 ( 
.A(n_2610),
.Y(n_3044)
);

XOR2xp5_ASAP7_75t_L g3045 ( 
.A(n_2356),
.B(n_1837),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2481),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2604),
.Y(n_3047)
);

XNOR2x2_ASAP7_75t_L g3048 ( 
.A(n_2356),
.B(n_810),
.Y(n_3048)
);

AOI21xp5_ASAP7_75t_L g3049 ( 
.A1(n_2449),
.A2(n_1861),
.B(n_1839),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2604),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2606),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2606),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2613),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2613),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2621),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2621),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2545),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2627),
.Y(n_3058)
);

INVx2_ASAP7_75t_SL g3059 ( 
.A(n_2614),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2627),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2557),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2632),
.Y(n_3062)
);

CKINVDCx5p33_ASAP7_75t_R g3063 ( 
.A(n_2614),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2632),
.Y(n_3064)
);

BUFx3_ASAP7_75t_L g3065 ( 
.A(n_2620),
.Y(n_3065)
);

BUFx2_ASAP7_75t_R g3066 ( 
.A(n_2446),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2636),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2636),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2312),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2321),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2322),
.Y(n_3071)
);

XOR2x2_ASAP7_75t_L g3072 ( 
.A(n_2456),
.B(n_1874),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2522),
.B(n_1814),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2400),
.B(n_1874),
.Y(n_3074)
);

BUFx8_ASAP7_75t_L g3075 ( 
.A(n_2652),
.Y(n_3075)
);

AND2x2_ASAP7_75t_SL g3076 ( 
.A(n_2641),
.B(n_1886),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2324),
.Y(n_3077)
);

INVx2_ASAP7_75t_SL g3078 ( 
.A(n_2620),
.Y(n_3078)
);

NOR2xp67_ASAP7_75t_L g3079 ( 
.A(n_2415),
.B(n_2580),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2539),
.B(n_1814),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2656),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2656),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2674),
.Y(n_3083)
);

INVx2_ASAP7_75t_SL g3084 ( 
.A(n_2705),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2674),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_2652),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2676),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2468),
.B(n_2057),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_2469),
.B(n_2391),
.Y(n_3089)
);

BUFx2_ASAP7_75t_L g3090 ( 
.A(n_2921),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_L g3091 ( 
.A1(n_2956),
.A2(n_2640),
.B1(n_2651),
.B2(n_2642),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_3079),
.B(n_2723),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_SL g3093 ( 
.A(n_2723),
.B(n_2367),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_SL g3094 ( 
.A(n_3089),
.B(n_2330),
.Y(n_3094)
);

NOR3xp33_ASAP7_75t_L g3095 ( 
.A(n_2763),
.B(n_2438),
.C(n_2423),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2717),
.Y(n_3096)
);

AOI22xp33_ASAP7_75t_L g3097 ( 
.A1(n_3048),
.A2(n_2828),
.B1(n_3089),
.B2(n_2763),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2877),
.B(n_2330),
.Y(n_3098)
);

AOI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2786),
.A2(n_2476),
.B1(n_2490),
.B2(n_2453),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2877),
.B(n_2640),
.Y(n_3100)
);

OR2x2_ASAP7_75t_L g3101 ( 
.A(n_2719),
.B(n_2653),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2938),
.B(n_2330),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2938),
.B(n_2642),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2965),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2709),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2949),
.B(n_2651),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2949),
.B(n_2482),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_2765),
.B(n_2331),
.Y(n_3108)
);

AOI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_2786),
.A2(n_2559),
.B1(n_2568),
.B2(n_2567),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2808),
.B(n_2326),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2720),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2941),
.B(n_2331),
.Y(n_3112)
);

AND2x4_ASAP7_75t_L g3113 ( 
.A(n_2832),
.B(n_2562),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2721),
.Y(n_3114)
);

INVx4_ASAP7_75t_L g3115 ( 
.A(n_2960),
.Y(n_3115)
);

O2A1O1Ixp33_ASAP7_75t_L g3116 ( 
.A1(n_2775),
.A2(n_2586),
.B(n_2617),
.C(n_2576),
.Y(n_3116)
);

INVx2_ASAP7_75t_SL g3117 ( 
.A(n_2974),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_2730),
.Y(n_3118)
);

AND2x4_ASAP7_75t_L g3119 ( 
.A(n_2849),
.B(n_2309),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2808),
.B(n_2597),
.Y(n_3120)
);

AOI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_3073),
.A2(n_2356),
.B1(n_2331),
.B2(n_2528),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_3088),
.B(n_2675),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_3088),
.B(n_2653),
.Y(n_3123)
);

OAI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2955),
.A2(n_2428),
.B1(n_2435),
.B2(n_2432),
.Y(n_3124)
);

BUFx3_ASAP7_75t_L g3125 ( 
.A(n_2889),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2766),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2955),
.B(n_2971),
.Y(n_3127)
);

NOR2xp67_ASAP7_75t_SL g3128 ( 
.A(n_2754),
.B(n_2309),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2971),
.B(n_2528),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2979),
.B(n_2528),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2809),
.B(n_2555),
.Y(n_3131)
);

INVx8_ASAP7_75t_L g3132 ( 
.A(n_2710),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2782),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2722),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2979),
.B(n_2555),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3047),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2874),
.B(n_2896),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_3050),
.Y(n_3138)
);

OAI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_2780),
.A2(n_2628),
.B1(n_2572),
.B2(n_2556),
.Y(n_3139)
);

NAND2xp33_ASAP7_75t_L g3140 ( 
.A(n_2960),
.B(n_2332),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2735),
.B(n_2605),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3051),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2789),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2874),
.B(n_2556),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2896),
.B(n_2572),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_L g3146 ( 
.A(n_2775),
.B(n_2600),
.Y(n_3146)
);

NAND2xp33_ASAP7_75t_L g3147 ( 
.A(n_2960),
.B(n_2332),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2900),
.B(n_2465),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2900),
.B(n_2465),
.Y(n_3149)
);

INVxp67_ASAP7_75t_L g3150 ( 
.A(n_2792),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2809),
.B(n_2364),
.Y(n_3151)
);

AOI22xp33_ASAP7_75t_L g3152 ( 
.A1(n_2785),
.A2(n_2332),
.B1(n_2465),
.B2(n_2462),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2736),
.B(n_2665),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2718),
.B(n_2669),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2806),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_3026),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2930),
.B(n_2439),
.Y(n_3157)
);

BUFx3_ASAP7_75t_L g3158 ( 
.A(n_2889),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2930),
.B(n_2447),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_3057),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2790),
.B(n_2457),
.Y(n_3161)
);

OAI22xp33_ASAP7_75t_L g3162 ( 
.A1(n_3052),
.A2(n_2473),
.B1(n_2479),
.B2(n_2477),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2756),
.B(n_2677),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_2799),
.A2(n_2332),
.B1(n_2462),
.B2(n_2461),
.Y(n_3164)
);

AOI22x1_ASAP7_75t_L g3165 ( 
.A1(n_2794),
.A2(n_2397),
.B1(n_2419),
.B2(n_2392),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3053),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3061),
.Y(n_3167)
);

INVx2_ASAP7_75t_SL g3168 ( 
.A(n_2908),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2718),
.B(n_2686),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2774),
.B(n_2332),
.Y(n_3170)
);

NAND2xp33_ASAP7_75t_SL g3171 ( 
.A(n_2817),
.B(n_2668),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3054),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2781),
.B(n_2332),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_3044),
.B(n_2431),
.Y(n_3174)
);

INVxp33_ASAP7_75t_SL g3175 ( 
.A(n_2746),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2963),
.B(n_2689),
.Y(n_3176)
);

OR2x2_ASAP7_75t_L g3177 ( 
.A(n_2730),
.B(n_2687),
.Y(n_3177)
);

AOI22xp5_ASAP7_75t_L g3178 ( 
.A1(n_3031),
.A2(n_2156),
.B1(n_2336),
.B2(n_2685),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2963),
.B(n_2697),
.Y(n_3179)
);

BUFx8_ASAP7_75t_L g3180 ( 
.A(n_2923),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3002),
.A2(n_2699),
.B1(n_2690),
.B2(n_2705),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3055),
.Y(n_3182)
);

NAND2xp33_ASAP7_75t_L g3183 ( 
.A(n_2985),
.B(n_2450),
.Y(n_3183)
);

INVx2_ASAP7_75t_SL g3184 ( 
.A(n_2892),
.Y(n_3184)
);

OAI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2737),
.A2(n_2340),
.B(n_2342),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_3063),
.B(n_2920),
.Y(n_3186)
);

INVx3_ASAP7_75t_L g3187 ( 
.A(n_2806),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3056),
.Y(n_3188)
);

INVx8_ASAP7_75t_L g3189 ( 
.A(n_2710),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2859),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_3058),
.B(n_2487),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3060),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2844),
.B(n_2340),
.Y(n_3193)
);

OR2x2_ASAP7_75t_SL g3194 ( 
.A(n_2969),
.B(n_1886),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2805),
.B(n_2487),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_SL g3196 ( 
.A(n_2985),
.B(n_2431),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2985),
.B(n_2431),
.Y(n_3197)
);

AOI22xp33_ASAP7_75t_L g3198 ( 
.A1(n_3027),
.A2(n_2471),
.B1(n_2480),
.B2(n_2472),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3062),
.B(n_3064),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_3067),
.B(n_2504),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2805),
.B(n_2504),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3068),
.B(n_2660),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2999),
.B(n_2660),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_SL g3204 ( 
.A(n_2918),
.B(n_2426),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3010),
.B(n_2807),
.Y(n_3205)
);

INVx2_ASAP7_75t_SL g3206 ( 
.A(n_2892),
.Y(n_3206)
);

AOI221xp5_ASAP7_75t_L g3207 ( 
.A1(n_3074),
.A2(n_1077),
.B1(n_824),
.B2(n_858),
.C(n_970),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2865),
.B(n_2951),
.Y(n_3208)
);

BUFx6f_ASAP7_75t_L g3209 ( 
.A(n_2806),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2814),
.B(n_2683),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2860),
.Y(n_3211)
);

AND2x6_ASAP7_75t_SL g3212 ( 
.A(n_3009),
.B(n_2846),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2975),
.B(n_2342),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_2871),
.B(n_2427),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_2975),
.B(n_2676),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2861),
.Y(n_3216)
);

NOR2xp33_ASAP7_75t_L g3217 ( 
.A(n_2751),
.B(n_2703),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2751),
.B(n_2511),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2977),
.B(n_2471),
.Y(n_3219)
);

O2A1O1Ixp5_ASAP7_75t_L g3220 ( 
.A1(n_2834),
.A2(n_2480),
.B(n_2484),
.C(n_2472),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2981),
.B(n_2484),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2848),
.B(n_2530),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_2878),
.B(n_2623),
.Y(n_3223)
);

BUFx3_ASAP7_75t_L g3224 ( 
.A(n_2976),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_2867),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_2732),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3033),
.B(n_2486),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2750),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2752),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2885),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3033),
.B(n_2486),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2853),
.B(n_2857),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3081),
.B(n_2557),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3082),
.B(n_2558),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2753),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2758),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2901),
.Y(n_3237)
);

BUFx4f_ASAP7_75t_L g3238 ( 
.A(n_2961),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2767),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2868),
.B(n_2392),
.Y(n_3240)
);

INVx1_ASAP7_75t_SL g3241 ( 
.A(n_2876),
.Y(n_3241)
);

INVxp67_ASAP7_75t_SL g3242 ( 
.A(n_2869),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_2780),
.B(n_2737),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_2994),
.A2(n_2635),
.B1(n_2450),
.B2(n_2061),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2997),
.A2(n_2450),
.B1(n_2062),
.B2(n_2071),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3083),
.B(n_2558),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2768),
.Y(n_3247)
);

INVx2_ASAP7_75t_SL g3248 ( 
.A(n_2715),
.Y(n_3248)
);

OAI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_3069),
.A2(n_2650),
.B1(n_992),
.B2(n_1010),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3085),
.B(n_2560),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2769),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3087),
.B(n_2560),
.Y(n_3252)
);

OAI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_2834),
.A2(n_2392),
.B1(n_2419),
.B2(n_2397),
.Y(n_3253)
);

BUFx3_ASAP7_75t_L g3254 ( 
.A(n_2976),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_2881),
.B(n_2623),
.Y(n_3255)
);

NAND3xp33_ASAP7_75t_L g3256 ( 
.A(n_2757),
.B(n_1685),
.C(n_2064),
.Y(n_3256)
);

INVxp67_ASAP7_75t_L g3257 ( 
.A(n_2792),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2991),
.B(n_2564),
.Y(n_3258)
);

OAI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_2858),
.A2(n_2397),
.B1(n_2419),
.B2(n_2429),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_SL g3260 ( 
.A(n_3059),
.B(n_2623),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3078),
.B(n_2369),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2992),
.B(n_2564),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2770),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2771),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2916),
.Y(n_3265)
);

A2O1A1Ixp33_ASAP7_75t_L g3266 ( 
.A1(n_2990),
.A2(n_2671),
.B(n_2429),
.C(n_2494),
.Y(n_3266)
);

NOR2xp33_ASAP7_75t_L g3267 ( 
.A(n_2922),
.B(n_3040),
.Y(n_3267)
);

AND2x2_ASAP7_75t_L g3268 ( 
.A(n_3030),
.B(n_1842),
.Y(n_3268)
);

NOR2xp67_ASAP7_75t_L g3269 ( 
.A(n_2742),
.B(n_2565),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_L g3270 ( 
.A(n_3021),
.B(n_2429),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2927),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2772),
.Y(n_3272)
);

NOR2xp33_ASAP7_75t_L g3273 ( 
.A(n_3086),
.B(n_2467),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2776),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3080),
.B(n_2565),
.Y(n_3275)
);

NOR2xp33_ASAP7_75t_L g3276 ( 
.A(n_3086),
.B(n_2467),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_3084),
.B(n_2369),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_2764),
.Y(n_3278)
);

INVx2_ASAP7_75t_L g3279 ( 
.A(n_3004),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_SL g3280 ( 
.A(n_2757),
.B(n_2411),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2990),
.B(n_2996),
.Y(n_3281)
);

HB1xp67_ASAP7_75t_L g3282 ( 
.A(n_2954),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2724),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2996),
.B(n_2566),
.Y(n_3284)
);

INVxp33_ASAP7_75t_L g3285 ( 
.A(n_2731),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_SL g3286 ( 
.A(n_2741),
.B(n_2411),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2778),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2725),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2779),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3070),
.B(n_2566),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2726),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3071),
.B(n_2569),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_2893),
.A2(n_2063),
.B1(n_2074),
.B2(n_2072),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3077),
.B(n_2569),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3022),
.B(n_2571),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_3038),
.B(n_2467),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2727),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_SL g3298 ( 
.A(n_2741),
.B(n_2411),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3023),
.B(n_3028),
.Y(n_3299)
);

A2O1A1Ixp33_ASAP7_75t_L g3300 ( 
.A1(n_2858),
.A2(n_2671),
.B(n_2494),
.C(n_2505),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2783),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2729),
.Y(n_3302)
);

NAND3xp33_ASAP7_75t_L g3303 ( 
.A(n_2800),
.B(n_2144),
.C(n_2064),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3029),
.B(n_2571),
.Y(n_3304)
);

INVx3_ASAP7_75t_L g3305 ( 
.A(n_2903),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2967),
.B(n_2863),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3036),
.B(n_2573),
.Y(n_3307)
);

NAND2xp33_ASAP7_75t_L g3308 ( 
.A(n_2903),
.B(n_2650),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2870),
.B(n_2494),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3041),
.B(n_2573),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3042),
.B(n_3043),
.Y(n_3311)
);

HB1xp67_ASAP7_75t_L g3312 ( 
.A(n_2801),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3046),
.B(n_2574),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2831),
.B(n_2574),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_2835),
.B(n_2578),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3014),
.B(n_1842),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2836),
.B(n_2578),
.Y(n_3317)
);

BUFx2_ASAP7_75t_L g3318 ( 
.A(n_2728),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2837),
.B(n_2579),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2784),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_3011),
.Y(n_3321)
);

AND2x6_ASAP7_75t_SL g3322 ( 
.A(n_3009),
.B(n_2961),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2838),
.B(n_2839),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2840),
.B(n_2579),
.Y(n_3324)
);

INVx8_ASAP7_75t_L g3325 ( 
.A(n_2894),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_2734),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2788),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2740),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2841),
.B(n_2585),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2791),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2845),
.B(n_2585),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_2803),
.B(n_2712),
.Y(n_3332)
);

OR2x2_ASAP7_75t_L g3333 ( 
.A(n_2716),
.B(n_2602),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2847),
.B(n_2587),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2793),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_2894),
.B(n_2411),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2850),
.B(n_2587),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_2852),
.B(n_2602),
.Y(n_3338)
);

OAI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_2904),
.A2(n_2650),
.B1(n_1017),
.B2(n_1039),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2854),
.B(n_2603),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2743),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2855),
.B(n_2603),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2744),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3020),
.B(n_2500),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2795),
.Y(n_3345)
);

OAI22xp5_ASAP7_75t_L g3346 ( 
.A1(n_2948),
.A2(n_2505),
.B1(n_2529),
.B2(n_2500),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_2822),
.A2(n_2948),
.B1(n_2797),
.B2(n_2798),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2907),
.B(n_2500),
.Y(n_3348)
);

INVx2_ASAP7_75t_SL g3349 ( 
.A(n_3065),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2796),
.B(n_2612),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2804),
.B(n_2612),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_2931),
.A2(n_2944),
.B1(n_3035),
.B2(n_3024),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2811),
.B(n_2616),
.Y(n_3353)
);

HB1xp67_ASAP7_75t_L g3354 ( 
.A(n_2903),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_SL g3355 ( 
.A(n_2897),
.B(n_2411),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2869),
.B(n_2616),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2886),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_2932),
.B(n_2505),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2745),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2887),
.Y(n_3360)
);

INVxp33_ASAP7_75t_L g3361 ( 
.A(n_2760),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_2872),
.B(n_2622),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2890),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2891),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_2872),
.B(n_2622),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2884),
.B(n_2633),
.Y(n_3366)
);

BUFx3_ASAP7_75t_L g3367 ( 
.A(n_3075),
.Y(n_3367)
);

OAI22xp5_ASAP7_75t_L g3368 ( 
.A1(n_2884),
.A2(n_2540),
.B1(n_2542),
.B2(n_2529),
.Y(n_3368)
);

INVx2_ASAP7_75t_SL g3369 ( 
.A(n_3075),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_2897),
.B(n_1280),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2895),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2747),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2748),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2812),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_2928),
.B(n_2489),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_2902),
.A2(n_1084),
.B1(n_1090),
.B2(n_1081),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2905),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_2909),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_2843),
.B(n_2529),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_2843),
.B(n_2540),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2910),
.B(n_2633),
.Y(n_3381)
);

BUFx12f_ASAP7_75t_SL g3382 ( 
.A(n_3009),
.Y(n_3382)
);

NOR2xp67_ASAP7_75t_SL g3383 ( 
.A(n_2833),
.B(n_2513),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2911),
.B(n_2634),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_2928),
.B(n_2489),
.Y(n_3385)
);

BUFx6f_ASAP7_75t_SL g3386 ( 
.A(n_2961),
.Y(n_3386)
);

INVx3_ASAP7_75t_L g3387 ( 
.A(n_2888),
.Y(n_3387)
);

HB1xp67_ASAP7_75t_L g3388 ( 
.A(n_2829),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2912),
.Y(n_3389)
);

AND2x2_ASAP7_75t_L g3390 ( 
.A(n_2988),
.B(n_1369),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2913),
.B(n_2634),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_SL g3392 ( 
.A1(n_2873),
.A2(n_2650),
.B1(n_1046),
.B2(n_1058),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_SL g3393 ( 
.A(n_2904),
.B(n_2489),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2914),
.B(n_2639),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_2815),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2917),
.Y(n_3396)
);

INVx2_ASAP7_75t_SL g3397 ( 
.A(n_2959),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_2919),
.B(n_2639),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_2924),
.B(n_2644),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_L g3400 ( 
.A(n_2958),
.B(n_2540),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3076),
.B(n_3032),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2816),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_2925),
.Y(n_3403)
);

O2A1O1Ixp5_ASAP7_75t_L g3404 ( 
.A1(n_2714),
.A2(n_2646),
.B(n_2647),
.C(n_2644),
.Y(n_3404)
);

NOR2xp33_ASAP7_75t_L g3405 ( 
.A(n_2964),
.B(n_2542),
.Y(n_3405)
);

AND2x4_ASAP7_75t_L g3406 ( 
.A(n_2959),
.B(n_2646),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2926),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2933),
.B(n_2647),
.Y(n_3408)
);

NOR2x1p5_ASAP7_75t_L g3409 ( 
.A(n_2755),
.B(n_2773),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3032),
.B(n_2489),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_2936),
.B(n_2542),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2818),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_2794),
.A2(n_2898),
.B1(n_2787),
.B2(n_2888),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_SL g3414 ( 
.A(n_3000),
.B(n_2489),
.Y(n_3414)
);

O2A1O1Ixp5_ASAP7_75t_L g3415 ( 
.A1(n_2714),
.A2(n_2649),
.B(n_2666),
.C(n_2662),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2935),
.Y(n_3416)
);

INVx3_ASAP7_75t_L g3417 ( 
.A(n_2945),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_2819),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2820),
.Y(n_3419)
);

OAI221xp5_ASAP7_75t_L g3420 ( 
.A1(n_3072),
.A2(n_835),
.B1(n_1112),
.B2(n_1106),
.C(n_1096),
.Y(n_3420)
);

OR2x2_ASAP7_75t_L g3421 ( 
.A(n_2762),
.B(n_2649),
.Y(n_3421)
);

NOR2xp33_ASAP7_75t_L g3422 ( 
.A(n_3045),
.B(n_2983),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2937),
.B(n_2608),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3283),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3137),
.B(n_2983),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3127),
.B(n_3000),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_3148),
.A2(n_2422),
.B(n_2693),
.Y(n_3427)
);

AND2x2_ASAP7_75t_L g3428 ( 
.A(n_3141),
.B(n_3003),
.Y(n_3428)
);

AND2x4_ASAP7_75t_L g3429 ( 
.A(n_3119),
.B(n_3003),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3288),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3281),
.B(n_2939),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3149),
.A2(n_2422),
.B(n_2693),
.Y(n_3432)
);

INVxp67_ASAP7_75t_L g3433 ( 
.A(n_3118),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3184),
.B(n_2873),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3208),
.B(n_2856),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3151),
.B(n_2862),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3120),
.A2(n_2422),
.B(n_2693),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3151),
.B(n_2875),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3136),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_3206),
.B(n_2987),
.Y(n_3440)
);

BUFx12f_ASAP7_75t_L g3441 ( 
.A(n_3180),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_3108),
.B(n_3109),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3108),
.B(n_1888),
.Y(n_3443)
);

A2O1A1Ixp33_ASAP7_75t_L g3444 ( 
.A1(n_3146),
.A2(n_2929),
.B(n_2940),
.C(n_2879),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3122),
.B(n_3205),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3107),
.B(n_2942),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3129),
.A2(n_2422),
.B(n_2654),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3210),
.B(n_3100),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3285),
.B(n_1888),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3103),
.B(n_2946),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3242),
.A2(n_2945),
.B1(n_2787),
.B2(n_2898),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3130),
.A2(n_2663),
.B(n_2655),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3155),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3213),
.A2(n_2548),
.B(n_2544),
.Y(n_3454)
);

INVx1_ASAP7_75t_SL g3455 ( 
.A(n_3118),
.Y(n_3455)
);

INVx4_ASAP7_75t_L g3456 ( 
.A(n_3155),
.Y(n_3456)
);

AND2x2_ASAP7_75t_L g3457 ( 
.A(n_3153),
.B(n_2777),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3291),
.Y(n_3458)
);

AO21x1_ASAP7_75t_L g3459 ( 
.A1(n_3093),
.A2(n_3193),
.B(n_3094),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3242),
.A2(n_2548),
.B(n_2544),
.Y(n_3460)
);

AOI21xp5_ASAP7_75t_L g3461 ( 
.A1(n_3144),
.A2(n_2630),
.B(n_2554),
.Y(n_3461)
);

AOI21xp5_ASAP7_75t_L g3462 ( 
.A1(n_3145),
.A2(n_2630),
.B(n_2554),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_3178),
.B(n_2899),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3138),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3404),
.A2(n_3017),
.B(n_2864),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3146),
.B(n_2738),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3297),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3106),
.A2(n_2593),
.B(n_2493),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3259),
.A2(n_3346),
.B(n_3185),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_3110),
.A2(n_3135),
.B(n_3157),
.Y(n_3470)
);

INVxp67_ASAP7_75t_L g3471 ( 
.A(n_3282),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3163),
.B(n_2739),
.Y(n_3472)
);

INVx2_ASAP7_75t_SL g3473 ( 
.A(n_3104),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3090),
.Y(n_3474)
);

AND2x6_ASAP7_75t_L g3475 ( 
.A(n_3387),
.B(n_2561),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3302),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3123),
.B(n_3176),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3179),
.B(n_2947),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3142),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_3101),
.B(n_2880),
.Y(n_3480)
);

OAI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3193),
.A2(n_2688),
.B(n_2950),
.Y(n_3481)
);

NAND2x1p5_ASAP7_75t_L g3482 ( 
.A(n_3383),
.B(n_2953),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3159),
.A2(n_2593),
.B(n_2493),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3097),
.A2(n_3005),
.B1(n_2923),
.B2(n_3037),
.Y(n_3484)
);

AOI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_3227),
.A2(n_2593),
.B(n_2493),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3231),
.A2(n_3266),
.B(n_3300),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_3413),
.A2(n_2593),
.B(n_2493),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3232),
.B(n_2957),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3306),
.B(n_2952),
.Y(n_3489)
);

OA21x2_ASAP7_75t_L g3490 ( 
.A1(n_3243),
.A2(n_2864),
.B(n_3017),
.Y(n_3490)
);

O2A1O1Ixp5_ASAP7_75t_L g3491 ( 
.A1(n_3092),
.A2(n_3049),
.B(n_3039),
.C(n_2823),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_3097),
.A2(n_2547),
.B1(n_2570),
.B2(n_2359),
.Y(n_3492)
);

AND2x2_ASAP7_75t_L g3493 ( 
.A(n_3370),
.B(n_2813),
.Y(n_3493)
);

O2A1O1Ixp33_ASAP7_75t_L g3494 ( 
.A1(n_3420),
.A2(n_2085),
.B(n_2088),
.C(n_2084),
.Y(n_3494)
);

AOI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3154),
.A2(n_2915),
.B1(n_2934),
.B2(n_2883),
.Y(n_3495)
);

OAI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_3116),
.A2(n_2966),
.B(n_2962),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3203),
.B(n_2968),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3183),
.A2(n_2593),
.B(n_2493),
.Y(n_3498)
);

AOI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_3169),
.A2(n_2092),
.B1(n_2094),
.B2(n_2093),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3215),
.B(n_2970),
.Y(n_3500)
);

AOI21x1_ASAP7_75t_L g3501 ( 
.A1(n_3243),
.A2(n_3049),
.B(n_3039),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3344),
.B(n_1437),
.Y(n_3502)
);

INVx4_ASAP7_75t_L g3503 ( 
.A(n_3155),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3154),
.B(n_2972),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_3326),
.Y(n_3505)
);

OAI321xp33_ASAP7_75t_L g3506 ( 
.A1(n_3339),
.A2(n_1102),
.A3(n_1090),
.B1(n_1104),
.B2(n_1099),
.C(n_1084),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3358),
.B(n_2943),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3169),
.B(n_2973),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3253),
.A2(n_2682),
.B(n_2598),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3140),
.A2(n_2682),
.B(n_2598),
.Y(n_3510)
);

NOR2xp33_ASAP7_75t_L g3511 ( 
.A(n_3306),
.B(n_3358),
.Y(n_3511)
);

INVxp67_ASAP7_75t_SL g3512 ( 
.A(n_3150),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3309),
.B(n_2978),
.Y(n_3513)
);

O2A1O1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_3131),
.A2(n_3095),
.B(n_3249),
.C(n_3339),
.Y(n_3514)
);

A2O1A1Ixp33_ASAP7_75t_L g3515 ( 
.A1(n_3309),
.A2(n_2982),
.B(n_2984),
.C(n_2980),
.Y(n_3515)
);

O2A1O1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_3095),
.A2(n_2105),
.B(n_2106),
.C(n_2096),
.Y(n_3516)
);

AOI21x1_ASAP7_75t_L g3517 ( 
.A1(n_3139),
.A2(n_2678),
.B(n_2670),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3268),
.B(n_2986),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3147),
.A2(n_2682),
.B(n_2598),
.Y(n_3519)
);

BUFx4f_ASAP7_75t_L g3520 ( 
.A(n_3132),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3344),
.B(n_2989),
.Y(n_3521)
);

AO21x1_ASAP7_75t_L g3522 ( 
.A1(n_3094),
.A2(n_2825),
.B(n_2821),
.Y(n_3522)
);

O2A1O1Ixp33_ASAP7_75t_L g3523 ( 
.A1(n_3249),
.A2(n_2114),
.B(n_2116),
.C(n_2112),
.Y(n_3523)
);

INVx3_ASAP7_75t_L g3524 ( 
.A(n_3387),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3308),
.A2(n_3221),
.B(n_3219),
.Y(n_3525)
);

NAND3xp33_ASAP7_75t_SL g3526 ( 
.A(n_3207),
.B(n_2993),
.C(n_2759),
.Y(n_3526)
);

A2O1A1Ixp33_ASAP7_75t_L g3527 ( 
.A1(n_3099),
.A2(n_2998),
.B(n_3001),
.C(n_2995),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3284),
.A2(n_2682),
.B(n_2598),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3152),
.A2(n_2682),
.B(n_2598),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_3392),
.B(n_2761),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3152),
.A2(n_2684),
.B(n_2551),
.Y(n_3531)
);

OAI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_3164),
.A2(n_2611),
.B1(n_3007),
.B2(n_3006),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3161),
.B(n_3008),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3328),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3341),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3112),
.B(n_2749),
.Y(n_3536)
);

BUFx3_ASAP7_75t_L g3537 ( 
.A(n_3117),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3166),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3270),
.B(n_3015),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3172),
.Y(n_3540)
);

O2A1O1Ixp5_ASAP7_75t_L g3541 ( 
.A1(n_3393),
.A2(n_2826),
.B(n_2830),
.C(n_2827),
.Y(n_3541)
);

OAI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_3121),
.A2(n_3013),
.B(n_3012),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3270),
.B(n_3016),
.Y(n_3543)
);

A2O1A1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3347),
.A2(n_3018),
.B(n_3019),
.C(n_2679),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3182),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3220),
.A2(n_2684),
.B(n_2551),
.Y(n_3546)
);

OR2x2_ASAP7_75t_L g3547 ( 
.A(n_3333),
.B(n_3034),
.Y(n_3547)
);

HB1xp67_ASAP7_75t_L g3548 ( 
.A(n_3282),
.Y(n_3548)
);

AOI33xp33_ASAP7_75t_L g3549 ( 
.A1(n_3392),
.A2(n_1140),
.A3(n_1125),
.B1(n_1418),
.B2(n_1420),
.B3(n_1417),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3220),
.A2(n_2684),
.B(n_2395),
.Y(n_3550)
);

AOI21xp5_ASAP7_75t_L g3551 ( 
.A1(n_3356),
.A2(n_2684),
.B(n_2395),
.Y(n_3551)
);

BUFx2_ASAP7_75t_L g3552 ( 
.A(n_3168),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3195),
.B(n_2829),
.Y(n_3553)
);

AOI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3362),
.A2(n_3366),
.B(n_3365),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3421),
.B(n_3390),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3170),
.A2(n_2684),
.B(n_2395),
.Y(n_3556)
);

NOR2xp67_ASAP7_75t_L g3557 ( 
.A(n_3267),
.B(n_2733),
.Y(n_3557)
);

O2A1O1Ixp33_ASAP7_75t_L g3558 ( 
.A1(n_3217),
.A2(n_2123),
.B(n_2124),
.C(n_2119),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3173),
.A2(n_2533),
.B(n_2380),
.Y(n_3559)
);

AOI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3165),
.A2(n_2533),
.B(n_2380),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_L g3561 ( 
.A(n_3112),
.B(n_2144),
.Y(n_3561)
);

AND2x2_ASAP7_75t_SL g3562 ( 
.A(n_3238),
.B(n_3066),
.Y(n_3562)
);

AOI21x1_ASAP7_75t_L g3563 ( 
.A1(n_3223),
.A2(n_2666),
.B(n_2662),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3195),
.B(n_2829),
.Y(n_3564)
);

OR2x2_ASAP7_75t_L g3565 ( 
.A(n_3241),
.B(n_3177),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3316),
.B(n_1445),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3332),
.B(n_2144),
.Y(n_3567)
);

AOI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3124),
.A2(n_2533),
.B(n_2380),
.Y(n_3568)
);

AND2x4_ASAP7_75t_L g3569 ( 
.A(n_3119),
.B(n_2843),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3124),
.A2(n_2551),
.B(n_2354),
.Y(n_3570)
);

INVx2_ASAP7_75t_SL g3571 ( 
.A(n_3321),
.Y(n_3571)
);

AOI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_3280),
.A2(n_2354),
.B(n_2325),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_3368),
.A2(n_2354),
.B(n_2325),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3343),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3201),
.B(n_2829),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3359),
.Y(n_3576)
);

OAI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3121),
.A2(n_2680),
.B(n_2673),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3372),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_SL g3579 ( 
.A(n_3113),
.B(n_2810),
.Y(n_3579)
);

INVx2_ASAP7_75t_SL g3580 ( 
.A(n_3349),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3098),
.A2(n_2354),
.B(n_2325),
.Y(n_3581)
);

AOI21xp5_ASAP7_75t_L g3582 ( 
.A1(n_3102),
.A2(n_2354),
.B(n_2325),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3201),
.B(n_2126),
.Y(n_3583)
);

O2A1O1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_3217),
.A2(n_2135),
.B(n_2140),
.C(n_2137),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3188),
.Y(n_3585)
);

OAI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3275),
.A2(n_3262),
.B(n_3258),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3192),
.Y(n_3587)
);

HB1xp67_ASAP7_75t_L g3588 ( 
.A(n_3150),
.Y(n_3588)
);

OAI22xp5_ASAP7_75t_L g3589 ( 
.A1(n_3164),
.A2(n_2594),
.B1(n_2561),
.B2(n_2608),
.Y(n_3589)
);

NOR2xp33_ASAP7_75t_SL g3590 ( 
.A(n_3175),
.B(n_3066),
.Y(n_3590)
);

BUFx6f_ASAP7_75t_L g3591 ( 
.A(n_3155),
.Y(n_3591)
);

AND2x2_ASAP7_75t_L g3592 ( 
.A(n_3411),
.B(n_1473),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3379),
.A2(n_2440),
.B(n_2325),
.Y(n_3593)
);

INVxp67_ASAP7_75t_L g3594 ( 
.A(n_3312),
.Y(n_3594)
);

A2O1A1Ixp33_ASAP7_75t_L g3595 ( 
.A1(n_3347),
.A2(n_2594),
.B(n_2561),
.C(n_2143),
.Y(n_3595)
);

CKINVDCx10_ASAP7_75t_R g3596 ( 
.A(n_3386),
.Y(n_3596)
);

INVx4_ASAP7_75t_L g3597 ( 
.A(n_3209),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3348),
.B(n_2141),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3348),
.B(n_2157),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3379),
.A2(n_2442),
.B(n_2440),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_3417),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3240),
.B(n_2164),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3240),
.B(n_2165),
.Y(n_3603)
);

OAI21xp33_ASAP7_75t_L g3604 ( 
.A1(n_3091),
.A2(n_2866),
.B(n_2802),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_SL g3605 ( 
.A(n_3113),
.B(n_2824),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3105),
.Y(n_3606)
);

OAI21xp33_ASAP7_75t_L g3607 ( 
.A1(n_3091),
.A2(n_856),
.B(n_853),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_3373),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3374),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3332),
.B(n_2711),
.Y(n_3610)
);

BUFx6f_ASAP7_75t_L g3611 ( 
.A(n_3209),
.Y(n_3611)
);

A2O1A1Ixp33_ASAP7_75t_L g3612 ( 
.A1(n_3400),
.A2(n_2594),
.B(n_2180),
.C(n_2181),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3181),
.B(n_2713),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3111),
.Y(n_3614)
);

AND2x4_ASAP7_75t_L g3615 ( 
.A(n_3397),
.B(n_2851),
.Y(n_3615)
);

A2O1A1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_3400),
.A2(n_2182),
.B(n_2183),
.C(n_2175),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3380),
.A2(n_2442),
.B(n_2440),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3114),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3209),
.Y(n_3619)
);

INVxp67_ASAP7_75t_L g3620 ( 
.A(n_3312),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3380),
.A2(n_2442),
.B(n_2440),
.Y(n_3621)
);

INVx3_ASAP7_75t_L g3622 ( 
.A(n_3417),
.Y(n_3622)
);

AOI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3405),
.A2(n_2185),
.B1(n_1029),
.B2(n_1044),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3411),
.B(n_2842),
.Y(n_3624)
);

BUFx6f_ASAP7_75t_L g3625 ( 
.A(n_3209),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_L g3626 ( 
.A(n_3296),
.B(n_2608),
.Y(n_3626)
);

BUFx12f_ASAP7_75t_L g3627 ( 
.A(n_3180),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3296),
.B(n_2618),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_SL g3629 ( 
.A(n_3352),
.B(n_3267),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_3255),
.A2(n_2442),
.B(n_2440),
.Y(n_3630)
);

AND2x4_ASAP7_75t_L g3631 ( 
.A(n_3115),
.B(n_2851),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3199),
.B(n_2618),
.Y(n_3632)
);

INVx3_ASAP7_75t_L g3633 ( 
.A(n_3115),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3405),
.A2(n_3025),
.B1(n_2631),
.B2(n_2618),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3134),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3260),
.A2(n_2508),
.B(n_2442),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3395),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3299),
.B(n_2631),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3202),
.A2(n_2508),
.B(n_2637),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3311),
.B(n_2631),
.Y(n_3640)
);

AOI21xp33_ASAP7_75t_L g3641 ( 
.A1(n_3218),
.A2(n_2842),
.B(n_2882),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3198),
.B(n_2673),
.Y(n_3642)
);

BUFx2_ASAP7_75t_SL g3643 ( 
.A(n_3125),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3198),
.B(n_3191),
.Y(n_3644)
);

OAI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3244),
.A2(n_2681),
.B(n_2680),
.Y(n_3645)
);

AND2x4_ASAP7_75t_L g3646 ( 
.A(n_3401),
.B(n_3406),
.Y(n_3646)
);

AOI21xp5_ASAP7_75t_L g3647 ( 
.A1(n_3200),
.A2(n_2508),
.B(n_2409),
.Y(n_3647)
);

OAI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3245),
.A2(n_2672),
.B1(n_2691),
.B2(n_2657),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_SL g3649 ( 
.A(n_3218),
.B(n_1876),
.Y(n_3649)
);

INVxp67_ASAP7_75t_L g3650 ( 
.A(n_3318),
.Y(n_3650)
);

BUFx2_ASAP7_75t_L g3651 ( 
.A(n_3257),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3273),
.B(n_2681),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3273),
.B(n_2692),
.Y(n_3653)
);

AOI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3381),
.A2(n_3391),
.B(n_3384),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3276),
.B(n_2692),
.Y(n_3655)
);

OAI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_3404),
.A2(n_2700),
.B(n_2695),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3276),
.B(n_2695),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3323),
.A2(n_2508),
.B(n_2409),
.Y(n_3658)
);

AOI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3415),
.A2(n_2508),
.B(n_2409),
.Y(n_3659)
);

AOI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_3415),
.A2(n_2381),
.B(n_1996),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3269),
.A2(n_3414),
.B(n_3410),
.Y(n_3661)
);

NOR2xp33_ASAP7_75t_L g3662 ( 
.A(n_3361),
.B(n_2842),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3228),
.B(n_2700),
.Y(n_3663)
);

AND2x2_ASAP7_75t_SL g3664 ( 
.A(n_3238),
.B(n_1099),
.Y(n_3664)
);

A2O1A1Ixp33_ASAP7_75t_L g3665 ( 
.A1(n_3293),
.A2(n_2706),
.B(n_2657),
.C(n_2691),
.Y(n_3665)
);

INVx4_ASAP7_75t_L g3666 ( 
.A(n_3132),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3402),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3162),
.A2(n_3315),
.B(n_3314),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3162),
.A2(n_2381),
.B(n_1996),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3229),
.B(n_2706),
.Y(n_3670)
);

NAND2xp33_ASAP7_75t_L g3671 ( 
.A(n_3132),
.B(n_3025),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3317),
.A2(n_2381),
.B(n_1996),
.Y(n_3672)
);

INVx1_ASAP7_75t_SL g3673 ( 
.A(n_3186),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3319),
.A2(n_1996),
.B(n_1979),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3235),
.B(n_3025),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_SL g3676 ( 
.A(n_3382),
.B(n_1876),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3324),
.A2(n_3331),
.B(n_3329),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_3334),
.A2(n_1981),
.B(n_1979),
.Y(n_3678)
);

OR2x2_ASAP7_75t_L g3679 ( 
.A(n_3257),
.B(n_2657),
.Y(n_3679)
);

AO21x1_ASAP7_75t_L g3680 ( 
.A1(n_3261),
.A2(n_2244),
.B(n_2240),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3128),
.B(n_1424),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3470),
.A2(n_3388),
.B(n_3197),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3439),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3464),
.Y(n_3684)
);

NOR2xp67_ASAP7_75t_L g3685 ( 
.A(n_3445),
.B(n_3412),
.Y(n_3685)
);

XOR2x2_ASAP7_75t_SL g3686 ( 
.A(n_3495),
.B(n_3248),
.Y(n_3686)
);

A2O1A1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3514),
.A2(n_3214),
.B(n_3256),
.C(n_3239),
.Y(n_3687)
);

O2A1O1Ixp5_ASAP7_75t_L g3688 ( 
.A1(n_3442),
.A2(n_3459),
.B(n_3530),
.C(n_3511),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3479),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3466),
.B(n_3226),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3538),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3448),
.B(n_3236),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3424),
.Y(n_3693)
);

OAI22xp5_ASAP7_75t_L g3694 ( 
.A1(n_3495),
.A2(n_3422),
.B1(n_3222),
.B2(n_3174),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3477),
.B(n_3502),
.Y(n_3695)
);

INVx3_ASAP7_75t_L g3696 ( 
.A(n_3631),
.Y(n_3696)
);

O2A1O1Ixp33_ASAP7_75t_L g3697 ( 
.A1(n_3463),
.A2(n_3222),
.B(n_3204),
.C(n_3422),
.Y(n_3697)
);

INVx3_ASAP7_75t_L g3698 ( 
.A(n_3631),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_R g3699 ( 
.A(n_3590),
.B(n_3171),
.Y(n_3699)
);

INVx2_ASAP7_75t_SL g3700 ( 
.A(n_3537),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3428),
.B(n_3406),
.Y(n_3701)
);

A2O1A1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3549),
.A2(n_3251),
.B(n_3263),
.C(n_3247),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3447),
.A2(n_3388),
.B(n_3196),
.Y(n_3703)
);

INVxp33_ASAP7_75t_SL g3704 ( 
.A(n_3590),
.Y(n_3704)
);

OAI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_3673),
.A2(n_3521),
.B1(n_3426),
.B2(n_3425),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_SL g3706 ( 
.A(n_3664),
.B(n_3303),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_SL g3707 ( 
.A(n_3673),
.B(n_3278),
.Y(n_3707)
);

INVx1_ASAP7_75t_SL g3708 ( 
.A(n_3565),
.Y(n_3708)
);

BUFx8_ASAP7_75t_L g3709 ( 
.A(n_3441),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3469),
.A2(n_3338),
.B(n_3337),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3567),
.B(n_3264),
.Y(n_3711)
);

BUFx2_ASAP7_75t_L g3712 ( 
.A(n_3474),
.Y(n_3712)
);

AO32x1_ASAP7_75t_L g3713 ( 
.A1(n_3532),
.A2(n_3363),
.A3(n_3364),
.B1(n_3360),
.B2(n_3357),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3555),
.B(n_3272),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3592),
.B(n_3274),
.Y(n_3715)
);

AOI22xp33_ASAP7_75t_L g3716 ( 
.A1(n_3526),
.A2(n_3386),
.B1(n_3325),
.B2(n_3189),
.Y(n_3716)
);

INVxp67_ASAP7_75t_L g3717 ( 
.A(n_3548),
.Y(n_3717)
);

AOI21x1_ASAP7_75t_L g3718 ( 
.A1(n_3669),
.A2(n_3398),
.B(n_3394),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_SL g3719 ( 
.A(n_3646),
.B(n_3287),
.Y(n_3719)
);

NOR2xp33_ASAP7_75t_L g3720 ( 
.A(n_3472),
.B(n_3194),
.Y(n_3720)
);

CKINVDCx20_ASAP7_75t_R g3721 ( 
.A(n_3457),
.Y(n_3721)
);

OAI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3489),
.A2(n_3289),
.B1(n_3320),
.B2(n_3301),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3566),
.B(n_3376),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_3554),
.A2(n_3342),
.B(n_3340),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3427),
.A2(n_3353),
.B(n_3350),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_3432),
.A2(n_3452),
.B(n_3525),
.Y(n_3726)
);

A2O1A1Ixp33_ASAP7_75t_L g3727 ( 
.A1(n_3506),
.A2(n_3330),
.B(n_3335),
.C(n_3327),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3604),
.A2(n_3325),
.B1(n_3189),
.B2(n_3418),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3540),
.Y(n_3729)
);

INVx4_ASAP7_75t_L g3730 ( 
.A(n_3520),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3646),
.B(n_3345),
.Y(n_3731)
);

NAND3xp33_ASAP7_75t_L g3732 ( 
.A(n_3623),
.B(n_3607),
.C(n_3604),
.Y(n_3732)
);

INVx2_ASAP7_75t_L g3733 ( 
.A(n_3430),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3465),
.A2(n_3408),
.B(n_3399),
.Y(n_3734)
);

A2O1A1Ixp33_ASAP7_75t_L g3735 ( 
.A1(n_3506),
.A2(n_3377),
.B(n_3378),
.C(n_3371),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3458),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3545),
.Y(n_3737)
);

A2O1A1Ixp33_ASAP7_75t_L g3738 ( 
.A1(n_3558),
.A2(n_3584),
.B(n_3494),
.C(n_3607),
.Y(n_3738)
);

BUFx2_ASAP7_75t_L g3739 ( 
.A(n_3552),
.Y(n_3739)
);

AOI21xp5_ASAP7_75t_L g3740 ( 
.A1(n_3437),
.A2(n_3351),
.B(n_3277),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3487),
.A2(n_3298),
.B(n_3286),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3629),
.B(n_3224),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3488),
.B(n_3376),
.Y(n_3743)
);

AND2x4_ASAP7_75t_L g3744 ( 
.A(n_3569),
.B(n_3409),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3486),
.A2(n_3336),
.B(n_3234),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3435),
.B(n_3419),
.Y(n_3746)
);

NAND2xp33_ASAP7_75t_R g3747 ( 
.A(n_3443),
.B(n_3187),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3493),
.B(n_3096),
.Y(n_3748)
);

INVx1_ASAP7_75t_SL g3749 ( 
.A(n_3455),
.Y(n_3749)
);

NOR2xp33_ASAP7_75t_SL g3750 ( 
.A(n_3562),
.B(n_3158),
.Y(n_3750)
);

OR2x6_ASAP7_75t_SL g3751 ( 
.A(n_3547),
.B(n_834),
.Y(n_3751)
);

OAI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3561),
.A2(n_3369),
.B1(n_3367),
.B2(n_3389),
.Y(n_3752)
);

BUFx3_ASAP7_75t_L g3753 ( 
.A(n_3473),
.Y(n_3753)
);

O2A1O1Ixp5_ASAP7_75t_L g3754 ( 
.A1(n_3434),
.A2(n_3375),
.B(n_3385),
.C(n_3355),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3585),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3504),
.B(n_3436),
.Y(n_3756)
);

A2O1A1Ixp33_ASAP7_75t_L g3757 ( 
.A1(n_3616),
.A2(n_3403),
.B(n_3407),
.C(n_3396),
.Y(n_3757)
);

AOI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3536),
.A2(n_3325),
.B1(n_3189),
.B2(n_1899),
.Y(n_3758)
);

AO32x1_ASAP7_75t_L g3759 ( 
.A1(n_3492),
.A2(n_3416),
.A3(n_1105),
.B1(n_1115),
.B2(n_1104),
.Y(n_3759)
);

CKINVDCx6p67_ASAP7_75t_R g3760 ( 
.A(n_3596),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3587),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3507),
.B(n_3254),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3677),
.A2(n_3246),
.B(n_3233),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_SL g3764 ( 
.A(n_3598),
.B(n_3290),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_3438),
.B(n_3126),
.Y(n_3765)
);

AO32x1_ASAP7_75t_L g3766 ( 
.A1(n_3451),
.A2(n_1115),
.A3(n_1121),
.B1(n_1105),
.B2(n_1102),
.Y(n_3766)
);

O2A1O1Ixp33_ASAP7_75t_L g3767 ( 
.A1(n_3649),
.A2(n_1124),
.B(n_1128),
.C(n_1121),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3599),
.A2(n_3294),
.B1(n_3292),
.B2(n_3313),
.Y(n_3768)
);

AOI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3660),
.A2(n_3423),
.B(n_3252),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3529),
.A2(n_3295),
.B(n_3250),
.Y(n_3770)
);

AO32x1_ASAP7_75t_L g3771 ( 
.A1(n_3648),
.A2(n_1128),
.A3(n_1133),
.B1(n_1129),
.B2(n_1124),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3531),
.A2(n_3307),
.B(n_3304),
.Y(n_3772)
);

AOI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3613),
.A2(n_859),
.B1(n_863),
.B2(n_861),
.Y(n_3773)
);

AOI21x1_ASAP7_75t_L g3774 ( 
.A1(n_3659),
.A2(n_3310),
.B(n_2240),
.Y(n_3774)
);

NOR2x1p5_ASAP7_75t_SL g3775 ( 
.A(n_3501),
.B(n_3133),
.Y(n_3775)
);

O2A1O1Ixp5_ASAP7_75t_L g3776 ( 
.A1(n_3522),
.A2(n_3305),
.B(n_3187),
.C(n_3156),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_R g3777 ( 
.A(n_3676),
.B(n_3212),
.Y(n_3777)
);

INVx3_ASAP7_75t_L g3778 ( 
.A(n_3569),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3467),
.Y(n_3779)
);

NOR2x1_ASAP7_75t_L g3780 ( 
.A(n_3666),
.B(n_3305),
.Y(n_3780)
);

OAI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3623),
.A2(n_3211),
.B1(n_3216),
.B2(n_3190),
.Y(n_3781)
);

CKINVDCx10_ASAP7_75t_R g3782 ( 
.A(n_3596),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3606),
.Y(n_3783)
);

OAI21xp33_ASAP7_75t_L g3784 ( 
.A1(n_3681),
.A2(n_870),
.B(n_866),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3460),
.A2(n_3354),
.B(n_2906),
.Y(n_3785)
);

OAI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3668),
.A2(n_3160),
.B(n_3143),
.Y(n_3786)
);

AO22x1_ASAP7_75t_L g3787 ( 
.A1(n_3662),
.A2(n_3512),
.B1(n_3624),
.B2(n_3449),
.Y(n_3787)
);

AOI21xp5_ASAP7_75t_L g3788 ( 
.A1(n_3560),
.A2(n_3354),
.B(n_2906),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3614),
.Y(n_3789)
);

INVx3_ASAP7_75t_L g3790 ( 
.A(n_3615),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3429),
.B(n_3167),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_SL g3792 ( 
.A(n_3455),
.B(n_3225),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3508),
.B(n_3230),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3618),
.Y(n_3794)
);

OAI22xp5_ASAP7_75t_L g3795 ( 
.A1(n_3484),
.A2(n_3265),
.B1(n_3271),
.B2(n_3237),
.Y(n_3795)
);

OA22x2_ASAP7_75t_L g3796 ( 
.A1(n_3433),
.A2(n_873),
.B1(n_875),
.B2(n_872),
.Y(n_3796)
);

INVx3_ASAP7_75t_L g3797 ( 
.A(n_3615),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3635),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3431),
.B(n_3279),
.Y(n_3799)
);

OAI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_3499),
.A2(n_2691),
.B1(n_2702),
.B2(n_2672),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3610),
.B(n_1430),
.Y(n_3801)
);

NAND2xp33_ASAP7_75t_L g3802 ( 
.A(n_3644),
.B(n_3025),
.Y(n_3802)
);

INVx2_ASAP7_75t_SL g3803 ( 
.A(n_3571),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3429),
.B(n_1432),
.Y(n_3804)
);

NOR2xp33_ASAP7_75t_SL g3805 ( 
.A(n_3520),
.B(n_1899),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3497),
.B(n_880),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3478),
.B(n_882),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_L g3808 ( 
.A(n_3650),
.B(n_3322),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3476),
.Y(n_3809)
);

HB1xp67_ASAP7_75t_L g3810 ( 
.A(n_3651),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3471),
.B(n_1610),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3634),
.A2(n_2702),
.B1(n_2672),
.B2(n_886),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3446),
.B(n_888),
.Y(n_3813)
);

BUFx8_ASAP7_75t_L g3814 ( 
.A(n_3627),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3533),
.B(n_893),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3505),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3647),
.A2(n_2906),
.B(n_2851),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3546),
.A2(n_2702),
.B(n_1996),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3534),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3550),
.A2(n_2004),
.B(n_1981),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3500),
.B(n_897),
.Y(n_3821)
);

A2O1A1Ixp33_ASAP7_75t_L g3822 ( 
.A1(n_3516),
.A2(n_1129),
.B(n_1143),
.C(n_1133),
.Y(n_3822)
);

AOI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3658),
.A2(n_2004),
.B(n_1981),
.Y(n_3823)
);

O2A1O1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_3612),
.A2(n_1143),
.B(n_1145),
.C(n_1123),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_3518),
.B(n_1022),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3676),
.B(n_1050),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3588),
.B(n_898),
.Y(n_3827)
);

CKINVDCx16_ASAP7_75t_R g3828 ( 
.A(n_3643),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3454),
.A2(n_3510),
.B(n_3498),
.Y(n_3829)
);

INVxp67_ASAP7_75t_L g3830 ( 
.A(n_3580),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_3480),
.B(n_3553),
.Y(n_3831)
);

AOI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3519),
.A2(n_2004),
.B(n_1981),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3539),
.B(n_900),
.Y(n_3833)
);

OAI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_3444),
.A2(n_2247),
.B(n_2237),
.Y(n_3834)
);

AOI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3481),
.A2(n_3450),
.B(n_3513),
.Y(n_3835)
);

O2A1O1Ixp33_ASAP7_75t_L g3836 ( 
.A1(n_3544),
.A2(n_1145),
.B(n_1436),
.C(n_1433),
.Y(n_3836)
);

NOR2xp67_ASAP7_75t_L g3837 ( 
.A(n_3666),
.B(n_2237),
.Y(n_3837)
);

OAI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3564),
.A2(n_901),
.B1(n_904),
.B2(n_902),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_L g3839 ( 
.A(n_3594),
.B(n_1610),
.Y(n_3839)
);

AOI22xp33_ASAP7_75t_L g3840 ( 
.A1(n_3641),
.A2(n_905),
.B1(n_907),
.B2(n_906),
.Y(n_3840)
);

AOI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3557),
.A2(n_3579),
.B1(n_3605),
.B2(n_3440),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3575),
.B(n_1052),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_3509),
.A2(n_2004),
.B(n_1981),
.Y(n_3843)
);

NOR2xp33_ASAP7_75t_L g3844 ( 
.A(n_3620),
.B(n_1053),
.Y(n_3844)
);

OAI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3583),
.A2(n_909),
.B1(n_914),
.B2(n_913),
.Y(n_3845)
);

A2O1A1Ixp33_ASAP7_75t_L g3846 ( 
.A1(n_3661),
.A2(n_1076),
.B(n_1087),
.C(n_1060),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3543),
.B(n_919),
.Y(n_3847)
);

INVx1_ASAP7_75t_SL g3848 ( 
.A(n_3679),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3535),
.B(n_3574),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3576),
.B(n_922),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3578),
.B(n_1088),
.Y(n_3851)
);

OAI22x1_ASAP7_75t_L g3852 ( 
.A1(n_3482),
.A2(n_3609),
.B1(n_3637),
.B2(n_3608),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3667),
.B(n_3602),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3603),
.B(n_931),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3586),
.B(n_1091),
.Y(n_3855)
);

O2A1O1Ixp33_ASAP7_75t_SL g3856 ( 
.A1(n_3595),
.A2(n_2248),
.B(n_2249),
.C(n_2247),
.Y(n_3856)
);

O2A1O1Ixp33_ASAP7_75t_L g3857 ( 
.A1(n_3515),
.A2(n_1441),
.B(n_1443),
.C(n_1442),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3626),
.B(n_3628),
.Y(n_3858)
);

O2A1O1Ixp33_ASAP7_75t_L g3859 ( 
.A1(n_3527),
.A2(n_1444),
.B(n_1448),
.C(n_1447),
.Y(n_3859)
);

O2A1O1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3523),
.A2(n_3496),
.B(n_3665),
.C(n_3491),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_3524),
.Y(n_3861)
);

NAND2x1p5_ASAP7_75t_L g3862 ( 
.A(n_3633),
.B(n_2217),
.Y(n_3862)
);

OAI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3461),
.A2(n_2249),
.B(n_2248),
.Y(n_3863)
);

INVx3_ASAP7_75t_L g3864 ( 
.A(n_3524),
.Y(n_3864)
);

O2A1O1Ixp5_ASAP7_75t_L g3865 ( 
.A1(n_3517),
.A2(n_2251),
.B(n_2253),
.C(n_2250),
.Y(n_3865)
);

AOI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3671),
.A2(n_1107),
.B1(n_1113),
.B2(n_1097),
.Y(n_3866)
);

OR2x2_ASAP7_75t_L g3867 ( 
.A(n_3663),
.B(n_3670),
.Y(n_3867)
);

O2A1O1Ixp33_ASAP7_75t_L g3868 ( 
.A1(n_3675),
.A2(n_1450),
.B(n_1455),
.C(n_1454),
.Y(n_3868)
);

A2O1A1Ixp33_ASAP7_75t_L g3869 ( 
.A1(n_3541),
.A2(n_1137),
.B(n_933),
.C(n_937),
.Y(n_3869)
);

INVx2_ASAP7_75t_SL g3870 ( 
.A(n_3453),
.Y(n_3870)
);

NOR2xp33_ASAP7_75t_L g3871 ( 
.A(n_3633),
.B(n_934),
.Y(n_3871)
);

AOI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3462),
.A2(n_2015),
.B(n_2004),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3652),
.B(n_939),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3468),
.A2(n_2028),
.B(n_2015),
.Y(n_3874)
);

AND2x2_ASAP7_75t_L g3875 ( 
.A(n_3456),
.B(n_1457),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3601),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_3653),
.B(n_940),
.Y(n_3877)
);

AOI22xp33_ASAP7_75t_L g3878 ( 
.A1(n_3542),
.A2(n_942),
.B1(n_944),
.B2(n_943),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3655),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3639),
.A2(n_2251),
.B(n_2250),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3601),
.Y(n_3881)
);

AOI21xp5_ASAP7_75t_L g3882 ( 
.A1(n_3483),
.A2(n_2028),
.B(n_2015),
.Y(n_3882)
);

AO21x1_ASAP7_75t_L g3883 ( 
.A1(n_3657),
.A2(n_2257),
.B(n_2253),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3622),
.Y(n_3884)
);

A2O1A1Ixp33_ASAP7_75t_SL g3885 ( 
.A1(n_3577),
.A2(n_2228),
.B(n_2256),
.C(n_2217),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3632),
.Y(n_3886)
);

OAI22xp5_ASAP7_75t_L g3887 ( 
.A1(n_3482),
.A2(n_3642),
.B1(n_3638),
.B2(n_3640),
.Y(n_3887)
);

INVx3_ASAP7_75t_L g3888 ( 
.A(n_3622),
.Y(n_3888)
);

AND2x2_ASAP7_75t_L g3889 ( 
.A(n_3456),
.B(n_1459),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3654),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3453),
.Y(n_3891)
);

AND2x4_ASAP7_75t_L g3892 ( 
.A(n_3503),
.B(n_2257),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3503),
.B(n_1460),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3597),
.B(n_3453),
.Y(n_3894)
);

O2A1O1Ixp33_ASAP7_75t_L g3895 ( 
.A1(n_3589),
.A2(n_1463),
.B(n_1465),
.C(n_1461),
.Y(n_3895)
);

OAI21x1_ASAP7_75t_L g3896 ( 
.A1(n_3656),
.A2(n_2264),
.B(n_2262),
.Y(n_3896)
);

AOI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3485),
.A2(n_2028),
.B(n_2015),
.Y(n_3897)
);

NOR2xp33_ASAP7_75t_L g3898 ( 
.A(n_3597),
.B(n_945),
.Y(n_3898)
);

A2O1A1Ixp33_ASAP7_75t_L g3899 ( 
.A1(n_3528),
.A2(n_947),
.B(n_952),
.C(n_950),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3591),
.Y(n_3900)
);

AOI21xp5_ASAP7_75t_L g3901 ( 
.A1(n_3551),
.A2(n_2028),
.B(n_2015),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3591),
.B(n_953),
.Y(n_3902)
);

INVx3_ASAP7_75t_L g3903 ( 
.A(n_3591),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3611),
.B(n_3619),
.Y(n_3904)
);

INVx5_ASAP7_75t_L g3905 ( 
.A(n_3611),
.Y(n_3905)
);

INVxp67_ASAP7_75t_L g3906 ( 
.A(n_3611),
.Y(n_3906)
);

NOR2xp33_ASAP7_75t_L g3907 ( 
.A(n_3619),
.B(n_954),
.Y(n_3907)
);

NOR2xp33_ASAP7_75t_L g3908 ( 
.A(n_3619),
.B(n_957),
.Y(n_3908)
);

HB1xp67_ASAP7_75t_L g3909 ( 
.A(n_3625),
.Y(n_3909)
);

AND2x4_ASAP7_75t_L g3910 ( 
.A(n_3625),
.B(n_2262),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_L g3911 ( 
.A(n_3625),
.B(n_958),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3645),
.B(n_2264),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3563),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3475),
.B(n_962),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3490),
.B(n_1468),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3568),
.A2(n_964),
.B1(n_971),
.B2(n_966),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3556),
.B(n_972),
.Y(n_3917)
);

OR2x2_ASAP7_75t_L g3918 ( 
.A(n_3708),
.B(n_3490),
.Y(n_3918)
);

AND2x2_ASAP7_75t_L g3919 ( 
.A(n_3701),
.B(n_1472),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3726),
.A2(n_3570),
.B(n_3672),
.Y(n_3920)
);

AOI21x1_ASAP7_75t_L g3921 ( 
.A1(n_3787),
.A2(n_3678),
.B(n_3674),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3695),
.B(n_974),
.Y(n_3922)
);

AOI21x1_ASAP7_75t_L g3923 ( 
.A1(n_3855),
.A2(n_3680),
.B(n_3582),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3683),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3705),
.B(n_975),
.Y(n_3925)
);

OAI21x1_ASAP7_75t_L g3926 ( 
.A1(n_3829),
.A2(n_3573),
.B(n_3559),
.Y(n_3926)
);

AOI211x1_ASAP7_75t_L g3927 ( 
.A1(n_3732),
.A2(n_1475),
.B(n_1479),
.C(n_1474),
.Y(n_3927)
);

NOR2xp33_ASAP7_75t_L g3928 ( 
.A(n_3690),
.B(n_976),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3756),
.B(n_978),
.Y(n_3929)
);

OAI21x1_ASAP7_75t_L g3930 ( 
.A1(n_3774),
.A2(n_3630),
.B(n_3572),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3684),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3817),
.A2(n_3581),
.B(n_3636),
.Y(n_3932)
);

AOI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3835),
.A2(n_3600),
.B(n_3593),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3689),
.Y(n_3934)
);

OAI21x1_ASAP7_75t_L g3935 ( 
.A1(n_3788),
.A2(n_3621),
.B(n_3617),
.Y(n_3935)
);

NOR2xp33_ASAP7_75t_L g3936 ( 
.A(n_3704),
.B(n_984),
.Y(n_3936)
);

NAND2xp33_ASAP7_75t_L g3937 ( 
.A(n_3777),
.B(n_3475),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_L g3938 ( 
.A(n_3753),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3691),
.Y(n_3939)
);

NOR2x1_ASAP7_75t_L g3940 ( 
.A(n_3685),
.B(n_1480),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3848),
.B(n_1482),
.Y(n_3941)
);

OAI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3688),
.A2(n_3475),
.B(n_2272),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3905),
.Y(n_3943)
);

AND2x2_ASAP7_75t_L g3944 ( 
.A(n_3748),
.B(n_1485),
.Y(n_3944)
);

OAI21x1_ASAP7_75t_L g3945 ( 
.A1(n_3865),
.A2(n_2272),
.B(n_2270),
.Y(n_3945)
);

OAI21x1_ASAP7_75t_L g3946 ( 
.A1(n_3823),
.A2(n_2277),
.B(n_2270),
.Y(n_3946)
);

OAI21x1_ASAP7_75t_L g3947 ( 
.A1(n_3785),
.A2(n_2285),
.B(n_2277),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3692),
.B(n_986),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3879),
.B(n_988),
.Y(n_3949)
);

OA21x2_ASAP7_75t_L g3950 ( 
.A1(n_3776),
.A2(n_1488),
.B(n_1487),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3853),
.B(n_989),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3746),
.B(n_990),
.Y(n_3952)
);

NOR2xp67_ASAP7_75t_SL g3953 ( 
.A(n_3828),
.B(n_1489),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_3782),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3724),
.A2(n_3475),
.B(n_2296),
.Y(n_3955)
);

OAI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3738),
.A2(n_2296),
.B(n_2285),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3729),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3763),
.A2(n_3710),
.B(n_3772),
.Y(n_3958)
);

BUFx3_ASAP7_75t_L g3959 ( 
.A(n_3712),
.Y(n_3959)
);

INVx3_ASAP7_75t_L g3960 ( 
.A(n_3730),
.Y(n_3960)
);

AOI21xp33_ASAP7_75t_L g3961 ( 
.A1(n_3916),
.A2(n_3697),
.B(n_3860),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3793),
.B(n_991),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3737),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_SL g3964 ( 
.A(n_3686),
.B(n_1491),
.Y(n_3964)
);

AOI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3725),
.A2(n_2298),
.B(n_2228),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_3770),
.A2(n_2298),
.B(n_2228),
.Y(n_3966)
);

NOR2xp33_ASAP7_75t_L g3967 ( 
.A(n_3711),
.B(n_994),
.Y(n_3967)
);

OAI21x1_ASAP7_75t_L g3968 ( 
.A1(n_3872),
.A2(n_1998),
.B(n_1992),
.Y(n_3968)
);

OA21x2_ASAP7_75t_L g3969 ( 
.A1(n_3734),
.A2(n_1494),
.B(n_1493),
.Y(n_3969)
);

INVxp67_ASAP7_75t_SL g3970 ( 
.A(n_3685),
.Y(n_3970)
);

OAI21x1_ASAP7_75t_SL g3971 ( 
.A1(n_3824),
.A2(n_1499),
.B(n_1497),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3714),
.B(n_996),
.Y(n_3972)
);

OAI21x1_ASAP7_75t_L g3973 ( 
.A1(n_3740),
.A2(n_1998),
.B(n_1992),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3765),
.B(n_1000),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3715),
.B(n_1003),
.Y(n_3975)
);

OAI21x1_ASAP7_75t_SL g3976 ( 
.A1(n_3741),
.A2(n_3745),
.B(n_3682),
.Y(n_3976)
);

OAI22xp5_ASAP7_75t_L g3977 ( 
.A1(n_3728),
.A2(n_1004),
.B1(n_1007),
.B2(n_1006),
.Y(n_3977)
);

AO21x1_ASAP7_75t_L g3978 ( 
.A1(n_3722),
.A2(n_1501),
.B(n_1500),
.Y(n_3978)
);

AOI21xp5_ASAP7_75t_L g3979 ( 
.A1(n_3764),
.A2(n_2256),
.B(n_2217),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3755),
.Y(n_3980)
);

OAI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3818),
.A2(n_1998),
.B(n_1992),
.Y(n_3981)
);

OAI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3687),
.A2(n_1503),
.B(n_1502),
.Y(n_3982)
);

OA22x2_ASAP7_75t_L g3983 ( 
.A1(n_3841),
.A2(n_1012),
.B1(n_1013),
.B2(n_1008),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_3799),
.B(n_1016),
.Y(n_3984)
);

INVxp67_ASAP7_75t_L g3985 ( 
.A(n_3810),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3761),
.Y(n_3986)
);

BUFx3_ASAP7_75t_L g3987 ( 
.A(n_3739),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3768),
.A2(n_2261),
.B(n_2256),
.Y(n_3988)
);

AOI21x1_ASAP7_75t_L g3989 ( 
.A1(n_3917),
.A2(n_1505),
.B(n_1504),
.Y(n_3989)
);

OAI22xp5_ASAP7_75t_L g3990 ( 
.A1(n_3723),
.A2(n_1020),
.B1(n_1026),
.B2(n_1019),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3749),
.B(n_1030),
.Y(n_3991)
);

OAI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3754),
.A2(n_3887),
.B(n_3869),
.Y(n_3992)
);

OR2x2_ASAP7_75t_L g3993 ( 
.A(n_3801),
.B(n_1506),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3886),
.B(n_3873),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3877),
.B(n_1032),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3693),
.Y(n_3996)
);

NOR2x1_ASAP7_75t_SL g3997 ( 
.A(n_3858),
.B(n_1508),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3791),
.B(n_3804),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3802),
.A2(n_2265),
.B(n_2261),
.Y(n_3999)
);

BUFx2_ASAP7_75t_L g4000 ( 
.A(n_3909),
.Y(n_4000)
);

OAI21x1_ASAP7_75t_L g4001 ( 
.A1(n_3820),
.A2(n_2012),
.B(n_2006),
.Y(n_4001)
);

OAI21x1_ASAP7_75t_L g4002 ( 
.A1(n_3863),
.A2(n_3896),
.B(n_3880),
.Y(n_4002)
);

OAI21x1_ASAP7_75t_L g4003 ( 
.A1(n_3843),
.A2(n_2012),
.B(n_2006),
.Y(n_4003)
);

OAI21x1_ASAP7_75t_L g4004 ( 
.A1(n_3703),
.A2(n_2012),
.B(n_2006),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3733),
.Y(n_4005)
);

AOI22xp33_ASAP7_75t_SL g4006 ( 
.A1(n_3694),
.A2(n_1036),
.B1(n_1042),
.B2(n_1034),
.Y(n_4006)
);

AOI221x1_ASAP7_75t_L g4007 ( 
.A1(n_3852),
.A2(n_1511),
.B1(n_1516),
.B2(n_1510),
.C(n_1509),
.Y(n_4007)
);

OAI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3786),
.A2(n_1518),
.B(n_1517),
.Y(n_4008)
);

AOI21x1_ASAP7_75t_SL g4009 ( 
.A1(n_3914),
.A2(n_686),
.B(n_1198),
.Y(n_4009)
);

BUFx2_ASAP7_75t_L g4010 ( 
.A(n_3894),
.Y(n_4010)
);

BUFx2_ASAP7_75t_SL g4011 ( 
.A(n_3721),
.Y(n_4011)
);

OAI21x1_ASAP7_75t_L g4012 ( 
.A1(n_3897),
.A2(n_2060),
.B(n_2032),
.Y(n_4012)
);

OAI22xp5_ASAP7_75t_L g4013 ( 
.A1(n_3716),
.A2(n_1033),
.B1(n_1051),
.B2(n_1048),
.Y(n_4013)
);

A2O1A1Ixp33_ASAP7_75t_L g4014 ( 
.A1(n_3742),
.A2(n_1524),
.B(n_1525),
.C(n_1521),
.Y(n_4014)
);

OAI21x1_ASAP7_75t_L g4015 ( 
.A1(n_3718),
.A2(n_2060),
.B(n_2032),
.Y(n_4015)
);

O2A1O1Ixp5_ASAP7_75t_L g4016 ( 
.A1(n_3706),
.A2(n_1527),
.B(n_1528),
.C(n_1526),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3783),
.Y(n_4017)
);

OAI21x1_ASAP7_75t_L g4018 ( 
.A1(n_3882),
.A2(n_2060),
.B(n_2032),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_SL g4019 ( 
.A1(n_3846),
.A2(n_686),
.B(n_1055),
.Y(n_4019)
);

OAI21x1_ASAP7_75t_L g4020 ( 
.A1(n_3901),
.A2(n_2200),
.B(n_2079),
.Y(n_4020)
);

OAI21x1_ASAP7_75t_L g4021 ( 
.A1(n_3769),
.A2(n_2200),
.B(n_2079),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_SL g4022 ( 
.A1(n_3730),
.A2(n_1063),
.B(n_1056),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3717),
.B(n_1064),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3885),
.A2(n_2265),
.B(n_2261),
.Y(n_4024)
);

NOR4xp25_ASAP7_75t_L g4025 ( 
.A(n_3822),
.B(n_1535),
.C(n_1539),
.D(n_1531),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3831),
.B(n_1540),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3890),
.A2(n_2269),
.B(n_2265),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3874),
.A2(n_2200),
.B(n_2079),
.Y(n_4028)
);

NAND3xp33_ASAP7_75t_L g4029 ( 
.A(n_3878),
.B(n_1066),
.C(n_1065),
.Y(n_4029)
);

INVx2_ASAP7_75t_SL g4030 ( 
.A(n_3700),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_L g4031 ( 
.A(n_3833),
.B(n_1067),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3847),
.B(n_1071),
.Y(n_4032)
);

OR2x2_ASAP7_75t_L g4033 ( 
.A(n_3789),
.B(n_1542),
.Y(n_4033)
);

OAI22xp5_ASAP7_75t_L g4034 ( 
.A1(n_3758),
.A2(n_1074),
.B1(n_1080),
.B2(n_1073),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_L g4035 ( 
.A(n_3743),
.B(n_1083),
.Y(n_4035)
);

BUFx12f_ASAP7_75t_L g4036 ( 
.A(n_3709),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3794),
.Y(n_4037)
);

AND2x4_ASAP7_75t_L g4038 ( 
.A(n_3719),
.B(n_471),
.Y(n_4038)
);

AOI21xp5_ASAP7_75t_L g4039 ( 
.A1(n_3713),
.A2(n_2288),
.B(n_2269),
.Y(n_4039)
);

OAI21x1_ASAP7_75t_L g4040 ( 
.A1(n_3832),
.A2(n_2288),
.B(n_2269),
.Y(n_4040)
);

OAI21x1_ASAP7_75t_L g4041 ( 
.A1(n_3834),
.A2(n_2297),
.B(n_2288),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_L g4042 ( 
.A(n_3821),
.B(n_1085),
.Y(n_4042)
);

OAI22xp5_ASAP7_75t_L g4043 ( 
.A1(n_3773),
.A2(n_1094),
.B1(n_1095),
.B2(n_1086),
.Y(n_4043)
);

OAI21x1_ASAP7_75t_L g4044 ( 
.A1(n_3915),
.A2(n_2305),
.B(n_2297),
.Y(n_4044)
);

BUFx3_ASAP7_75t_L g4045 ( 
.A(n_3744),
.Y(n_4045)
);

NAND2x1_ASAP7_75t_L g4046 ( 
.A(n_3861),
.B(n_2297),
.Y(n_4046)
);

INVx8_ASAP7_75t_L g4047 ( 
.A(n_3905),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3807),
.B(n_1098),
.Y(n_4048)
);

BUFx3_ASAP7_75t_L g4049 ( 
.A(n_3744),
.Y(n_4049)
);

AO31x2_ASAP7_75t_L g4050 ( 
.A1(n_3883),
.A2(n_1545),
.A3(n_1550),
.B(n_1543),
.Y(n_4050)
);

OAI21x1_ASAP7_75t_L g4051 ( 
.A1(n_3913),
.A2(n_2305),
.B(n_1552),
.Y(n_4051)
);

OR2x2_ASAP7_75t_L g4052 ( 
.A(n_3798),
.B(n_1551),
.Y(n_4052)
);

A2O1A1Ixp33_ASAP7_75t_L g4053 ( 
.A1(n_3836),
.A2(n_3784),
.B(n_3702),
.C(n_3899),
.Y(n_4053)
);

AO31x2_ASAP7_75t_L g4054 ( 
.A1(n_3757),
.A2(n_1556),
.A3(n_1558),
.B(n_1554),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3859),
.A2(n_2305),
.B(n_1560),
.Y(n_4055)
);

BUFx3_ASAP7_75t_L g4056 ( 
.A(n_3803),
.Y(n_4056)
);

AO31x2_ASAP7_75t_L g4057 ( 
.A1(n_3735),
.A2(n_3727),
.A3(n_3800),
.B(n_3781),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3736),
.B(n_1100),
.Y(n_4058)
);

CKINVDCx11_ASAP7_75t_R g4059 ( 
.A(n_3760),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3875),
.B(n_1559),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3857),
.A2(n_1564),
.B(n_1562),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3779),
.B(n_1101),
.Y(n_4062)
);

OAI21x1_ASAP7_75t_L g4063 ( 
.A1(n_3861),
.A2(n_1565),
.B(n_1470),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3809),
.B(n_3816),
.Y(n_4064)
);

INVx4_ASAP7_75t_L g4065 ( 
.A(n_3905),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3819),
.B(n_1110),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3813),
.B(n_1116),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3849),
.Y(n_4068)
);

INVx4_ASAP7_75t_L g4069 ( 
.A(n_3903),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_SL g4070 ( 
.A1(n_3842),
.A2(n_1127),
.B(n_1118),
.Y(n_4070)
);

OAI21x1_ASAP7_75t_L g4071 ( 
.A1(n_3864),
.A2(n_1470),
.B(n_1456),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_3752),
.B(n_1130),
.Y(n_4072)
);

OAI21xp5_ASAP7_75t_L g4073 ( 
.A1(n_3825),
.A2(n_1486),
.B(n_1476),
.Y(n_4073)
);

OAI21xp33_ASAP7_75t_L g4074 ( 
.A1(n_3773),
.A2(n_1135),
.B(n_1132),
.Y(n_4074)
);

CKINVDCx11_ASAP7_75t_R g4075 ( 
.A(n_3751),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_3713),
.A2(n_2243),
.B(n_2233),
.Y(n_4076)
);

A2O1A1Ixp33_ASAP7_75t_L g4077 ( 
.A1(n_3767),
.A2(n_1139),
.B(n_1138),
.C(n_1136),
.Y(n_4077)
);

INVx3_ASAP7_75t_L g4078 ( 
.A(n_3903),
.Y(n_4078)
);

OAI21x1_ASAP7_75t_L g4079 ( 
.A1(n_3864),
.A2(n_1486),
.B(n_1476),
.Y(n_4079)
);

OAI21x1_ASAP7_75t_L g4080 ( 
.A1(n_3888),
.A2(n_1523),
.B(n_1496),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_3889),
.B(n_472),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3713),
.A2(n_3856),
.B(n_3912),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3806),
.B(n_1141),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3893),
.B(n_479),
.Y(n_4084)
);

OAI21xp5_ASAP7_75t_L g4085 ( 
.A1(n_3795),
.A2(n_3868),
.B(n_3912),
.Y(n_4085)
);

NAND2xp33_ASAP7_75t_L g4086 ( 
.A(n_3699),
.B(n_1142),
.Y(n_4086)
);

BUFx3_ASAP7_75t_L g4087 ( 
.A(n_3709),
.Y(n_4087)
);

AOI21x1_ASAP7_75t_L g4088 ( 
.A1(n_3792),
.A2(n_1523),
.B(n_1496),
.Y(n_4088)
);

OAI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_3895),
.A2(n_1541),
.B(n_1536),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3815),
.B(n_1144),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3867),
.B(n_1808),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3775),
.Y(n_4092)
);

OAI21x1_ASAP7_75t_L g4093 ( 
.A1(n_3888),
.A2(n_1541),
.B(n_1536),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3876),
.Y(n_4094)
);

OAI21x1_ASAP7_75t_SL g4095 ( 
.A1(n_3881),
.A2(n_1563),
.B(n_1549),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3731),
.A2(n_2066),
.B(n_2028),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_SL g4097 ( 
.A(n_3762),
.B(n_2045),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3884),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3778),
.B(n_482),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3854),
.B(n_1808),
.Y(n_4100)
);

O2A1O1Ixp5_ASAP7_75t_L g4101 ( 
.A1(n_3707),
.A2(n_1563),
.B(n_1549),
.C(n_7),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_SL g4102 ( 
.A1(n_3826),
.A2(n_2056),
.B(n_2045),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_3871),
.B(n_1808),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3891),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3837),
.A2(n_1898),
.B(n_1808),
.Y(n_4105)
);

NOR4xp25_ASAP7_75t_L g4106 ( 
.A(n_3840),
.B(n_7),
.C(n_3),
.D(n_6),
.Y(n_4106)
);

OAI21x1_ASAP7_75t_L g4107 ( 
.A1(n_3837),
.A2(n_1898),
.B(n_2066),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3900),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3778),
.B(n_3790),
.Y(n_4109)
);

OAI21x1_ASAP7_75t_L g4110 ( 
.A1(n_3780),
.A2(n_1898),
.B(n_2066),
.Y(n_4110)
);

AND2x4_ASAP7_75t_L g4111 ( 
.A(n_3696),
.B(n_486),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3910),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3790),
.B(n_3),
.Y(n_4113)
);

OAI22xp5_ASAP7_75t_L g4114 ( 
.A1(n_3808),
.A2(n_10),
.B1(n_6),
.B2(n_9),
.Y(n_4114)
);

AOI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3750),
.A2(n_2056),
.B1(n_2113),
.B2(n_2045),
.Y(n_4115)
);

OAI21x1_ASAP7_75t_L g4116 ( 
.A1(n_3904),
.A2(n_2078),
.B(n_2066),
.Y(n_4116)
);

BUFx3_ASAP7_75t_L g4117 ( 
.A(n_3814),
.Y(n_4117)
);

OAI21x1_ASAP7_75t_L g4118 ( 
.A1(n_3812),
.A2(n_2078),
.B(n_2066),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3805),
.B(n_2045),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3766),
.Y(n_4120)
);

OAI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_3720),
.A2(n_2113),
.B1(n_2125),
.B2(n_2056),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3797),
.B(n_9),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3797),
.B(n_12),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3759),
.A2(n_3766),
.B(n_3771),
.Y(n_4124)
);

NAND2x1p5_ASAP7_75t_L g4125 ( 
.A(n_3696),
.B(n_2056),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3766),
.Y(n_4126)
);

AO31x2_ASAP7_75t_L g4127 ( 
.A1(n_3759),
.A2(n_492),
.A3(n_493),
.B(n_488),
.Y(n_4127)
);

BUFx6f_ASAP7_75t_L g4128 ( 
.A(n_3870),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_3698),
.B(n_13),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3759),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3698),
.B(n_15),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3850),
.Y(n_4132)
);

OAI21x1_ASAP7_75t_L g4133 ( 
.A1(n_3862),
.A2(n_2086),
.B(n_2078),
.Y(n_4133)
);

OAI21x1_ASAP7_75t_L g4134 ( 
.A1(n_3851),
.A2(n_2086),
.B(n_2078),
.Y(n_4134)
);

NOR2x1_ASAP7_75t_L g4135 ( 
.A(n_3910),
.B(n_2113),
.Y(n_4135)
);

AO32x2_ASAP7_75t_L g4136 ( 
.A1(n_3838),
.A2(n_19),
.A3(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_3771),
.A2(n_2086),
.B(n_2078),
.Y(n_4137)
);

INVx4_ASAP7_75t_L g4138 ( 
.A(n_3892),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_3771),
.A2(n_2150),
.B(n_2086),
.Y(n_4139)
);

OAI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_3866),
.A2(n_1752),
.B(n_1751),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3844),
.B(n_16),
.Y(n_4141)
);

OAI21x1_ASAP7_75t_L g4142 ( 
.A1(n_3902),
.A2(n_2150),
.B(n_2086),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3906),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3845),
.B(n_21),
.Y(n_4144)
);

OAI21x1_ASAP7_75t_L g4145 ( 
.A1(n_3911),
.A2(n_2168),
.B(n_2150),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3907),
.B(n_21),
.Y(n_4146)
);

OAI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3898),
.A2(n_1752),
.B(n_1751),
.Y(n_4147)
);

AOI21x1_ASAP7_75t_L g4148 ( 
.A1(n_3892),
.A2(n_2125),
.B(n_2113),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3827),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_3908),
.Y(n_4150)
);

OAI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3811),
.A2(n_1752),
.B(n_1751),
.Y(n_4151)
);

BUFx6f_ASAP7_75t_L g4152 ( 
.A(n_3839),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3796),
.B(n_498),
.Y(n_4153)
);

OAI21x1_ASAP7_75t_L g4154 ( 
.A1(n_3747),
.A2(n_2168),
.B(n_2150),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3830),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3814),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3924),
.Y(n_4157)
);

AOI21xp5_ASAP7_75t_L g4158 ( 
.A1(n_3958),
.A2(n_2168),
.B(n_2150),
.Y(n_4158)
);

INVxp67_ASAP7_75t_SL g4159 ( 
.A(n_3918),
.Y(n_4159)
);

AOI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_4140),
.A2(n_3920),
.B(n_4147),
.Y(n_4160)
);

NAND2x1p5_ASAP7_75t_L g4161 ( 
.A(n_4065),
.B(n_2125),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_4140),
.A2(n_2176),
.B(n_2168),
.Y(n_4162)
);

O2A1O1Ixp33_ASAP7_75t_L g4163 ( 
.A1(n_3961),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_4163)
);

OAI21x1_ASAP7_75t_L g4164 ( 
.A1(n_3933),
.A2(n_3930),
.B(n_3926),
.Y(n_4164)
);

INVx3_ASAP7_75t_L g4165 ( 
.A(n_4069),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4104),
.Y(n_4166)
);

INVx3_ASAP7_75t_L g4167 ( 
.A(n_4069),
.Y(n_4167)
);

BUFx2_ASAP7_75t_L g4168 ( 
.A(n_4010),
.Y(n_4168)
);

OAI22xp5_ASAP7_75t_L g4169 ( 
.A1(n_4006),
.A2(n_3782),
.B1(n_2127),
.B2(n_2189),
.Y(n_4169)
);

HB1xp67_ASAP7_75t_L g4170 ( 
.A(n_3985),
.Y(n_4170)
);

INVxp67_ASAP7_75t_L g4171 ( 
.A(n_4155),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3931),
.Y(n_4172)
);

CKINVDCx5p33_ASAP7_75t_R g4173 ( 
.A(n_4059),
.Y(n_4173)
);

INVx3_ASAP7_75t_L g4174 ( 
.A(n_3943),
.Y(n_4174)
);

BUFx6f_ASAP7_75t_L g4175 ( 
.A(n_3938),
.Y(n_4175)
);

NOR2xp33_ASAP7_75t_SL g4176 ( 
.A(n_4036),
.B(n_2125),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3934),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_3994),
.B(n_22),
.Y(n_4178)
);

CKINVDCx5p33_ASAP7_75t_R g4179 ( 
.A(n_3954),
.Y(n_4179)
);

BUFx2_ASAP7_75t_L g4180 ( 
.A(n_4000),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_3998),
.B(n_24),
.Y(n_4181)
);

INVx1_ASAP7_75t_SL g4182 ( 
.A(n_3959),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_3939),
.B(n_26),
.Y(n_4183)
);

AOI22xp33_ASAP7_75t_L g4184 ( 
.A1(n_3983),
.A2(n_2189),
.B1(n_2192),
.B2(n_2127),
.Y(n_4184)
);

O2A1O1Ixp5_ASAP7_75t_SL g4185 ( 
.A1(n_4114),
.A2(n_4097),
.B(n_4092),
.C(n_4120),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_3938),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_4068),
.B(n_27),
.Y(n_4187)
);

BUFx6f_ASAP7_75t_L g4188 ( 
.A(n_3938),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4108),
.Y(n_4189)
);

AND2x4_ASAP7_75t_L g4190 ( 
.A(n_3957),
.B(n_500),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_4132),
.B(n_27),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3963),
.Y(n_4192)
);

OAI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_4029),
.A2(n_2189),
.B1(n_2192),
.B2(n_2127),
.Y(n_4193)
);

AND2x4_ASAP7_75t_L g4194 ( 
.A(n_3980),
.B(n_3986),
.Y(n_4194)
);

INVx3_ASAP7_75t_L g4195 ( 
.A(n_3943),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4017),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4037),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3996),
.Y(n_4198)
);

OAI21xp33_ASAP7_75t_SL g4199 ( 
.A1(n_4106),
.A2(n_28),
.B(n_29),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_4005),
.B(n_28),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4094),
.Y(n_4201)
);

CKINVDCx11_ASAP7_75t_R g4202 ( 
.A(n_4087),
.Y(n_4202)
);

BUFx3_ASAP7_75t_L g4203 ( 
.A(n_4056),
.Y(n_4203)
);

AOI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_4029),
.A2(n_2189),
.B1(n_2192),
.B2(n_2127),
.Y(n_4204)
);

BUFx3_ASAP7_75t_L g4205 ( 
.A(n_3987),
.Y(n_4205)
);

AOI21xp5_ASAP7_75t_L g4206 ( 
.A1(n_4147),
.A2(n_2176),
.B(n_2168),
.Y(n_4206)
);

BUFx6f_ASAP7_75t_L g4207 ( 
.A(n_3943),
.Y(n_4207)
);

AOI21xp5_ASAP7_75t_L g4208 ( 
.A1(n_3976),
.A2(n_2222),
.B(n_2176),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4149),
.B(n_29),
.Y(n_4209)
);

OR2x2_ASAP7_75t_L g4210 ( 
.A(n_3941),
.B(n_30),
.Y(n_4210)
);

INVx2_ASAP7_75t_SL g4211 ( 
.A(n_4030),
.Y(n_4211)
);

INVx5_ASAP7_75t_L g4212 ( 
.A(n_4047),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_3970),
.B(n_501),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_4114),
.A2(n_2192),
.B1(n_2306),
.B2(n_2222),
.Y(n_4214)
);

AOI221xp5_ASAP7_75t_L g4215 ( 
.A1(n_4106),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.C(n_33),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4064),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_4143),
.B(n_32),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4130),
.Y(n_4218)
);

CKINVDCx5p33_ASAP7_75t_R g4219 ( 
.A(n_4011),
.Y(n_4219)
);

INVx1_ASAP7_75t_SL g4220 ( 
.A(n_4150),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4054),
.Y(n_4221)
);

INVx2_ASAP7_75t_L g4222 ( 
.A(n_4098),
.Y(n_4222)
);

INVx2_ASAP7_75t_SL g4223 ( 
.A(n_4128),
.Y(n_4223)
);

AND2x4_ASAP7_75t_L g4224 ( 
.A(n_4045),
.B(n_502),
.Y(n_4224)
);

O2A1O1Ixp33_ASAP7_75t_L g4225 ( 
.A1(n_4053),
.A2(n_38),
.B(n_34),
.C(n_35),
.Y(n_4225)
);

BUFx12f_ASAP7_75t_L g4226 ( 
.A(n_4150),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3944),
.B(n_34),
.Y(n_4227)
);

INVx4_ASAP7_75t_L g4228 ( 
.A(n_4047),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_3928),
.B(n_39),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_4035),
.B(n_41),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4033),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3919),
.B(n_41),
.Y(n_4232)
);

O2A1O1Ixp5_ASAP7_75t_L g4233 ( 
.A1(n_3992),
.A2(n_3978),
.B(n_4085),
.C(n_3925),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_4078),
.Y(n_4234)
);

AND2x4_ASAP7_75t_L g4235 ( 
.A(n_4049),
.B(n_503),
.Y(n_4235)
);

AOI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4150),
.A2(n_2306),
.B1(n_2222),
.B2(n_2227),
.Y(n_4236)
);

OAI22xp5_ASAP7_75t_L g4237 ( 
.A1(n_4144),
.A2(n_2306),
.B1(n_2222),
.B2(n_2227),
.Y(n_4237)
);

AO31x2_ASAP7_75t_L g4238 ( 
.A1(n_4082),
.A2(n_44),
.A3(n_42),
.B(n_43),
.Y(n_4238)
);

AND2x4_ASAP7_75t_L g4239 ( 
.A(n_3960),
.B(n_4138),
.Y(n_4239)
);

AND2x4_ASAP7_75t_L g4240 ( 
.A(n_3960),
.B(n_504),
.Y(n_4240)
);

INVx3_ASAP7_75t_L g4241 ( 
.A(n_4047),
.Y(n_4241)
);

NOR2xp33_ASAP7_75t_L g4242 ( 
.A(n_3936),
.B(n_44),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_4117),
.Y(n_4243)
);

AND2x4_ASAP7_75t_L g4244 ( 
.A(n_4138),
.B(n_509),
.Y(n_4244)
);

OR2x6_ASAP7_75t_L g4245 ( 
.A(n_4102),
.B(n_1698),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4112),
.B(n_45),
.Y(n_4246)
);

O2A1O1Ixp5_ASAP7_75t_L g4247 ( 
.A1(n_3992),
.A2(n_4085),
.B(n_3964),
.C(n_3982),
.Y(n_4247)
);

NOR3xp33_ASAP7_75t_L g4248 ( 
.A(n_4074),
.B(n_45),
.C(n_46),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_3948),
.B(n_47),
.Y(n_4249)
);

CKINVDCx20_ASAP7_75t_R g4250 ( 
.A(n_4075),
.Y(n_4250)
);

NOR2x1_ASAP7_75t_SL g4251 ( 
.A(n_3921),
.B(n_2306),
.Y(n_4251)
);

AND2x4_ASAP7_75t_L g4252 ( 
.A(n_4078),
.B(n_517),
.Y(n_4252)
);

BUFx12f_ASAP7_75t_L g4253 ( 
.A(n_4152),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4109),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_4019),
.A2(n_2222),
.B(n_2176),
.Y(n_4255)
);

AOI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_3955),
.A2(n_2227),
.B(n_2176),
.Y(n_4256)
);

CKINVDCx14_ASAP7_75t_R g4257 ( 
.A(n_4156),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_4152),
.B(n_47),
.Y(n_4258)
);

NAND2x1_ASAP7_75t_L g4259 ( 
.A(n_4065),
.B(n_2227),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4052),
.Y(n_4260)
);

NOR2xp67_ASAP7_75t_L g4261 ( 
.A(n_4026),
.B(n_48),
.Y(n_4261)
);

INVx2_ASAP7_75t_SL g4262 ( 
.A(n_4128),
.Y(n_4262)
);

O2A1O1Ixp33_ASAP7_75t_L g4263 ( 
.A1(n_4077),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4152),
.B(n_51),
.Y(n_4264)
);

INVx3_ASAP7_75t_L g4265 ( 
.A(n_4128),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4060),
.B(n_53),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3962),
.B(n_54),
.Y(n_4267)
);

HB1xp67_ASAP7_75t_L g4268 ( 
.A(n_4154),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_4153),
.B(n_56),
.Y(n_4269)
);

AND2x2_ASAP7_75t_L g4270 ( 
.A(n_4081),
.B(n_56),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3974),
.B(n_59),
.Y(n_4271)
);

INVx2_ASAP7_75t_SL g4272 ( 
.A(n_4111),
.Y(n_4272)
);

AOI22xp33_ASAP7_75t_L g4273 ( 
.A1(n_4074),
.A2(n_2233),
.B1(n_2243),
.B2(n_2227),
.Y(n_4273)
);

BUFx3_ASAP7_75t_L g4274 ( 
.A(n_4111),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4084),
.B(n_60),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_3942),
.A2(n_2243),
.B(n_2233),
.Y(n_4276)
);

INVx2_ASAP7_75t_SL g4277 ( 
.A(n_4099),
.Y(n_4277)
);

INVx1_ASAP7_75t_SL g4278 ( 
.A(n_3991),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3929),
.B(n_60),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4054),
.Y(n_4280)
);

BUFx12f_ASAP7_75t_L g4281 ( 
.A(n_3993),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4054),
.Y(n_4282)
);

AND2x6_ASAP7_75t_L g4283 ( 
.A(n_4038),
.B(n_2233),
.Y(n_4283)
);

AOI21xp5_ASAP7_75t_L g4284 ( 
.A1(n_3942),
.A2(n_2243),
.B(n_2233),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4136),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_3951),
.B(n_3984),
.Y(n_4286)
);

BUFx2_ASAP7_75t_L g4287 ( 
.A(n_4135),
.Y(n_4287)
);

A2O1A1Ixp33_ASAP7_75t_L g4288 ( 
.A1(n_3967),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_4288)
);

INVxp67_ASAP7_75t_SL g4289 ( 
.A(n_3997),
.Y(n_4289)
);

OA21x2_ASAP7_75t_L g4290 ( 
.A1(n_4007),
.A2(n_63),
.B(n_65),
.Y(n_4290)
);

HB1xp67_ASAP7_75t_L g4291 ( 
.A(n_4057),
.Y(n_4291)
);

BUFx6f_ASAP7_75t_L g4292 ( 
.A(n_4038),
.Y(n_4292)
);

AND2x4_ASAP7_75t_L g4293 ( 
.A(n_4135),
.B(n_519),
.Y(n_4293)
);

NOR2xp33_ASAP7_75t_L g4294 ( 
.A(n_4141),
.B(n_65),
.Y(n_4294)
);

O2A1O1Ixp33_ASAP7_75t_L g4295 ( 
.A1(n_4146),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_4295)
);

BUFx3_ASAP7_75t_L g4296 ( 
.A(n_4023),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4116),
.Y(n_4297)
);

AND2x2_ASAP7_75t_L g4298 ( 
.A(n_4113),
.B(n_68),
.Y(n_4298)
);

INVx2_ASAP7_75t_SL g4299 ( 
.A(n_4129),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_SL g4300 ( 
.A(n_3953),
.B(n_2243),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4122),
.B(n_70),
.Y(n_4301)
);

O2A1O1Ixp33_ASAP7_75t_SL g4302 ( 
.A1(n_4119),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_4131),
.Y(n_4303)
);

INVx2_ASAP7_75t_SL g4304 ( 
.A(n_4123),
.Y(n_4304)
);

BUFx6f_ASAP7_75t_L g4305 ( 
.A(n_4125),
.Y(n_4305)
);

O2A1O1Ixp33_ASAP7_75t_L g4306 ( 
.A1(n_3990),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_4306)
);

NAND2x1p5_ASAP7_75t_L g4307 ( 
.A(n_3940),
.B(n_4115),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_4151),
.A2(n_2259),
.B(n_2255),
.Y(n_4308)
);

INVx2_ASAP7_75t_SL g4309 ( 
.A(n_4046),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_L g4310 ( 
.A(n_3922),
.B(n_73),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3952),
.B(n_74),
.Y(n_4311)
);

INVx3_ASAP7_75t_L g4312 ( 
.A(n_4142),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4145),
.Y(n_4313)
);

INVx5_ASAP7_75t_L g4314 ( 
.A(n_3940),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4136),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_4151),
.A2(n_2259),
.B(n_2255),
.Y(n_4316)
);

BUFx2_ASAP7_75t_L g4317 ( 
.A(n_4134),
.Y(n_4317)
);

INVx3_ASAP7_75t_L g4318 ( 
.A(n_4133),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4136),
.Y(n_4319)
);

NOR2xp33_ASAP7_75t_L g4320 ( 
.A(n_4031),
.B(n_74),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_3950),
.Y(n_4321)
);

INVx2_ASAP7_75t_SL g4322 ( 
.A(n_4058),
.Y(n_4322)
);

INVx1_ASAP7_75t_SL g4323 ( 
.A(n_3972),
.Y(n_4323)
);

HB1xp67_ASAP7_75t_L g4324 ( 
.A(n_4057),
.Y(n_4324)
);

INVx4_ASAP7_75t_L g4325 ( 
.A(n_3950),
.Y(n_4325)
);

AND2x4_ASAP7_75t_L g4326 ( 
.A(n_3932),
.B(n_520),
.Y(n_4326)
);

AOI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_4096),
.A2(n_2259),
.B(n_2255),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3975),
.B(n_75),
.Y(n_4328)
);

AOI22xp5_ASAP7_75t_L g4329 ( 
.A1(n_4034),
.A2(n_2259),
.B1(n_2276),
.B2(n_2255),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_3949),
.B(n_77),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4057),
.B(n_77),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3927),
.B(n_78),
.Y(n_4332)
);

AOI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_3937),
.A2(n_2259),
.B(n_2255),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4008),
.A2(n_2284),
.B(n_2276),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_3927),
.B(n_78),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_4126),
.Y(n_4336)
);

AOI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_4008),
.A2(n_2284),
.B(n_2276),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4050),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_3990),
.B(n_79),
.Y(n_4339)
);

OR2x2_ASAP7_75t_L g4340 ( 
.A(n_4062),
.B(n_80),
.Y(n_4340)
);

OR2x2_ASAP7_75t_L g4341 ( 
.A(n_4066),
.B(n_80),
.Y(n_4341)
);

AOI22xp33_ASAP7_75t_L g4342 ( 
.A1(n_4072),
.A2(n_2284),
.B1(n_2276),
.B2(n_1713),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3995),
.B(n_4032),
.Y(n_4343)
);

AOI22xp33_ASAP7_75t_L g4344 ( 
.A1(n_3971),
.A2(n_2284),
.B1(n_2276),
.B2(n_1713),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_4050),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4115),
.B(n_81),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4050),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4042),
.B(n_4048),
.Y(n_4348)
);

A2O1A1Ixp33_ASAP7_75t_L g4349 ( 
.A1(n_3982),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_4349)
);

AND2x4_ASAP7_75t_L g4350 ( 
.A(n_3935),
.B(n_522),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4067),
.B(n_84),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4127),
.Y(n_4352)
);

INVx2_ASAP7_75t_L g4353 ( 
.A(n_4127),
.Y(n_4353)
);

INVx5_ASAP7_75t_L g4354 ( 
.A(n_4009),
.Y(n_4354)
);

INVx5_ASAP7_75t_L g4355 ( 
.A(n_3923),
.Y(n_4355)
);

OAI22xp33_ASAP7_75t_L g4356 ( 
.A1(n_4103),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_4356)
);

CKINVDCx6p67_ASAP7_75t_R g4357 ( 
.A(n_4083),
.Y(n_4357)
);

AOI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3965),
.A2(n_3956),
.B(n_3988),
.Y(n_4358)
);

OAI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_4101),
.A2(n_1752),
.B(n_1751),
.Y(n_4359)
);

NOR2xp33_ASAP7_75t_L g4360 ( 
.A(n_4090),
.B(n_85),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4091),
.B(n_4118),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3969),
.Y(n_4362)
);

BUFx6f_ASAP7_75t_L g4363 ( 
.A(n_4148),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4121),
.Y(n_4364)
);

AOI21xp5_ASAP7_75t_L g4365 ( 
.A1(n_3956),
.A2(n_2284),
.B(n_1713),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4127),
.Y(n_4366)
);

INVx2_ASAP7_75t_SL g4367 ( 
.A(n_4063),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3969),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_4086),
.B(n_88),
.Y(n_4369)
);

HB1xp67_ASAP7_75t_L g4370 ( 
.A(n_4044),
.Y(n_4370)
);

AND2x4_ASAP7_75t_L g4371 ( 
.A(n_4015),
.B(n_4021),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_L g4372 ( 
.A(n_4025),
.B(n_89),
.Y(n_4372)
);

OAI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_4043),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_4373)
);

INVxp67_ASAP7_75t_SL g4374 ( 
.A(n_4051),
.Y(n_4374)
);

AOI22xp33_ASAP7_75t_L g4375 ( 
.A1(n_4100),
.A2(n_1718),
.B1(n_1725),
.B2(n_1698),
.Y(n_4375)
);

A2O1A1Ixp33_ASAP7_75t_SL g4376 ( 
.A1(n_4022),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_4376)
);

AOI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_3966),
.A2(n_1718),
.B(n_1698),
.Y(n_4377)
);

INVx1_ASAP7_75t_SL g4378 ( 
.A(n_3979),
.Y(n_4378)
);

BUFx2_ASAP7_75t_L g4379 ( 
.A(n_4110),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4014),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4025),
.B(n_93),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4002),
.B(n_94),
.Y(n_4382)
);

BUFx12f_ASAP7_75t_L g4383 ( 
.A(n_4070),
.Y(n_4383)
);

CKINVDCx8_ASAP7_75t_R g4384 ( 
.A(n_4013),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_3977),
.B(n_95),
.Y(n_4385)
);

BUFx3_ASAP7_75t_L g4386 ( 
.A(n_4095),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_3968),
.Y(n_4387)
);

INVx3_ASAP7_75t_L g4388 ( 
.A(n_4040),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_4027),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4041),
.B(n_96),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_4124),
.B(n_96),
.Y(n_4391)
);

BUFx3_ASAP7_75t_L g4392 ( 
.A(n_4107),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3945),
.Y(n_4393)
);

CKINVDCx11_ASAP7_75t_R g4394 ( 
.A(n_4250),
.Y(n_4394)
);

OAI22xp5_ASAP7_75t_L g4395 ( 
.A1(n_4384),
.A2(n_3989),
.B1(n_3999),
.B2(n_4088),
.Y(n_4395)
);

BUFx2_ASAP7_75t_L g4396 ( 
.A(n_4180),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4157),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_SL g4398 ( 
.A1(n_4199),
.A2(n_4061),
.B1(n_4073),
.B2(n_4055),
.Y(n_4398)
);

BUFx6f_ASAP7_75t_L g4399 ( 
.A(n_4175),
.Y(n_4399)
);

BUFx10_ASAP7_75t_L g4400 ( 
.A(n_4173),
.Y(n_4400)
);

INVx4_ASAP7_75t_L g4401 ( 
.A(n_4212),
.Y(n_4401)
);

AOI22xp33_ASAP7_75t_L g4402 ( 
.A1(n_4248),
.A2(n_4073),
.B1(n_4089),
.B2(n_4024),
.Y(n_4402)
);

BUFx10_ASAP7_75t_L g4403 ( 
.A(n_4179),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4194),
.Y(n_4404)
);

OAI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_4349),
.A2(n_4039),
.B1(n_4076),
.B2(n_4137),
.Y(n_4405)
);

AOI21xp5_ASAP7_75t_L g4406 ( 
.A1(n_4160),
.A2(n_4139),
.B(n_4089),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4172),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4177),
.Y(n_4408)
);

HB1xp67_ASAP7_75t_L g4409 ( 
.A(n_4159),
.Y(n_4409)
);

OAI22xp5_ASAP7_75t_L g4410 ( 
.A1(n_4288),
.A2(n_4016),
.B1(n_4105),
.B2(n_101),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4194),
.Y(n_4411)
);

BUFx3_ASAP7_75t_L g4412 ( 
.A(n_4226),
.Y(n_4412)
);

AOI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_4229),
.A2(n_3947),
.B1(n_4079),
.B2(n_4071),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_4215),
.A2(n_4093),
.B1(n_4080),
.B2(n_4004),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4192),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4197),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4166),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4196),
.Y(n_4418)
);

AOI22xp5_ASAP7_75t_L g4419 ( 
.A1(n_4242),
.A2(n_4020),
.B1(n_4003),
.B2(n_4018),
.Y(n_4419)
);

INVxp67_ASAP7_75t_L g4420 ( 
.A(n_4170),
.Y(n_4420)
);

AOI22xp33_ASAP7_75t_L g4421 ( 
.A1(n_4369),
.A2(n_4028),
.B1(n_4012),
.B2(n_3981),
.Y(n_4421)
);

CKINVDCx20_ASAP7_75t_R g4422 ( 
.A(n_4202),
.Y(n_4422)
);

OAI22xp5_ASAP7_75t_SL g4423 ( 
.A1(n_4257),
.A2(n_4219),
.B1(n_4294),
.B2(n_4339),
.Y(n_4423)
);

INVx6_ASAP7_75t_L g4424 ( 
.A(n_4253),
.Y(n_4424)
);

AOI22xp33_ASAP7_75t_L g4425 ( 
.A1(n_4281),
.A2(n_4360),
.B1(n_4320),
.B2(n_4357),
.Y(n_4425)
);

CKINVDCx14_ASAP7_75t_R g4426 ( 
.A(n_4243),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4189),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4162),
.A2(n_3973),
.B(n_4001),
.Y(n_4428)
);

CKINVDCx20_ASAP7_75t_R g4429 ( 
.A(n_4205),
.Y(n_4429)
);

INVx1_ASAP7_75t_SL g4430 ( 
.A(n_4220),
.Y(n_4430)
);

AOI22xp33_ASAP7_75t_SL g4431 ( 
.A1(n_4331),
.A2(n_3946),
.B1(n_102),
.B2(n_97),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_L g4432 ( 
.A1(n_4184),
.A2(n_103),
.B1(n_97),
.B2(n_98),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4198),
.Y(n_4433)
);

BUFx2_ASAP7_75t_L g4434 ( 
.A(n_4168),
.Y(n_4434)
);

AOI22xp33_ASAP7_75t_L g4435 ( 
.A1(n_4303),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4254),
.Y(n_4436)
);

CKINVDCx6p67_ASAP7_75t_R g4437 ( 
.A(n_4203),
.Y(n_4437)
);

BUFx2_ASAP7_75t_L g4438 ( 
.A(n_4303),
.Y(n_4438)
);

INVx4_ASAP7_75t_L g4439 ( 
.A(n_4212),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_4175),
.Y(n_4440)
);

OAI22xp5_ASAP7_75t_L g4441 ( 
.A1(n_4214),
.A2(n_109),
.B1(n_104),
.B2(n_106),
.Y(n_4441)
);

INVxp67_ASAP7_75t_SL g4442 ( 
.A(n_4291),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4216),
.Y(n_4443)
);

CKINVDCx5p33_ASAP7_75t_R g4444 ( 
.A(n_4175),
.Y(n_4444)
);

BUFx3_ASAP7_75t_L g4445 ( 
.A(n_4186),
.Y(n_4445)
);

CKINVDCx20_ASAP7_75t_R g4446 ( 
.A(n_4296),
.Y(n_4446)
);

AOI22xp33_ASAP7_75t_SL g4447 ( 
.A1(n_4292),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4201),
.Y(n_4448)
);

OAI22xp33_ASAP7_75t_L g4449 ( 
.A1(n_4381),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_4449)
);

INVx2_ASAP7_75t_SL g4450 ( 
.A(n_4186),
.Y(n_4450)
);

AOI22xp33_ASAP7_75t_L g4451 ( 
.A1(n_4303),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4171),
.B(n_116),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4299),
.B(n_116),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4222),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4218),
.Y(n_4455)
);

INVx8_ASAP7_75t_L g4456 ( 
.A(n_4213),
.Y(n_4456)
);

AOI22xp33_ASAP7_75t_SL g4457 ( 
.A1(n_4292),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_4457)
);

INVx6_ASAP7_75t_L g4458 ( 
.A(n_4186),
.Y(n_4458)
);

INVx1_ASAP7_75t_SL g4459 ( 
.A(n_4278),
.Y(n_4459)
);

BUFx12f_ASAP7_75t_L g4460 ( 
.A(n_4383),
.Y(n_4460)
);

INVx3_ASAP7_75t_L g4461 ( 
.A(n_4188),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_4310),
.A2(n_121),
.B1(n_117),
.B2(n_120),
.Y(n_4462)
);

BUFx6f_ASAP7_75t_L g4463 ( 
.A(n_4188),
.Y(n_4463)
);

AOI22xp33_ASAP7_75t_SL g4464 ( 
.A1(n_4292),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_4464)
);

INVx1_ASAP7_75t_SL g4465 ( 
.A(n_4182),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4218),
.Y(n_4466)
);

INVx1_ASAP7_75t_SL g4467 ( 
.A(n_4188),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4260),
.Y(n_4468)
);

CKINVDCx11_ASAP7_75t_R g4469 ( 
.A(n_4323),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_4211),
.Y(n_4470)
);

AOI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4169),
.A2(n_1725),
.B1(n_1726),
.B2(n_1718),
.Y(n_4471)
);

OAI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_4225),
.A2(n_125),
.B1(n_122),
.B2(n_124),
.Y(n_4472)
);

OAI22xp33_ASAP7_75t_L g4473 ( 
.A1(n_4372),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_4473)
);

INVx4_ASAP7_75t_L g4474 ( 
.A(n_4212),
.Y(n_4474)
);

OAI22xp33_ASAP7_75t_SL g4475 ( 
.A1(n_4391),
.A2(n_129),
.B1(n_126),
.B2(n_127),
.Y(n_4475)
);

INVx3_ASAP7_75t_L g4476 ( 
.A(n_4239),
.Y(n_4476)
);

BUFx6f_ASAP7_75t_L g4477 ( 
.A(n_4207),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4336),
.Y(n_4478)
);

CKINVDCx11_ASAP7_75t_R g4479 ( 
.A(n_4207),
.Y(n_4479)
);

INVx1_ASAP7_75t_SL g4480 ( 
.A(n_4322),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_4385),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_4481)
);

CKINVDCx20_ASAP7_75t_R g4482 ( 
.A(n_4274),
.Y(n_4482)
);

CKINVDCx11_ASAP7_75t_R g4483 ( 
.A(n_4207),
.Y(n_4483)
);

OAI21xp33_ASAP7_75t_L g4484 ( 
.A1(n_4295),
.A2(n_4373),
.B(n_4306),
.Y(n_4484)
);

INVx6_ASAP7_75t_L g4485 ( 
.A(n_4228),
.Y(n_4485)
);

BUFx2_ASAP7_75t_L g4486 ( 
.A(n_4239),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4336),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4234),
.Y(n_4488)
);

AOI22xp33_ASAP7_75t_L g4489 ( 
.A1(n_4380),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_4489)
);

AOI22xp33_ASAP7_75t_L g4490 ( 
.A1(n_4269),
.A2(n_136),
.B1(n_132),
.B2(n_133),
.Y(n_4490)
);

BUFx2_ASAP7_75t_R g4491 ( 
.A(n_4286),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4231),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4324),
.Y(n_4493)
);

INVx6_ASAP7_75t_L g4494 ( 
.A(n_4228),
.Y(n_4494)
);

OAI21xp33_ASAP7_75t_L g4495 ( 
.A1(n_4163),
.A2(n_133),
.B(n_136),
.Y(n_4495)
);

OAI22x1_ASAP7_75t_L g4496 ( 
.A1(n_4285),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_4496)
);

OAI22xp5_ASAP7_75t_L g4497 ( 
.A1(n_4289),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_4497)
);

AOI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4283),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_4265),
.Y(n_4499)
);

INVx3_ASAP7_75t_L g4500 ( 
.A(n_4265),
.Y(n_4500)
);

INVx3_ASAP7_75t_L g4501 ( 
.A(n_4165),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_SL g4502 ( 
.A1(n_4343),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4502)
);

CKINVDCx11_ASAP7_75t_R g4503 ( 
.A(n_4305),
.Y(n_4503)
);

INVx2_ASAP7_75t_SL g4504 ( 
.A(n_4223),
.Y(n_4504)
);

BUFx2_ASAP7_75t_L g4505 ( 
.A(n_4241),
.Y(n_4505)
);

BUFx12f_ASAP7_75t_L g4506 ( 
.A(n_4210),
.Y(n_4506)
);

INVx2_ASAP7_75t_SL g4507 ( 
.A(n_4262),
.Y(n_4507)
);

INVx8_ASAP7_75t_L g4508 ( 
.A(n_4213),
.Y(n_4508)
);

INVx5_ASAP7_75t_L g4509 ( 
.A(n_4245),
.Y(n_4509)
);

AOI22xp33_ASAP7_75t_L g4510 ( 
.A1(n_4283),
.A2(n_149),
.B1(n_145),
.B2(n_146),
.Y(n_4510)
);

OAI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_4300),
.A2(n_149),
.B1(n_145),
.B2(n_146),
.Y(n_4511)
);

NAND2x1p5_ASAP7_75t_L g4512 ( 
.A(n_4314),
.B(n_1725),
.Y(n_4512)
);

AND2x2_ASAP7_75t_L g4513 ( 
.A(n_4304),
.B(n_151),
.Y(n_4513)
);

BUFx2_ASAP7_75t_L g4514 ( 
.A(n_4241),
.Y(n_4514)
);

AOI22xp33_ASAP7_75t_L g4515 ( 
.A1(n_4283),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_4515)
);

BUFx10_ASAP7_75t_L g4516 ( 
.A(n_4240),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_L g4517 ( 
.A1(n_4283),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_4517)
);

NAND2x1p5_ASAP7_75t_L g4518 ( 
.A(n_4314),
.B(n_1726),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4287),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4221),
.Y(n_4520)
);

AOI22xp33_ASAP7_75t_L g4521 ( 
.A1(n_4348),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_4174),
.Y(n_4522)
);

INVx8_ASAP7_75t_L g4523 ( 
.A(n_4240),
.Y(n_4523)
);

BUFx10_ASAP7_75t_L g4524 ( 
.A(n_4244),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4313),
.Y(n_4525)
);

AOI22xp33_ASAP7_75t_SL g4526 ( 
.A1(n_4346),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4526)
);

CKINVDCx5p33_ASAP7_75t_R g4527 ( 
.A(n_4174),
.Y(n_4527)
);

CKINVDCx5p33_ASAP7_75t_R g4528 ( 
.A(n_4195),
.Y(n_4528)
);

OAI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4307),
.A2(n_162),
.B1(n_158),
.B2(n_160),
.Y(n_4529)
);

AOI22xp33_ASAP7_75t_SL g4530 ( 
.A1(n_4290),
.A2(n_163),
.B1(n_160),
.B2(n_162),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4297),
.Y(n_4531)
);

AOI22xp33_ASAP7_75t_SL g4532 ( 
.A1(n_4290),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_4532)
);

INVx4_ASAP7_75t_L g4533 ( 
.A(n_4314),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_SL g4534 ( 
.A1(n_4332),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4312),
.Y(n_4535)
);

INVx6_ASAP7_75t_L g4536 ( 
.A(n_4258),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4221),
.Y(n_4537)
);

INVx3_ASAP7_75t_L g4538 ( 
.A(n_4165),
.Y(n_4538)
);

BUFx6f_ASAP7_75t_L g4539 ( 
.A(n_4195),
.Y(n_4539)
);

BUFx2_ASAP7_75t_SL g4540 ( 
.A(n_4261),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4282),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4238),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_SL g4543 ( 
.A1(n_4335),
.A2(n_169),
.B1(n_166),
.B2(n_167),
.Y(n_4543)
);

BUFx2_ASAP7_75t_L g4544 ( 
.A(n_4167),
.Y(n_4544)
);

BUFx8_ASAP7_75t_L g4545 ( 
.A(n_4264),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4312),
.Y(n_4546)
);

OAI22xp33_ASAP7_75t_L g4547 ( 
.A1(n_4329),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_4547)
);

INVx8_ASAP7_75t_L g4548 ( 
.A(n_4244),
.Y(n_4548)
);

OAI22xp33_ASAP7_75t_L g4549 ( 
.A1(n_4315),
.A2(n_4319),
.B1(n_4176),
.B2(n_4272),
.Y(n_4549)
);

AOI22xp33_ASAP7_75t_L g4550 ( 
.A1(n_4382),
.A2(n_4301),
.B1(n_4298),
.B2(n_4386),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_4167),
.Y(n_4551)
);

INVx6_ASAP7_75t_L g4552 ( 
.A(n_4224),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4238),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_4356),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_4554)
);

AOI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4389),
.A2(n_1730),
.B1(n_1726),
.B2(n_175),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4277),
.B(n_173),
.Y(n_4556)
);

BUFx8_ASAP7_75t_SL g4557 ( 
.A(n_4181),
.Y(n_4557)
);

OAI22xp33_ASAP7_75t_L g4558 ( 
.A1(n_4230),
.A2(n_4209),
.B1(n_4279),
.B2(n_4191),
.Y(n_4558)
);

AOI22xp33_ASAP7_75t_L g4559 ( 
.A1(n_4270),
.A2(n_179),
.B1(n_174),
.B2(n_176),
.Y(n_4559)
);

CKINVDCx20_ASAP7_75t_R g4560 ( 
.A(n_4275),
.Y(n_4560)
);

CKINVDCx20_ASAP7_75t_R g4561 ( 
.A(n_4232),
.Y(n_4561)
);

INVx2_ASAP7_75t_L g4562 ( 
.A(n_4268),
.Y(n_4562)
);

AOI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_4190),
.A2(n_1730),
.B1(n_181),
.B2(n_179),
.Y(n_4563)
);

INVx11_ASAP7_75t_L g4564 ( 
.A(n_4246),
.Y(n_4564)
);

INVx2_ASAP7_75t_L g4565 ( 
.A(n_4280),
.Y(n_4565)
);

INVx2_ASAP7_75t_SL g4566 ( 
.A(n_4305),
.Y(n_4566)
);

CKINVDCx5p33_ASAP7_75t_R g4567 ( 
.A(n_4266),
.Y(n_4567)
);

BUFx12f_ASAP7_75t_L g4568 ( 
.A(n_4340),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4238),
.Y(n_4569)
);

OAI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4263),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4317),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4190),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_4572)
);

CKINVDCx5p33_ASAP7_75t_R g4573 ( 
.A(n_4351),
.Y(n_4573)
);

AOI22xp5_ASAP7_75t_L g4574 ( 
.A1(n_4224),
.A2(n_1730),
.B1(n_187),
.B2(n_183),
.Y(n_4574)
);

OAI22xp5_ASAP7_75t_L g4575 ( 
.A1(n_4273),
.A2(n_188),
.B1(n_184),
.B2(n_187),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4361),
.B(n_188),
.Y(n_4576)
);

BUFx3_ASAP7_75t_L g4577 ( 
.A(n_4235),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4486),
.B(n_4434),
.Y(n_4578)
);

INVxp33_ASAP7_75t_L g4579 ( 
.A(n_4394),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4455),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4455),
.Y(n_4581)
);

O2A1O1Ixp33_ASAP7_75t_L g4582 ( 
.A1(n_4475),
.A2(n_4484),
.B(n_4472),
.C(n_4473),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4420),
.B(n_4378),
.Y(n_4583)
);

INVx2_ASAP7_75t_L g4584 ( 
.A(n_4519),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_4409),
.Y(n_4585)
);

HB1xp67_ASAP7_75t_L g4586 ( 
.A(n_4571),
.Y(n_4586)
);

AOI21x1_ASAP7_75t_SL g4587 ( 
.A1(n_4576),
.A2(n_4330),
.B(n_4178),
.Y(n_4587)
);

OR2x2_ASAP7_75t_L g4588 ( 
.A(n_4404),
.B(n_4338),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4466),
.Y(n_4589)
);

OR2x2_ASAP7_75t_L g4590 ( 
.A(n_4411),
.B(n_4345),
.Y(n_4590)
);

OR2x2_ASAP7_75t_L g4591 ( 
.A(n_4396),
.B(n_4352),
.Y(n_4591)
);

CKINVDCx16_ASAP7_75t_R g4592 ( 
.A(n_4422),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4478),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_4438),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4487),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4443),
.B(n_4364),
.Y(n_4596)
);

OAI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4534),
.A2(n_4204),
.B1(n_4333),
.B2(n_4236),
.Y(n_4597)
);

CKINVDCx5p33_ASAP7_75t_R g4598 ( 
.A(n_4469),
.Y(n_4598)
);

INVx3_ASAP7_75t_L g4599 ( 
.A(n_4476),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4468),
.B(n_4390),
.Y(n_4600)
);

OAI22xp5_ASAP7_75t_L g4601 ( 
.A1(n_4543),
.A2(n_4510),
.B1(n_4515),
.B2(n_4498),
.Y(n_4601)
);

AND2x2_ASAP7_75t_L g4602 ( 
.A(n_4476),
.B(n_4370),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4544),
.B(n_4379),
.Y(n_4603)
);

AND2x4_ASAP7_75t_L g4604 ( 
.A(n_4501),
.B(n_4318),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4397),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4407),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4436),
.B(n_4217),
.Y(n_4607)
);

AOI221xp5_ASAP7_75t_L g4608 ( 
.A1(n_4502),
.A2(n_4233),
.B1(n_4247),
.B2(n_4249),
.C(n_4267),
.Y(n_4608)
);

NOR2xp67_ASAP7_75t_R g4609 ( 
.A(n_4401),
.B(n_4355),
.Y(n_4609)
);

OR2x2_ASAP7_75t_L g4610 ( 
.A(n_4492),
.B(n_4353),
.Y(n_4610)
);

OA21x2_ASAP7_75t_L g4611 ( 
.A1(n_4542),
.A2(n_4366),
.B(n_4164),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_4459),
.Y(n_4612)
);

AOI21xp5_ASAP7_75t_L g4613 ( 
.A1(n_4406),
.A2(n_4206),
.B(n_4334),
.Y(n_4613)
);

AOI21xp33_ASAP7_75t_L g4614 ( 
.A1(n_4558),
.A2(n_4341),
.B(n_4311),
.Y(n_4614)
);

BUFx2_ASAP7_75t_L g4615 ( 
.A(n_4522),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4499),
.B(n_4183),
.Y(n_4616)
);

OA22x2_ASAP7_75t_L g4617 ( 
.A1(n_4496),
.A2(n_4187),
.B1(n_4227),
.B2(n_4271),
.Y(n_4617)
);

O2A1O1Ixp5_ASAP7_75t_L g4618 ( 
.A1(n_4449),
.A2(n_4570),
.B(n_4481),
.C(n_4549),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4505),
.B(n_4355),
.Y(n_4619)
);

OR2x2_ASAP7_75t_L g4620 ( 
.A(n_4427),
.B(n_4347),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4408),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4514),
.B(n_4355),
.Y(n_4622)
);

BUFx6f_ASAP7_75t_L g4623 ( 
.A(n_4503),
.Y(n_4623)
);

INVx2_ASAP7_75t_L g4624 ( 
.A(n_4415),
.Y(n_4624)
);

AOI21x1_ASAP7_75t_SL g4625 ( 
.A1(n_4453),
.A2(n_4328),
.B(n_4200),
.Y(n_4625)
);

BUFx4f_ASAP7_75t_L g4626 ( 
.A(n_4460),
.Y(n_4626)
);

OA21x2_ASAP7_75t_L g4627 ( 
.A1(n_4553),
.A2(n_4208),
.B(n_4158),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4418),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4448),
.B(n_4362),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4430),
.B(n_4392),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4433),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4520),
.Y(n_4632)
);

OR2x2_ASAP7_75t_L g4633 ( 
.A(n_4562),
.B(n_4368),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4537),
.Y(n_4634)
);

O2A1O1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4495),
.A2(n_4376),
.B(n_4302),
.C(n_4237),
.Y(n_4635)
);

AOI21x1_ASAP7_75t_SL g4636 ( 
.A1(n_4452),
.A2(n_4350),
.B(n_4326),
.Y(n_4636)
);

NOR2xp67_ASAP7_75t_L g4637 ( 
.A(n_4533),
.B(n_4325),
.Y(n_4637)
);

OAI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4517),
.A2(n_4245),
.B1(n_4293),
.B2(n_4342),
.Y(n_4638)
);

O2A1O1Ixp33_ASAP7_75t_L g4639 ( 
.A1(n_4529),
.A2(n_4358),
.B(n_4193),
.C(n_4365),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4541),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4416),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4417),
.Y(n_4642)
);

AOI221x1_ASAP7_75t_SL g4643 ( 
.A1(n_4497),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.C(n_194),
.Y(n_4643)
);

INVx2_ASAP7_75t_L g4644 ( 
.A(n_4488),
.Y(n_4644)
);

NOR2xp33_ASAP7_75t_SL g4645 ( 
.A(n_4491),
.B(n_4308),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4480),
.B(n_4318),
.Y(n_4646)
);

AOI21xp5_ASAP7_75t_L g4647 ( 
.A1(n_4410),
.A2(n_4337),
.B(n_4316),
.Y(n_4647)
);

O2A1O1Ixp33_ASAP7_75t_L g4648 ( 
.A1(n_4547),
.A2(n_4284),
.B(n_4276),
.C(n_4359),
.Y(n_4648)
);

OA21x2_ASAP7_75t_L g4649 ( 
.A1(n_4569),
.A2(n_4327),
.B(n_4256),
.Y(n_4649)
);

AOI21xp5_ASAP7_75t_L g4650 ( 
.A1(n_4395),
.A2(n_4402),
.B(n_4405),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4454),
.B(n_4551),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4493),
.Y(n_4652)
);

OA21x2_ASAP7_75t_L g4653 ( 
.A1(n_4535),
.A2(n_4321),
.B(n_4377),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4465),
.B(n_4501),
.Y(n_4654)
);

AND2x2_ASAP7_75t_L g4655 ( 
.A(n_4538),
.B(n_4536),
.Y(n_4655)
);

BUFx4f_ASAP7_75t_SL g4656 ( 
.A(n_4429),
.Y(n_4656)
);

INVx2_ASAP7_75t_SL g4657 ( 
.A(n_4424),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4538),
.B(n_4325),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4536),
.B(n_4388),
.Y(n_4659)
);

NAND2xp5_ASAP7_75t_L g4660 ( 
.A(n_4550),
.B(n_4350),
.Y(n_4660)
);

OA21x2_ASAP7_75t_L g4661 ( 
.A1(n_4546),
.A2(n_4374),
.B(n_4393),
.Y(n_4661)
);

OA21x2_ASAP7_75t_L g4662 ( 
.A1(n_4442),
.A2(n_4393),
.B(n_4255),
.Y(n_4662)
);

AOI21xp5_ASAP7_75t_SL g4663 ( 
.A1(n_4401),
.A2(n_4326),
.B(n_4293),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4437),
.B(n_4388),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4525),
.Y(n_4665)
);

AND2x4_ASAP7_75t_L g4666 ( 
.A(n_4500),
.B(n_4309),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4531),
.Y(n_4667)
);

OAI22xp5_ASAP7_75t_L g4668 ( 
.A1(n_4530),
.A2(n_4354),
.B1(n_4344),
.B2(n_4235),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4426),
.B(n_4251),
.Y(n_4669)
);

OAI22xp5_ASAP7_75t_L g4670 ( 
.A1(n_4532),
.A2(n_4354),
.B1(n_4305),
.B2(n_4161),
.Y(n_4670)
);

AOI21x1_ASAP7_75t_SL g4671 ( 
.A1(n_4513),
.A2(n_4252),
.B(n_4371),
.Y(n_4671)
);

O2A1O1Ixp5_ASAP7_75t_L g4672 ( 
.A1(n_4533),
.A2(n_4259),
.B(n_4252),
.C(n_4387),
.Y(n_4672)
);

INVx1_ASAP7_75t_SL g4673 ( 
.A(n_4458),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4412),
.B(n_4251),
.Y(n_4674)
);

NAND4xp25_ASAP7_75t_L g4675 ( 
.A(n_4462),
.B(n_4375),
.C(n_196),
.D(n_191),
.Y(n_4675)
);

AND2x4_ASAP7_75t_L g4676 ( 
.A(n_4500),
.B(n_4371),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4467),
.B(n_4185),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4565),
.Y(n_4678)
);

AOI21x1_ASAP7_75t_SL g4679 ( 
.A1(n_4556),
.A2(n_4354),
.B(n_195),
.Y(n_4679)
);

A2O1A1Ixp33_ASAP7_75t_L g4680 ( 
.A1(n_4555),
.A2(n_4367),
.B(n_197),
.C(n_195),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4539),
.Y(n_4681)
);

OR2x2_ASAP7_75t_L g4682 ( 
.A(n_4504),
.B(n_4363),
.Y(n_4682)
);

CKINVDCx5p33_ASAP7_75t_R g4683 ( 
.A(n_4479),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4554),
.A2(n_4363),
.B1(n_198),
.B2(n_196),
.Y(n_4684)
);

O2A1O1Ixp5_ASAP7_75t_L g4685 ( 
.A1(n_4511),
.A2(n_199),
.B(n_197),
.C(n_198),
.Y(n_4685)
);

OAI211xp5_ASAP7_75t_L g4686 ( 
.A1(n_4526),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4507),
.B(n_4363),
.Y(n_4687)
);

OAI22xp5_ASAP7_75t_L g4688 ( 
.A1(n_4563),
.A2(n_205),
.B1(n_200),
.B2(n_202),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4461),
.B(n_205),
.Y(n_4689)
);

A2O1A1Ixp33_ASAP7_75t_SL g4690 ( 
.A1(n_4521),
.A2(n_209),
.B(n_206),
.C(n_207),
.Y(n_4690)
);

OR2x2_ASAP7_75t_L g4691 ( 
.A(n_4461),
.B(n_206),
.Y(n_4691)
);

OR2x2_ASAP7_75t_L g4692 ( 
.A(n_4450),
.B(n_4566),
.Y(n_4692)
);

OAI22xp5_ASAP7_75t_L g4693 ( 
.A1(n_4574),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_4693)
);

OR2x2_ASAP7_75t_L g4694 ( 
.A(n_4440),
.B(n_211),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4539),
.Y(n_4695)
);

HB1xp67_ASAP7_75t_L g4696 ( 
.A(n_4539),
.Y(n_4696)
);

CKINVDCx20_ASAP7_75t_R g4697 ( 
.A(n_4446),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4445),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_4483),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4458),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4527),
.B(n_213),
.Y(n_4701)
);

AOI211xp5_ASAP7_75t_L g4702 ( 
.A1(n_4423),
.A2(n_216),
.B(n_213),
.C(n_215),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_4573),
.B(n_216),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4399),
.B(n_219),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4528),
.B(n_220),
.Y(n_4705)
);

AOI21x1_ASAP7_75t_SL g4706 ( 
.A1(n_4540),
.A2(n_221),
.B(n_222),
.Y(n_4706)
);

OR2x2_ASAP7_75t_L g4707 ( 
.A(n_4577),
.B(n_222),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4399),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4482),
.B(n_223),
.Y(n_4709)
);

OAI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4447),
.A2(n_228),
.B1(n_225),
.B2(n_226),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4399),
.B(n_225),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4398),
.A2(n_1764),
.B(n_524),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4463),
.Y(n_4713)
);

NAND2xp5_ASAP7_75t_L g4714 ( 
.A(n_4463),
.B(n_4425),
.Y(n_4714)
);

AOI21x1_ASAP7_75t_SL g4715 ( 
.A1(n_4400),
.A2(n_228),
.B(n_229),
.Y(n_4715)
);

AOI21x1_ASAP7_75t_SL g4716 ( 
.A1(n_4400),
.A2(n_229),
.B(n_230),
.Y(n_4716)
);

AOI21xp5_ASAP7_75t_SL g4717 ( 
.A1(n_4439),
.A2(n_230),
.B(n_231),
.Y(n_4717)
);

O2A1O1Ixp33_ASAP7_75t_L g4718 ( 
.A1(n_4432),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4568),
.B(n_234),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_SL g4720 ( 
.A1(n_4439),
.A2(n_236),
.B(n_237),
.Y(n_4720)
);

NAND2x1_ASAP7_75t_L g4721 ( 
.A(n_4615),
.B(n_4474),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4632),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4596),
.B(n_4419),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4578),
.B(n_4444),
.Y(n_4724)
);

INVx2_ASAP7_75t_SL g4725 ( 
.A(n_4623),
.Y(n_4725)
);

INVx1_ASAP7_75t_SL g4726 ( 
.A(n_4656),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_4592),
.Y(n_4727)
);

AND2x4_ASAP7_75t_L g4728 ( 
.A(n_4664),
.B(n_4474),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4585),
.B(n_4463),
.Y(n_4729)
);

XNOR2xp5_ASAP7_75t_L g4730 ( 
.A(n_4697),
.B(n_4560),
.Y(n_4730)
);

OR2x6_ASAP7_75t_L g4731 ( 
.A(n_4663),
.B(n_4456),
.Y(n_4731)
);

NOR3xp33_ASAP7_75t_SL g4732 ( 
.A(n_4683),
.B(n_4470),
.C(n_4567),
.Y(n_4732)
);

INVx8_ASAP7_75t_L g4733 ( 
.A(n_4623),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4580),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4581),
.Y(n_4735)
);

INVx1_ASAP7_75t_L g4736 ( 
.A(n_4634),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4640),
.Y(n_4737)
);

OAI21xp5_ASAP7_75t_L g4738 ( 
.A1(n_4650),
.A2(n_4431),
.B(n_4457),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4589),
.Y(n_4739)
);

OAI22xp5_ASAP7_75t_L g4740 ( 
.A1(n_4702),
.A2(n_4552),
.B1(n_4471),
.B2(n_4572),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_L g4741 ( 
.A1(n_4601),
.A2(n_4506),
.B1(n_4464),
.B2(n_4575),
.Y(n_4741)
);

AND2x2_ASAP7_75t_L g4742 ( 
.A(n_4655),
.B(n_4424),
.Y(n_4742)
);

NAND2xp33_ASAP7_75t_R g4743 ( 
.A(n_4598),
.B(n_4699),
.Y(n_4743)
);

AOI22xp33_ASAP7_75t_L g4744 ( 
.A1(n_4608),
.A2(n_4490),
.B1(n_4489),
.B2(n_4561),
.Y(n_4744)
);

BUFx6f_ASAP7_75t_SL g4745 ( 
.A(n_4623),
.Y(n_4745)
);

INVx3_ASAP7_75t_L g4746 ( 
.A(n_4604),
.Y(n_4746)
);

AO31x2_ASAP7_75t_L g4747 ( 
.A1(n_4677),
.A2(n_4428),
.A3(n_4441),
.B(n_4485),
.Y(n_4747)
);

BUFx2_ASAP7_75t_L g4748 ( 
.A(n_4586),
.Y(n_4748)
);

AND2x2_ASAP7_75t_L g4749 ( 
.A(n_4659),
.B(n_4485),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4616),
.B(n_4594),
.Y(n_4750)
);

CKINVDCx16_ASAP7_75t_R g4751 ( 
.A(n_4645),
.Y(n_4751)
);

AOI22xp33_ASAP7_75t_L g4752 ( 
.A1(n_4712),
.A2(n_4688),
.B1(n_4647),
.B2(n_4668),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4602),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4593),
.Y(n_4754)
);

OAI21xp33_ASAP7_75t_L g4755 ( 
.A1(n_4680),
.A2(n_4559),
.B(n_4451),
.Y(n_4755)
);

AND2x4_ASAP7_75t_SL g4756 ( 
.A(n_4669),
.B(n_4403),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4612),
.B(n_4646),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4591),
.Y(n_4758)
);

HB1xp67_ASAP7_75t_L g4759 ( 
.A(n_4652),
.Y(n_4759)
);

AND2x4_ASAP7_75t_L g4760 ( 
.A(n_4674),
.B(n_4477),
.Y(n_4760)
);

CKINVDCx16_ASAP7_75t_R g4761 ( 
.A(n_4645),
.Y(n_4761)
);

BUFx6f_ASAP7_75t_L g4762 ( 
.A(n_4626),
.Y(n_4762)
);

NAND3xp33_ASAP7_75t_L g4763 ( 
.A(n_4582),
.B(n_4435),
.C(n_4414),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4612),
.B(n_4494),
.Y(n_4764)
);

NOR2xp33_ASAP7_75t_R g4765 ( 
.A(n_4626),
.B(n_4403),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4657),
.Y(n_4766)
);

BUFx2_ASAP7_75t_SL g4767 ( 
.A(n_4719),
.Y(n_4767)
);

CKINVDCx5p33_ASAP7_75t_R g4768 ( 
.A(n_4673),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4583),
.B(n_4600),
.Y(n_4769)
);

OR2x2_ASAP7_75t_L g4770 ( 
.A(n_4654),
.B(n_4477),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4595),
.Y(n_4771)
);

BUFx3_ASAP7_75t_L g4772 ( 
.A(n_4698),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4631),
.B(n_4477),
.Y(n_4773)
);

INVxp67_ASAP7_75t_SL g4774 ( 
.A(n_4658),
.Y(n_4774)
);

AO31x2_ASAP7_75t_L g4775 ( 
.A1(n_4613),
.A2(n_4494),
.A3(n_4509),
.B(n_4524),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4629),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4628),
.Y(n_4777)
);

NOR2xp33_ASAP7_75t_L g4778 ( 
.A(n_4579),
.B(n_4557),
.Y(n_4778)
);

O2A1O1Ixp33_ASAP7_75t_L g4779 ( 
.A1(n_4702),
.A2(n_4512),
.B(n_4518),
.C(n_4421),
.Y(n_4779)
);

NAND2xp33_ASAP7_75t_SL g4780 ( 
.A(n_4707),
.B(n_4456),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4599),
.B(n_4552),
.Y(n_4781)
);

HB1xp67_ASAP7_75t_L g4782 ( 
.A(n_4588),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4605),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4590),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4606),
.Y(n_4785)
);

CKINVDCx16_ASAP7_75t_R g4786 ( 
.A(n_4709),
.Y(n_4786)
);

AOI22xp33_ASAP7_75t_L g4787 ( 
.A1(n_4688),
.A2(n_4508),
.B1(n_4545),
.B2(n_4548),
.Y(n_4787)
);

AOI22xp33_ASAP7_75t_L g4788 ( 
.A1(n_4668),
.A2(n_4508),
.B1(n_4545),
.B2(n_4548),
.Y(n_4788)
);

AND2x2_ASAP7_75t_L g4789 ( 
.A(n_4599),
.B(n_4524),
.Y(n_4789)
);

AOI22xp33_ASAP7_75t_L g4790 ( 
.A1(n_4693),
.A2(n_4523),
.B1(n_4516),
.B2(n_4413),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4696),
.B(n_4516),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4621),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4624),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4633),
.Y(n_4794)
);

BUFx3_ASAP7_75t_L g4795 ( 
.A(n_4700),
.Y(n_4795)
);

BUFx2_ASAP7_75t_L g4796 ( 
.A(n_4666),
.Y(n_4796)
);

AOI22xp33_ASAP7_75t_SL g4797 ( 
.A1(n_4670),
.A2(n_4523),
.B1(n_4509),
.B2(n_4564),
.Y(n_4797)
);

BUFx3_ASAP7_75t_L g4798 ( 
.A(n_4701),
.Y(n_4798)
);

AND2x2_ASAP7_75t_SL g4799 ( 
.A(n_4660),
.B(n_4509),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4610),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_4603),
.Y(n_4801)
);

OAI22xp5_ASAP7_75t_L g4802 ( 
.A1(n_4617),
.A2(n_240),
.B1(n_236),
.B2(n_238),
.Y(n_4802)
);

AOI21xp5_ASAP7_75t_L g4803 ( 
.A1(n_4639),
.A2(n_238),
.B(n_240),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4678),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_L g4805 ( 
.A1(n_4675),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4630),
.B(n_244),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_4665),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4667),
.Y(n_4808)
);

AO31x2_ASAP7_75t_L g4809 ( 
.A1(n_4695),
.A2(n_247),
.A3(n_245),
.B(n_246),
.Y(n_4809)
);

AND2x4_ASAP7_75t_L g4810 ( 
.A(n_4676),
.B(n_245),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4619),
.B(n_248),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4641),
.Y(n_4812)
);

INVx1_ASAP7_75t_L g4813 ( 
.A(n_4642),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4620),
.Y(n_4814)
);

NAND3xp33_ASAP7_75t_SL g4815 ( 
.A(n_4618),
.B(n_248),
.C(n_250),
.Y(n_4815)
);

AND2x2_ASAP7_75t_SL g4816 ( 
.A(n_4714),
.B(n_251),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4644),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_4673),
.Y(n_4818)
);

OAI22xp33_ASAP7_75t_L g4819 ( 
.A1(n_4675),
.A2(n_4597),
.B1(n_4638),
.B2(n_4710),
.Y(n_4819)
);

AND2x2_ASAP7_75t_L g4820 ( 
.A(n_4622),
.B(n_252),
.Y(n_4820)
);

INVx2_ASAP7_75t_L g4821 ( 
.A(n_4584),
.Y(n_4821)
);

NAND3xp33_ASAP7_75t_L g4822 ( 
.A(n_4720),
.B(n_253),
.C(n_255),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4682),
.Y(n_4823)
);

NAND3xp33_ASAP7_75t_SL g4824 ( 
.A(n_4635),
.B(n_253),
.C(n_256),
.Y(n_4824)
);

AND2x4_ASAP7_75t_L g4825 ( 
.A(n_4676),
.B(n_256),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4651),
.Y(n_4826)
);

NAND2xp33_ASAP7_75t_R g4827 ( 
.A(n_4705),
.B(n_258),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4681),
.B(n_259),
.Y(n_4828)
);

INVx2_ASAP7_75t_L g4829 ( 
.A(n_4604),
.Y(n_4829)
);

NOR3xp33_ASAP7_75t_SL g4830 ( 
.A(n_4686),
.B(n_259),
.C(n_261),
.Y(n_4830)
);

NAND2xp33_ASAP7_75t_R g4831 ( 
.A(n_4703),
.B(n_262),
.Y(n_4831)
);

OR2x2_ASAP7_75t_L g4832 ( 
.A(n_4607),
.B(n_262),
.Y(n_4832)
);

NAND2xp33_ASAP7_75t_SL g4833 ( 
.A(n_4694),
.B(n_263),
.Y(n_4833)
);

BUFx3_ASAP7_75t_L g4834 ( 
.A(n_4692),
.Y(n_4834)
);

BUFx2_ASAP7_75t_L g4835 ( 
.A(n_4666),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4691),
.Y(n_4836)
);

NOR2xp33_ASAP7_75t_R g4837 ( 
.A(n_4704),
.B(n_263),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4708),
.B(n_264),
.Y(n_4838)
);

CKINVDCx16_ASAP7_75t_R g4839 ( 
.A(n_4710),
.Y(n_4839)
);

BUFx4f_ASAP7_75t_SL g4840 ( 
.A(n_4713),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_4614),
.B(n_264),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_L g4842 ( 
.A(n_4687),
.B(n_265),
.Y(n_4842)
);

OAI22xp5_ASAP7_75t_L g4843 ( 
.A1(n_4717),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_R g4844 ( 
.A(n_4711),
.B(n_266),
.Y(n_4844)
);

NOR2xp33_ASAP7_75t_R g4845 ( 
.A(n_4689),
.B(n_267),
.Y(n_4845)
);

BUFx4f_ASAP7_75t_SL g4846 ( 
.A(n_4625),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4661),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4661),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4648),
.B(n_270),
.Y(n_4849)
);

AND2x4_ASAP7_75t_L g4850 ( 
.A(n_4637),
.B(n_271),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4637),
.B(n_272),
.Y(n_4851)
);

OR2x6_ASAP7_75t_L g4852 ( 
.A(n_4609),
.B(n_272),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4611),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4672),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4662),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4611),
.Y(n_4856)
);

BUFx2_ASAP7_75t_L g4857 ( 
.A(n_4662),
.Y(n_4857)
);

AND2x2_ASAP7_75t_L g4858 ( 
.A(n_4728),
.B(n_4653),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4819),
.A2(n_4690),
.B(n_4685),
.Y(n_4859)
);

AOI22xp33_ASAP7_75t_L g4860 ( 
.A1(n_4839),
.A2(n_4684),
.B1(n_4643),
.B2(n_4649),
.Y(n_4860)
);

OA21x2_ASAP7_75t_L g4861 ( 
.A1(n_4855),
.A2(n_4609),
.B(n_4684),
.Y(n_4861)
);

INVx2_ASAP7_75t_SL g4862 ( 
.A(n_4733),
.Y(n_4862)
);

BUFx3_ASAP7_75t_L g4863 ( 
.A(n_4733),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4836),
.Y(n_4864)
);

INVx1_ASAP7_75t_L g4865 ( 
.A(n_4722),
.Y(n_4865)
);

INVx5_ASAP7_75t_L g4866 ( 
.A(n_4762),
.Y(n_4866)
);

OAI322xp33_ASAP7_75t_L g4867 ( 
.A1(n_4802),
.A2(n_4718),
.A3(n_4643),
.B1(n_4715),
.B2(n_4716),
.C1(n_4706),
.C2(n_4587),
.Y(n_4867)
);

OR2x6_ASAP7_75t_L g4868 ( 
.A(n_4852),
.B(n_4649),
.Y(n_4868)
);

OR2x2_ASAP7_75t_L g4869 ( 
.A(n_4769),
.B(n_4653),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4722),
.Y(n_4870)
);

INVx3_ASAP7_75t_L g4871 ( 
.A(n_4721),
.Y(n_4871)
);

INVx2_ASAP7_75t_L g4872 ( 
.A(n_4836),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4836),
.Y(n_4873)
);

AND2x4_ASAP7_75t_L g4874 ( 
.A(n_4731),
.B(n_4671),
.Y(n_4874)
);

BUFx3_ASAP7_75t_L g4875 ( 
.A(n_4762),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4754),
.Y(n_4876)
);

OR2x2_ASAP7_75t_L g4877 ( 
.A(n_4784),
.B(n_4627),
.Y(n_4877)
);

AO21x2_ASAP7_75t_L g4878 ( 
.A1(n_4847),
.A2(n_4636),
.B(n_4679),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4776),
.B(n_4627),
.Y(n_4879)
);

OAI21xp5_ASAP7_75t_L g4880 ( 
.A1(n_4815),
.A2(n_273),
.B(n_274),
.Y(n_4880)
);

AO21x2_ASAP7_75t_L g4881 ( 
.A1(n_4847),
.A2(n_4848),
.B(n_4854),
.Y(n_4881)
);

BUFx6f_ASAP7_75t_L g4882 ( 
.A(n_4762),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4754),
.Y(n_4883)
);

AO21x2_ASAP7_75t_L g4884 ( 
.A1(n_4848),
.A2(n_274),
.B(n_275),
.Y(n_4884)
);

INVx1_ASAP7_75t_SL g4885 ( 
.A(n_4846),
.Y(n_4885)
);

INVx3_ASAP7_75t_L g4886 ( 
.A(n_4728),
.Y(n_4886)
);

OR2x6_ASAP7_75t_L g4887 ( 
.A(n_4852),
.B(n_275),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4771),
.Y(n_4888)
);

INVx2_ASAP7_75t_L g4889 ( 
.A(n_4796),
.Y(n_4889)
);

BUFx2_ASAP7_75t_L g4890 ( 
.A(n_4731),
.Y(n_4890)
);

INVx4_ASAP7_75t_L g4891 ( 
.A(n_4745),
.Y(n_4891)
);

OAI211xp5_ASAP7_75t_L g4892 ( 
.A1(n_4824),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_4892)
);

INVx2_ASAP7_75t_L g4893 ( 
.A(n_4835),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4771),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4799),
.B(n_276),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4759),
.Y(n_4896)
);

OAI221xp5_ASAP7_75t_SL g4897 ( 
.A1(n_4805),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.C(n_281),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4736),
.Y(n_4898)
);

AO21x2_ASAP7_75t_L g4899 ( 
.A1(n_4853),
.A2(n_279),
.B(n_284),
.Y(n_4899)
);

HB1xp67_ASAP7_75t_L g4900 ( 
.A(n_4857),
.Y(n_4900)
);

OR2x2_ASAP7_75t_L g4901 ( 
.A(n_4723),
.B(n_284),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4756),
.B(n_285),
.Y(n_4902)
);

OR2x6_ASAP7_75t_L g4903 ( 
.A(n_4767),
.B(n_286),
.Y(n_4903)
);

OR2x2_ASAP7_75t_L g4904 ( 
.A(n_4823),
.B(n_287),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4829),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4826),
.B(n_287),
.Y(n_4906)
);

AOI21xp5_ASAP7_75t_SL g4907 ( 
.A1(n_4822),
.A2(n_289),
.B(n_290),
.Y(n_4907)
);

INVxp67_ASAP7_75t_L g4908 ( 
.A(n_4827),
.Y(n_4908)
);

INVxp67_ASAP7_75t_L g4909 ( 
.A(n_4831),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4781),
.B(n_291),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4749),
.B(n_292),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4739),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4757),
.B(n_4789),
.Y(n_4913)
);

INVx2_ASAP7_75t_SL g4914 ( 
.A(n_4725),
.Y(n_4914)
);

AOI22xp33_ASAP7_75t_L g4915 ( 
.A1(n_4752),
.A2(n_299),
.B1(n_296),
.B2(n_297),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4734),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4737),
.Y(n_4917)
);

HB1xp67_ASAP7_75t_L g4918 ( 
.A(n_4776),
.Y(n_4918)
);

NOR2xp33_ASAP7_75t_L g4919 ( 
.A(n_4745),
.B(n_296),
.Y(n_4919)
);

INVx2_ASAP7_75t_L g4920 ( 
.A(n_4834),
.Y(n_4920)
);

AO21x2_ASAP7_75t_L g4921 ( 
.A1(n_4853),
.A2(n_299),
.B(n_300),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4777),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4764),
.B(n_301),
.Y(n_4923)
);

BUFx3_ASAP7_75t_L g4924 ( 
.A(n_4727),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4804),
.Y(n_4925)
);

BUFx2_ASAP7_75t_L g4926 ( 
.A(n_4765),
.Y(n_4926)
);

AND2x4_ASAP7_75t_SL g4927 ( 
.A(n_4732),
.B(n_4724),
.Y(n_4927)
);

NAND3xp33_ASAP7_75t_L g4928 ( 
.A(n_4849),
.B(n_302),
.C(n_303),
.Y(n_4928)
);

AO21x2_ASAP7_75t_L g4929 ( 
.A1(n_4856),
.A2(n_304),
.B(n_305),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4808),
.Y(n_4930)
);

HB1xp67_ASAP7_75t_L g4931 ( 
.A(n_4748),
.Y(n_4931)
);

OR2x2_ASAP7_75t_L g4932 ( 
.A(n_4826),
.B(n_305),
.Y(n_4932)
);

OR2x6_ASAP7_75t_L g4933 ( 
.A(n_4850),
.B(n_306),
.Y(n_4933)
);

OR2x2_ASAP7_75t_L g4934 ( 
.A(n_4794),
.B(n_4774),
.Y(n_4934)
);

INVxp67_ASAP7_75t_SL g4935 ( 
.A(n_4851),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4742),
.B(n_307),
.Y(n_4936)
);

OAI22xp33_ASAP7_75t_L g4937 ( 
.A1(n_4751),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4758),
.B(n_308),
.Y(n_4938)
);

OR2x2_ASAP7_75t_L g4939 ( 
.A(n_4782),
.B(n_311),
.Y(n_4939)
);

OR2x2_ASAP7_75t_L g4940 ( 
.A(n_4800),
.B(n_311),
.Y(n_4940)
);

OA21x2_ASAP7_75t_L g4941 ( 
.A1(n_4785),
.A2(n_312),
.B(n_313),
.Y(n_4941)
);

AND2x2_ASAP7_75t_L g4942 ( 
.A(n_4791),
.B(n_312),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4801),
.B(n_313),
.Y(n_4943)
);

AOI22xp5_ASAP7_75t_L g4944 ( 
.A1(n_4763),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_4778),
.B(n_314),
.Y(n_4945)
);

BUFx3_ASAP7_75t_L g4946 ( 
.A(n_4766),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4735),
.Y(n_4947)
);

HB1xp67_ASAP7_75t_L g4948 ( 
.A(n_4785),
.Y(n_4948)
);

BUFx3_ASAP7_75t_L g4949 ( 
.A(n_4768),
.Y(n_4949)
);

OR2x2_ASAP7_75t_L g4950 ( 
.A(n_4814),
.B(n_315),
.Y(n_4950)
);

INVx2_ASAP7_75t_L g4951 ( 
.A(n_4746),
.Y(n_4951)
);

AOI221xp5_ASAP7_75t_L g4952 ( 
.A1(n_4738),
.A2(n_4755),
.B1(n_4843),
.B2(n_4841),
.C(n_4803),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4760),
.B(n_316),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_SL g4954 ( 
.A1(n_4850),
.A2(n_4779),
.B(n_4810),
.Y(n_4954)
);

INVx2_ASAP7_75t_L g4955 ( 
.A(n_4746),
.Y(n_4955)
);

AO21x2_ASAP7_75t_L g4956 ( 
.A1(n_4845),
.A2(n_318),
.B(n_319),
.Y(n_4956)
);

AOI221xp5_ASAP7_75t_L g4957 ( 
.A1(n_4741),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.C(n_322),
.Y(n_4957)
);

AO21x2_ASAP7_75t_L g4958 ( 
.A1(n_4837),
.A2(n_322),
.B(n_325),
.Y(n_4958)
);

AO21x2_ASAP7_75t_L g4959 ( 
.A1(n_4844),
.A2(n_326),
.B(n_327),
.Y(n_4959)
);

BUFx3_ASAP7_75t_L g4960 ( 
.A(n_4818),
.Y(n_4960)
);

INVx2_ASAP7_75t_SL g4961 ( 
.A(n_4840),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4821),
.Y(n_4962)
);

INVx4_ASAP7_75t_SL g4963 ( 
.A(n_4809),
.Y(n_4963)
);

HB1xp67_ASAP7_75t_L g4964 ( 
.A(n_4817),
.Y(n_4964)
);

BUFx6f_ASAP7_75t_L g4965 ( 
.A(n_4891),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4865),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4890),
.B(n_4797),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4935),
.B(n_4816),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4935),
.B(n_4952),
.Y(n_4969)
);

OAI22xp5_ASAP7_75t_L g4970 ( 
.A1(n_4860),
.A2(n_4761),
.B1(n_4788),
.B2(n_4790),
.Y(n_4970)
);

AND2x2_ASAP7_75t_L g4971 ( 
.A(n_4886),
.B(n_4760),
.Y(n_4971)
);

INVx1_ASAP7_75t_L g4972 ( 
.A(n_4870),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4963),
.Y(n_4973)
);

INVx2_ASAP7_75t_L g4974 ( 
.A(n_4963),
.Y(n_4974)
);

INVxp67_ASAP7_75t_L g4975 ( 
.A(n_4908),
.Y(n_4975)
);

AND2x2_ASAP7_75t_L g4976 ( 
.A(n_4886),
.B(n_4750),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4963),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4952),
.B(n_4811),
.Y(n_4978)
);

AOI22xp33_ASAP7_75t_L g4979 ( 
.A1(n_4859),
.A2(n_4744),
.B1(n_4833),
.B2(n_4740),
.Y(n_4979)
);

INVxp67_ASAP7_75t_L g4980 ( 
.A(n_4908),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4876),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4864),
.B(n_4820),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4913),
.B(n_4795),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4874),
.B(n_4786),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4874),
.B(n_4753),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4883),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4888),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4894),
.Y(n_4988)
);

BUFx2_ASAP7_75t_L g4989 ( 
.A(n_4903),
.Y(n_4989)
);

BUFx3_ASAP7_75t_L g4990 ( 
.A(n_4866),
.Y(n_4990)
);

AND2x4_ASAP7_75t_L g4991 ( 
.A(n_4871),
.B(n_4775),
.Y(n_4991)
);

INVx3_ASAP7_75t_L g4992 ( 
.A(n_4891),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4948),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4948),
.Y(n_4994)
);

INVx2_ASAP7_75t_SL g4995 ( 
.A(n_4866),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4964),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4964),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4872),
.B(n_4810),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4881),
.Y(n_4999)
);

INVxp67_ASAP7_75t_SL g5000 ( 
.A(n_4909),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4916),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_4881),
.Y(n_5002)
);

AND2x4_ASAP7_75t_L g5003 ( 
.A(n_4871),
.B(n_4775),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4873),
.B(n_4828),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4898),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4912),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4914),
.B(n_4825),
.Y(n_5007)
);

BUFx4f_ASAP7_75t_SL g5008 ( 
.A(n_4882),
.Y(n_5008)
);

AOI22xp33_ASAP7_75t_L g5009 ( 
.A1(n_4859),
.A2(n_4957),
.B1(n_4909),
.B2(n_4928),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4878),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4917),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4922),
.Y(n_5012)
);

NAND3xp33_ASAP7_75t_L g5013 ( 
.A(n_4944),
.B(n_4957),
.C(n_4928),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4925),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4889),
.B(n_4825),
.Y(n_5015)
);

AOI22xp5_ASAP7_75t_L g5016 ( 
.A1(n_4944),
.A2(n_4780),
.B1(n_4830),
.B2(n_4787),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4893),
.B(n_4772),
.Y(n_5017)
);

INVx2_ASAP7_75t_SL g5018 ( 
.A(n_4866),
.Y(n_5018)
);

BUFx3_ASAP7_75t_L g5019 ( 
.A(n_4863),
.Y(n_5019)
);

INVx2_ASAP7_75t_L g5020 ( 
.A(n_4878),
.Y(n_5020)
);

OR2x2_ASAP7_75t_L g5021 ( 
.A(n_4934),
.B(n_4747),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_4931),
.B(n_4747),
.Y(n_5022)
);

AOI22xp33_ASAP7_75t_SL g5023 ( 
.A1(n_4956),
.A2(n_4798),
.B1(n_4806),
.B2(n_4832),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_4903),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4920),
.B(n_4770),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_4930),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4918),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4918),
.Y(n_5028)
);

INVx2_ASAP7_75t_L g5029 ( 
.A(n_4903),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4901),
.B(n_4838),
.Y(n_5030)
);

AND2x2_ASAP7_75t_L g5031 ( 
.A(n_4926),
.B(n_4885),
.Y(n_5031)
);

INVxp67_ASAP7_75t_L g5032 ( 
.A(n_4958),
.Y(n_5032)
);

NAND2x1_ASAP7_75t_L g5033 ( 
.A(n_4868),
.B(n_4792),
.Y(n_5033)
);

AOI22xp33_ASAP7_75t_SL g5034 ( 
.A1(n_4956),
.A2(n_4842),
.B1(n_4726),
.B2(n_4747),
.Y(n_5034)
);

AND2x4_ASAP7_75t_L g5035 ( 
.A(n_4951),
.B(n_4775),
.Y(n_5035)
);

OR2x6_ASAP7_75t_L g5036 ( 
.A(n_5018),
.B(n_4907),
.Y(n_5036)
);

AND4x1_ASAP7_75t_L g5037 ( 
.A(n_5009),
.B(n_4954),
.C(n_4880),
.D(n_4895),
.Y(n_5037)
);

HB1xp67_ASAP7_75t_L g5038 ( 
.A(n_4989),
.Y(n_5038)
);

AOI22xp33_ASAP7_75t_L g5039 ( 
.A1(n_4979),
.A2(n_4861),
.B1(n_4868),
.B2(n_4885),
.Y(n_5039)
);

AOI33xp33_ASAP7_75t_L g5040 ( 
.A1(n_5009),
.A2(n_4937),
.A3(n_4915),
.B1(n_4896),
.B2(n_4927),
.B3(n_4862),
.Y(n_5040)
);

AOI22xp33_ASAP7_75t_L g5041 ( 
.A1(n_4979),
.A2(n_4861),
.B1(n_4868),
.B2(n_4880),
.Y(n_5041)
);

AOI22xp33_ASAP7_75t_L g5042 ( 
.A1(n_5013),
.A2(n_4875),
.B1(n_4882),
.B2(n_4958),
.Y(n_5042)
);

INVxp67_ASAP7_75t_L g5043 ( 
.A(n_5000),
.Y(n_5043)
);

BUFx2_ASAP7_75t_L g5044 ( 
.A(n_5000),
.Y(n_5044)
);

HB1xp67_ASAP7_75t_L g5045 ( 
.A(n_4975),
.Y(n_5045)
);

AOI22xp33_ASAP7_75t_L g5046 ( 
.A1(n_4969),
.A2(n_4882),
.B1(n_4959),
.B2(n_4867),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4993),
.Y(n_5047)
);

NOR2x1_ASAP7_75t_L g5048 ( 
.A(n_4990),
.B(n_4959),
.Y(n_5048)
);

OAI221xp5_ASAP7_75t_L g5049 ( 
.A1(n_5034),
.A2(n_4892),
.B1(n_4887),
.B2(n_4897),
.C(n_4945),
.Y(n_5049)
);

AOI221xp5_ASAP7_75t_L g5050 ( 
.A1(n_5032),
.A2(n_4867),
.B1(n_4892),
.B2(n_4897),
.C(n_4900),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4984),
.B(n_4955),
.Y(n_5051)
);

OAI31xp33_ASAP7_75t_L g5052 ( 
.A1(n_4970),
.A2(n_4900),
.A3(n_4919),
.B(n_4939),
.Y(n_5052)
);

INVx2_ASAP7_75t_L g5053 ( 
.A(n_4990),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_5033),
.A2(n_4879),
.B(n_4858),
.Y(n_5054)
);

OR2x2_ASAP7_75t_L g5055 ( 
.A(n_5032),
.B(n_4947),
.Y(n_5055)
);

AOI33xp33_ASAP7_75t_L g5056 ( 
.A1(n_5034),
.A2(n_4943),
.A3(n_4923),
.B1(n_4953),
.B2(n_4961),
.B3(n_4936),
.Y(n_5056)
);

OR2x2_ASAP7_75t_L g5057 ( 
.A(n_4968),
.B(n_4905),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_5031),
.B(n_4962),
.Y(n_5058)
);

AND2x2_ASAP7_75t_L g5059 ( 
.A(n_4971),
.B(n_4869),
.Y(n_5059)
);

CKINVDCx5p33_ASAP7_75t_R g5060 ( 
.A(n_4965),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_5018),
.Y(n_5061)
);

OAI221xp5_ASAP7_75t_L g5062 ( 
.A1(n_4975),
.A2(n_4887),
.B1(n_4933),
.B2(n_4949),
.C(n_4960),
.Y(n_5062)
);

HB1xp67_ASAP7_75t_L g5063 ( 
.A(n_4980),
.Y(n_5063)
);

OAI31xp33_ASAP7_75t_L g5064 ( 
.A1(n_4980),
.A2(n_4902),
.A3(n_4932),
.B(n_4906),
.Y(n_5064)
);

AOI22xp33_ASAP7_75t_L g5065 ( 
.A1(n_4967),
.A2(n_4992),
.B1(n_4965),
.B2(n_4978),
.Y(n_5065)
);

OAI22xp5_ASAP7_75t_L g5066 ( 
.A1(n_5023),
.A2(n_4887),
.B1(n_4933),
.B2(n_4941),
.Y(n_5066)
);

AND2x2_ASAP7_75t_L g5067 ( 
.A(n_4976),
.B(n_4946),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_5023),
.B(n_4904),
.Y(n_5068)
);

AOI22xp33_ASAP7_75t_L g5069 ( 
.A1(n_4992),
.A2(n_4884),
.B1(n_4921),
.B2(n_4899),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_4994),
.Y(n_5070)
);

OR2x2_ASAP7_75t_L g5071 ( 
.A(n_5027),
.B(n_4879),
.Y(n_5071)
);

INVx2_ASAP7_75t_L g5072 ( 
.A(n_4999),
.Y(n_5072)
);

OAI221xp5_ASAP7_75t_L g5073 ( 
.A1(n_5016),
.A2(n_4933),
.B1(n_4938),
.B2(n_4924),
.C(n_4940),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_L g5074 ( 
.A(n_5024),
.B(n_4911),
.Y(n_5074)
);

INVx2_ASAP7_75t_L g5075 ( 
.A(n_4999),
.Y(n_5075)
);

AOI222xp33_ASAP7_75t_L g5076 ( 
.A1(n_5024),
.A2(n_4942),
.B1(n_4910),
.B2(n_4730),
.C1(n_4884),
.C2(n_4921),
.Y(n_5076)
);

OA21x2_ASAP7_75t_L g5077 ( 
.A1(n_5010),
.A2(n_4877),
.B(n_4950),
.Y(n_5077)
);

NAND3xp33_ASAP7_75t_L g5078 ( 
.A(n_5010),
.B(n_4941),
.C(n_4813),
.Y(n_5078)
);

BUFx12f_ASAP7_75t_L g5079 ( 
.A(n_4965),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_4965),
.A2(n_4899),
.B1(n_4929),
.B2(n_4807),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_4985),
.B(n_4793),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_5067),
.B(n_5038),
.Y(n_5082)
);

AND2x4_ASAP7_75t_L g5083 ( 
.A(n_5044),
.B(n_5020),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5045),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_5067),
.B(n_4995),
.Y(n_5085)
);

AND2x2_ASAP7_75t_L g5086 ( 
.A(n_5051),
.B(n_5058),
.Y(n_5086)
);

HB1xp67_ASAP7_75t_L g5087 ( 
.A(n_5063),
.Y(n_5087)
);

HB1xp67_ASAP7_75t_L g5088 ( 
.A(n_5043),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_5055),
.Y(n_5089)
);

INVxp67_ASAP7_75t_SL g5090 ( 
.A(n_5048),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_5055),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_5036),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_5051),
.B(n_5029),
.Y(n_5093)
);

INVx2_ASAP7_75t_L g5094 ( 
.A(n_5036),
.Y(n_5094)
);

OR2x2_ASAP7_75t_L g5095 ( 
.A(n_5068),
.B(n_5028),
.Y(n_5095)
);

AND2x2_ASAP7_75t_L g5096 ( 
.A(n_5058),
.B(n_5029),
.Y(n_5096)
);

AND2x2_ASAP7_75t_L g5097 ( 
.A(n_5053),
.B(n_5019),
.Y(n_5097)
);

AND2x2_ASAP7_75t_L g5098 ( 
.A(n_5053),
.B(n_5019),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_5072),
.Y(n_5099)
);

INVx2_ASAP7_75t_L g5100 ( 
.A(n_5036),
.Y(n_5100)
);

AND2x2_ASAP7_75t_SL g5101 ( 
.A(n_5037),
.B(n_5020),
.Y(n_5101)
);

INVx2_ASAP7_75t_L g5102 ( 
.A(n_5036),
.Y(n_5102)
);

AND2x2_ASAP7_75t_L g5103 ( 
.A(n_5059),
.B(n_5017),
.Y(n_5103)
);

HB1xp67_ASAP7_75t_L g5104 ( 
.A(n_5077),
.Y(n_5104)
);

AND2x2_ASAP7_75t_L g5105 ( 
.A(n_5059),
.B(n_4983),
.Y(n_5105)
);

AND2x2_ASAP7_75t_L g5106 ( 
.A(n_5061),
.B(n_5025),
.Y(n_5106)
);

AND2x2_ASAP7_75t_L g5107 ( 
.A(n_5061),
.B(n_5015),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5072),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_5077),
.Y(n_5109)
);

AND2x2_ASAP7_75t_L g5110 ( 
.A(n_5081),
.B(n_5065),
.Y(n_5110)
);

INVx1_ASAP7_75t_SL g5111 ( 
.A(n_5060),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_5050),
.B(n_5001),
.Y(n_5112)
);

AND2x4_ASAP7_75t_SL g5113 ( 
.A(n_5046),
.B(n_5007),
.Y(n_5113)
);

AND2x2_ASAP7_75t_L g5114 ( 
.A(n_5081),
.B(n_4973),
.Y(n_5114)
);

INVx2_ASAP7_75t_L g5115 ( 
.A(n_5077),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_5060),
.B(n_4973),
.Y(n_5116)
);

OR2x2_ASAP7_75t_L g5117 ( 
.A(n_5104),
.B(n_5066),
.Y(n_5117)
);

BUFx3_ASAP7_75t_L g5118 ( 
.A(n_5097),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_5087),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_5111),
.B(n_5062),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_5082),
.B(n_5079),
.Y(n_5121)
);

AND2x2_ASAP7_75t_L g5122 ( 
.A(n_5082),
.B(n_5079),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_5104),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_5109),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_5085),
.B(n_5056),
.Y(n_5125)
);

AND2x2_ASAP7_75t_L g5126 ( 
.A(n_5085),
.B(n_5056),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5083),
.Y(n_5127)
);

AND2x2_ASAP7_75t_L g5128 ( 
.A(n_5097),
.B(n_5042),
.Y(n_5128)
);

AND2x2_ASAP7_75t_L g5129 ( 
.A(n_5098),
.B(n_4974),
.Y(n_5129)
);

NOR2xp33_ASAP7_75t_L g5130 ( 
.A(n_5111),
.B(n_5073),
.Y(n_5130)
);

INVxp67_ASAP7_75t_SL g5131 ( 
.A(n_5090),
.Y(n_5131)
);

INVxp67_ASAP7_75t_L g5132 ( 
.A(n_5098),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_5086),
.B(n_4974),
.Y(n_5133)
);

INVxp67_ASAP7_75t_L g5134 ( 
.A(n_5093),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5083),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_5086),
.B(n_4977),
.Y(n_5136)
);

AND2x4_ASAP7_75t_L g5137 ( 
.A(n_5090),
.B(n_4977),
.Y(n_5137)
);

NAND2xp5_ASAP7_75t_L g5138 ( 
.A(n_5093),
.B(n_5052),
.Y(n_5138)
);

OR2x2_ASAP7_75t_L g5139 ( 
.A(n_5095),
.B(n_5074),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_5105),
.B(n_5076),
.Y(n_5140)
);

INVx2_ASAP7_75t_L g5141 ( 
.A(n_5118),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_5118),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5127),
.Y(n_5143)
);

OR2x2_ASAP7_75t_L g5144 ( 
.A(n_5139),
.B(n_5095),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5135),
.Y(n_5145)
);

OR2x2_ASAP7_75t_L g5146 ( 
.A(n_5132),
.B(n_5084),
.Y(n_5146)
);

NAND2xp5_ASAP7_75t_L g5147 ( 
.A(n_5131),
.B(n_5084),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_5125),
.B(n_5096),
.Y(n_5148)
);

INVx1_ASAP7_75t_L g5149 ( 
.A(n_5123),
.Y(n_5149)
);

OR2x2_ASAP7_75t_L g5150 ( 
.A(n_5134),
.B(n_5088),
.Y(n_5150)
);

CKINVDCx16_ASAP7_75t_R g5151 ( 
.A(n_5121),
.Y(n_5151)
);

INVx2_ASAP7_75t_SL g5152 ( 
.A(n_5121),
.Y(n_5152)
);

AND2x2_ASAP7_75t_L g5153 ( 
.A(n_5122),
.B(n_5105),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5124),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_5133),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_5140),
.B(n_5112),
.Y(n_5156)
);

NAND2x1_ASAP7_75t_L g5157 ( 
.A(n_5122),
.B(n_5083),
.Y(n_5157)
);

INVxp67_ASAP7_75t_SL g5158 ( 
.A(n_5117),
.Y(n_5158)
);

NAND2x1_ASAP7_75t_L g5159 ( 
.A(n_5137),
.B(n_5083),
.Y(n_5159)
);

INVxp67_ASAP7_75t_SL g5160 ( 
.A(n_5117),
.Y(n_5160)
);

OAI21xp5_ASAP7_75t_L g5161 ( 
.A1(n_5138),
.A2(n_5101),
.B(n_5049),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_5140),
.B(n_5125),
.Y(n_5162)
);

AND2x2_ASAP7_75t_L g5163 ( 
.A(n_5128),
.B(n_5103),
.Y(n_5163)
);

OR2x2_ASAP7_75t_L g5164 ( 
.A(n_5119),
.B(n_5096),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5159),
.Y(n_5165)
);

INVx2_ASAP7_75t_L g5166 ( 
.A(n_5157),
.Y(n_5166)
);

INVx4_ASAP7_75t_L g5167 ( 
.A(n_5141),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_5155),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_5164),
.Y(n_5169)
);

INVx1_ASAP7_75t_SL g5170 ( 
.A(n_5163),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5158),
.B(n_5126),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_5160),
.B(n_5126),
.Y(n_5172)
);

AOI32xp33_ASAP7_75t_L g5173 ( 
.A1(n_5156),
.A2(n_5039),
.A3(n_5041),
.B1(n_5113),
.B2(n_5112),
.Y(n_5173)
);

HB1xp67_ASAP7_75t_L g5174 ( 
.A(n_5151),
.Y(n_5174)
);

NOR2xp67_ASAP7_75t_L g5175 ( 
.A(n_5152),
.B(n_5115),
.Y(n_5175)
);

INVx2_ASAP7_75t_SL g5176 ( 
.A(n_5153),
.Y(n_5176)
);

BUFx2_ASAP7_75t_L g5177 ( 
.A(n_5142),
.Y(n_5177)
);

OAI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_5156),
.A2(n_5069),
.B1(n_5080),
.B2(n_5101),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_5146),
.Y(n_5179)
);

INVxp67_ASAP7_75t_SL g5180 ( 
.A(n_5144),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_5148),
.B(n_5110),
.Y(n_5181)
);

HB1xp67_ASAP7_75t_L g5182 ( 
.A(n_5175),
.Y(n_5182)
);

INVx1_ASAP7_75t_SL g5183 ( 
.A(n_5170),
.Y(n_5183)
);

OR2x2_ASAP7_75t_L g5184 ( 
.A(n_5170),
.B(n_5162),
.Y(n_5184)
);

INVxp33_ASAP7_75t_L g5185 ( 
.A(n_5174),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5175),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5180),
.Y(n_5187)
);

INVx1_ASAP7_75t_SL g5188 ( 
.A(n_5177),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_5176),
.B(n_5129),
.Y(n_5189)
);

NOR2x1_ASAP7_75t_L g5190 ( 
.A(n_5166),
.B(n_5147),
.Y(n_5190)
);

INVx4_ASAP7_75t_L g5191 ( 
.A(n_5167),
.Y(n_5191)
);

BUFx2_ASAP7_75t_L g5192 ( 
.A(n_5165),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_5167),
.Y(n_5193)
);

OR2x2_ASAP7_75t_L g5194 ( 
.A(n_5184),
.B(n_5171),
.Y(n_5194)
);

NOR2xp33_ASAP7_75t_L g5195 ( 
.A(n_5185),
.B(n_5130),
.Y(n_5195)
);

AOI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_5189),
.A2(n_5161),
.B(n_5178),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5182),
.Y(n_5197)
);

AOI22xp5_ASAP7_75t_L g5198 ( 
.A1(n_5188),
.A2(n_5162),
.B1(n_5161),
.B2(n_5120),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_5186),
.Y(n_5199)
);

OAI31xp33_ASAP7_75t_L g5200 ( 
.A1(n_5183),
.A2(n_5113),
.A3(n_5172),
.B(n_5128),
.Y(n_5200)
);

AOI21xp33_ASAP7_75t_L g5201 ( 
.A1(n_5187),
.A2(n_5101),
.B(n_5147),
.Y(n_5201)
);

AND2x4_ASAP7_75t_L g5202 ( 
.A(n_5191),
.B(n_5143),
.Y(n_5202)
);

INVxp67_ASAP7_75t_L g5203 ( 
.A(n_5190),
.Y(n_5203)
);

NOR2xp33_ASAP7_75t_L g5204 ( 
.A(n_5191),
.B(n_5150),
.Y(n_5204)
);

OAI321xp33_ASAP7_75t_L g5205 ( 
.A1(n_5192),
.A2(n_5173),
.A3(n_5169),
.B1(n_5181),
.B2(n_5145),
.C(n_5179),
.Y(n_5205)
);

OAI322xp33_ASAP7_75t_L g5206 ( 
.A1(n_5193),
.A2(n_5154),
.A3(n_5149),
.B1(n_5091),
.B2(n_5089),
.C1(n_5168),
.C2(n_5092),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_L g5207 ( 
.A(n_5183),
.B(n_5129),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5207),
.Y(n_5208)
);

NAND3x2_ASAP7_75t_L g5209 ( 
.A(n_5194),
.B(n_5116),
.C(n_5137),
.Y(n_5209)
);

NAND2xp5_ASAP7_75t_L g5210 ( 
.A(n_5198),
.B(n_5116),
.Y(n_5210)
);

AOI322xp5_ASAP7_75t_L g5211 ( 
.A1(n_5195),
.A2(n_5110),
.A3(n_5107),
.B1(n_5091),
.B2(n_5089),
.C1(n_5106),
.C2(n_5133),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5202),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5202),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_5197),
.B(n_5107),
.Y(n_5214)
);

AOI21xp5_ASAP7_75t_L g5215 ( 
.A1(n_5203),
.A2(n_5115),
.B(n_5094),
.Y(n_5215)
);

NAND2x1p5_ASAP7_75t_L g5216 ( 
.A(n_5204),
.B(n_5092),
.Y(n_5216)
);

AOI211xp5_ASAP7_75t_L g5217 ( 
.A1(n_5201),
.A2(n_5094),
.B(n_5100),
.C(n_5092),
.Y(n_5217)
);

OR2x2_ASAP7_75t_L g5218 ( 
.A(n_5209),
.B(n_5200),
.Y(n_5218)
);

NOR2xp33_ASAP7_75t_L g5219 ( 
.A(n_5210),
.B(n_5206),
.Y(n_5219)
);

OR2x2_ASAP7_75t_L g5220 ( 
.A(n_5216),
.B(n_5094),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_L g5221 ( 
.A(n_5211),
.B(n_5196),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_5214),
.B(n_5136),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_5212),
.Y(n_5223)
);

NOR2xp33_ASAP7_75t_SL g5224 ( 
.A(n_5213),
.B(n_5008),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_5217),
.B(n_5199),
.Y(n_5225)
);

AND2x2_ASAP7_75t_L g5226 ( 
.A(n_5208),
.B(n_5136),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_5215),
.A2(n_5113),
.B1(n_5100),
.B2(n_5102),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_SL g5228 ( 
.A(n_5227),
.B(n_5100),
.Y(n_5228)
);

NOR4xp25_ASAP7_75t_L g5229 ( 
.A(n_5221),
.B(n_5205),
.C(n_5102),
.D(n_5115),
.Y(n_5229)
);

AND4x1_ASAP7_75t_L g5230 ( 
.A(n_5224),
.B(n_5040),
.C(n_5106),
.D(n_5064),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5222),
.Y(n_5231)
);

NAND3xp33_ASAP7_75t_L g5232 ( 
.A(n_5219),
.B(n_5102),
.C(n_5137),
.Y(n_5232)
);

NAND4xp25_ASAP7_75t_L g5233 ( 
.A(n_5218),
.B(n_5225),
.C(n_5226),
.D(n_5223),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_5220),
.B(n_5103),
.Y(n_5234)
);

AOI22xp5_ASAP7_75t_L g5235 ( 
.A1(n_5224),
.A2(n_5114),
.B1(n_5099),
.B2(n_5108),
.Y(n_5235)
);

AOI221xp5_ASAP7_75t_L g5236 ( 
.A1(n_5219),
.A2(n_5108),
.B1(n_5099),
.B2(n_5070),
.C(n_5047),
.Y(n_5236)
);

NOR2xp33_ASAP7_75t_L g5237 ( 
.A(n_5224),
.B(n_5008),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_5222),
.B(n_5040),
.Y(n_5238)
);

NAND2x1_ASAP7_75t_L g5239 ( 
.A(n_5222),
.B(n_5114),
.Y(n_5239)
);

NAND3xp33_ASAP7_75t_L g5240 ( 
.A(n_5224),
.B(n_5075),
.C(n_5071),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_5220),
.Y(n_5241)
);

INVx1_ASAP7_75t_SL g5242 ( 
.A(n_5222),
.Y(n_5242)
);

AOI22xp5_ASAP7_75t_L g5243 ( 
.A1(n_5224),
.A2(n_5075),
.B1(n_5057),
.B2(n_4996),
.Y(n_5243)
);

NOR2xp33_ASAP7_75t_L g5244 ( 
.A(n_5224),
.B(n_5071),
.Y(n_5244)
);

CKINVDCx5p33_ASAP7_75t_R g5245 ( 
.A(n_5219),
.Y(n_5245)
);

OAI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_5232),
.A2(n_5054),
.B(n_5002),
.Y(n_5246)
);

AOI21xp33_ASAP7_75t_SL g5247 ( 
.A1(n_5229),
.A2(n_5054),
.B(n_5078),
.Y(n_5247)
);

OR2x2_ASAP7_75t_L g5248 ( 
.A(n_5239),
.B(n_5021),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_5240),
.A2(n_5002),
.B(n_5022),
.Y(n_5249)
);

AND4x1_ASAP7_75t_L g5250 ( 
.A(n_5237),
.B(n_4997),
.C(n_5030),
.D(n_5006),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_SL g5251 ( 
.A(n_5235),
.B(n_4991),
.Y(n_5251)
);

NAND5xp2_ASAP7_75t_L g5252 ( 
.A(n_5236),
.B(n_4998),
.C(n_5014),
.D(n_5012),
.E(n_5011),
.Y(n_5252)
);

AOI221xp5_ASAP7_75t_L g5253 ( 
.A1(n_5228),
.A2(n_5026),
.B1(n_5005),
.B2(n_4991),
.C(n_5003),
.Y(n_5253)
);

NOR2x1_ASAP7_75t_L g5254 ( 
.A(n_5233),
.B(n_4991),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_5230),
.B(n_4966),
.Y(n_5255)
);

AND4x1_ASAP7_75t_L g5256 ( 
.A(n_5231),
.B(n_4972),
.C(n_4986),
.D(n_4981),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5242),
.B(n_5003),
.Y(n_5257)
);

HB1xp67_ASAP7_75t_L g5258 ( 
.A(n_5241),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_5244),
.A2(n_5003),
.B1(n_5035),
.B2(n_4987),
.Y(n_5259)
);

NOR2x1_ASAP7_75t_L g5260 ( 
.A(n_5234),
.B(n_4988),
.Y(n_5260)
);

O2A1O1Ixp33_ASAP7_75t_L g5261 ( 
.A1(n_5238),
.A2(n_5035),
.B(n_4929),
.C(n_5004),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5243),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_L g5263 ( 
.A(n_5245),
.B(n_4982),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5234),
.Y(n_5264)
);

AND2x2_ASAP7_75t_L g5265 ( 
.A(n_5242),
.B(n_5035),
.Y(n_5265)
);

NOR4xp25_ASAP7_75t_L g5266 ( 
.A(n_5232),
.B(n_4729),
.C(n_330),
.D(n_328),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5234),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5234),
.Y(n_5268)
);

NOR2x1_ASAP7_75t_L g5269 ( 
.A(n_5232),
.B(n_4743),
.Y(n_5269)
);

BUFx3_ASAP7_75t_L g5270 ( 
.A(n_5239),
.Y(n_5270)
);

NOR2xp33_ASAP7_75t_L g5271 ( 
.A(n_5258),
.B(n_329),
.Y(n_5271)
);

AOI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_5269),
.A2(n_4773),
.B(n_4817),
.Y(n_5272)
);

AOI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_5263),
.A2(n_4812),
.B(n_330),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5248),
.Y(n_5274)
);

OR2x2_ASAP7_75t_L g5275 ( 
.A(n_5266),
.B(n_4809),
.Y(n_5275)
);

NOR3x1_ASAP7_75t_SL g5276 ( 
.A(n_5270),
.B(n_331),
.C(n_332),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_5257),
.B(n_4809),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_5265),
.B(n_4783),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5254),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_5247),
.B(n_331),
.Y(n_5280)
);

AOI311xp33_ASAP7_75t_L g5281 ( 
.A1(n_5262),
.A2(n_332),
.A3(n_333),
.B(n_334),
.C(n_335),
.Y(n_5281)
);

AND2x4_ASAP7_75t_L g5282 ( 
.A(n_5260),
.B(n_335),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_5255),
.Y(n_5283)
);

OR2x2_ASAP7_75t_L g5284 ( 
.A(n_5252),
.B(n_337),
.Y(n_5284)
);

AOI221xp5_ASAP7_75t_L g5285 ( 
.A1(n_5253),
.A2(n_338),
.B1(n_339),
.B2(n_341),
.C(n_342),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5251),
.Y(n_5286)
);

OAI21xp5_ASAP7_75t_L g5287 ( 
.A1(n_5264),
.A2(n_338),
.B(n_339),
.Y(n_5287)
);

AO21x1_ASAP7_75t_L g5288 ( 
.A1(n_5267),
.A2(n_341),
.B(n_344),
.Y(n_5288)
);

NAND4xp75_ASAP7_75t_L g5289 ( 
.A(n_5268),
.B(n_345),
.C(n_347),
.D(n_348),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_5246),
.A2(n_347),
.B(n_349),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_5250),
.Y(n_5291)
);

NOR3x1_ASAP7_75t_L g5292 ( 
.A(n_5249),
.B(n_5256),
.C(n_5261),
.Y(n_5292)
);

NOR3xp33_ASAP7_75t_L g5293 ( 
.A(n_5259),
.B(n_349),
.C(n_352),
.Y(n_5293)
);

NAND3xp33_ASAP7_75t_L g5294 ( 
.A(n_5259),
.B(n_353),
.C(n_354),
.Y(n_5294)
);

INVxp67_ASAP7_75t_L g5295 ( 
.A(n_5258),
.Y(n_5295)
);

NAND4xp25_ASAP7_75t_L g5296 ( 
.A(n_5269),
.B(n_355),
.C(n_356),
.D(n_357),
.Y(n_5296)
);

NAND5xp2_ASAP7_75t_L g5297 ( 
.A(n_5253),
.B(n_356),
.C(n_357),
.D(n_358),
.E(n_359),
.Y(n_5297)
);

NOR3xp33_ASAP7_75t_L g5298 ( 
.A(n_5295),
.B(n_360),
.C(n_361),
.Y(n_5298)
);

OR2x2_ASAP7_75t_L g5299 ( 
.A(n_5297),
.B(n_360),
.Y(n_5299)
);

AND4x1_ASAP7_75t_L g5300 ( 
.A(n_5271),
.B(n_362),
.C(n_363),
.D(n_364),
.Y(n_5300)
);

OAI22xp33_ASAP7_75t_L g5301 ( 
.A1(n_5275),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_5301)
);

NOR4xp25_ASAP7_75t_L g5302 ( 
.A(n_5280),
.B(n_366),
.C(n_368),
.D(n_369),
.Y(n_5302)
);

NAND3xp33_ASAP7_75t_L g5303 ( 
.A(n_5285),
.B(n_368),
.C(n_370),
.Y(n_5303)
);

INVxp33_ASAP7_75t_L g5304 ( 
.A(n_5296),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_5279),
.B(n_5282),
.Y(n_5305)
);

NOR3x1_ASAP7_75t_L g5306 ( 
.A(n_5294),
.B(n_5286),
.C(n_5284),
.Y(n_5306)
);

NOR3xp33_ASAP7_75t_L g5307 ( 
.A(n_5274),
.B(n_5291),
.C(n_5283),
.Y(n_5307)
);

AOI221x1_ASAP7_75t_L g5308 ( 
.A1(n_5293),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.C(n_373),
.Y(n_5308)
);

NAND4xp25_ASAP7_75t_L g5309 ( 
.A(n_5292),
.B(n_372),
.C(n_373),
.D(n_374),
.Y(n_5309)
);

AOI211x1_ASAP7_75t_SL g5310 ( 
.A1(n_5290),
.A2(n_377),
.B(n_378),
.C(n_379),
.Y(n_5310)
);

AOI221xp5_ASAP7_75t_L g5311 ( 
.A1(n_5273),
.A2(n_379),
.B1(n_380),
.B2(n_381),
.C(n_382),
.Y(n_5311)
);

NAND3xp33_ASAP7_75t_L g5312 ( 
.A(n_5281),
.B(n_383),
.C(n_384),
.Y(n_5312)
);

AND4x1_ASAP7_75t_L g5313 ( 
.A(n_5287),
.B(n_5276),
.C(n_5277),
.D(n_5272),
.Y(n_5313)
);

OAI211xp5_ASAP7_75t_L g5314 ( 
.A1(n_5278),
.A2(n_383),
.B(n_384),
.C(n_385),
.Y(n_5314)
);

NOR2x1_ASAP7_75t_L g5315 ( 
.A(n_5289),
.B(n_5282),
.Y(n_5315)
);

O2A1O1Ixp33_ASAP7_75t_SL g5316 ( 
.A1(n_5288),
.A2(n_385),
.B(n_386),
.C(n_387),
.Y(n_5316)
);

NAND4xp25_ASAP7_75t_L g5317 ( 
.A(n_5297),
.B(n_386),
.C(n_388),
.D(n_390),
.Y(n_5317)
);

NAND4xp25_ASAP7_75t_L g5318 ( 
.A(n_5297),
.B(n_388),
.C(n_390),
.D(n_391),
.Y(n_5318)
);

AOI221x1_ASAP7_75t_L g5319 ( 
.A1(n_5279),
.A2(n_392),
.B1(n_394),
.B2(n_396),
.C(n_397),
.Y(n_5319)
);

NOR2x1_ASAP7_75t_L g5320 ( 
.A(n_5289),
.B(n_392),
.Y(n_5320)
);

OAI21xp5_ASAP7_75t_L g5321 ( 
.A1(n_5295),
.A2(n_396),
.B(n_398),
.Y(n_5321)
);

HB1xp67_ASAP7_75t_L g5322 ( 
.A(n_5300),
.Y(n_5322)
);

NOR3x1_ASAP7_75t_L g5323 ( 
.A(n_5312),
.B(n_5309),
.C(n_5303),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_5302),
.B(n_398),
.Y(n_5324)
);

NOR2x1p5_ASAP7_75t_L g5325 ( 
.A(n_5299),
.B(n_399),
.Y(n_5325)
);

INVxp67_ASAP7_75t_L g5326 ( 
.A(n_5315),
.Y(n_5326)
);

AOI21xp5_ASAP7_75t_L g5327 ( 
.A1(n_5305),
.A2(n_399),
.B(n_400),
.Y(n_5327)
);

NAND3x1_ASAP7_75t_SL g5328 ( 
.A(n_5320),
.B(n_400),
.C(n_401),
.Y(n_5328)
);

HB1xp67_ASAP7_75t_L g5329 ( 
.A(n_5319),
.Y(n_5329)
);

OAI322xp33_ASAP7_75t_L g5330 ( 
.A1(n_5301),
.A2(n_401),
.A3(n_402),
.B1(n_403),
.B2(n_404),
.C1(n_406),
.C2(n_408),
.Y(n_5330)
);

AOI222xp33_ASAP7_75t_L g5331 ( 
.A1(n_5304),
.A2(n_406),
.B1(n_411),
.B2(n_412),
.C1(n_413),
.C2(n_414),
.Y(n_5331)
);

AOI211x1_ASAP7_75t_L g5332 ( 
.A1(n_5313),
.A2(n_412),
.B(n_413),
.C(n_415),
.Y(n_5332)
);

HB1xp67_ASAP7_75t_L g5333 ( 
.A(n_5308),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_5298),
.B(n_416),
.Y(n_5334)
);

INVx1_ASAP7_75t_SL g5335 ( 
.A(n_5321),
.Y(n_5335)
);

NOR2xp33_ASAP7_75t_L g5336 ( 
.A(n_5317),
.B(n_5318),
.Y(n_5336)
);

AND2x2_ASAP7_75t_L g5337 ( 
.A(n_5306),
.B(n_417),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_R g5338 ( 
.A1(n_5310),
.A2(n_417),
.B1(n_418),
.B2(n_420),
.Y(n_5338)
);

BUFx6f_ASAP7_75t_L g5339 ( 
.A(n_5307),
.Y(n_5339)
);

INVx3_ASAP7_75t_L g5340 ( 
.A(n_5339),
.Y(n_5340)
);

INVxp33_ASAP7_75t_SL g5341 ( 
.A(n_5322),
.Y(n_5341)
);

NOR2x1_ASAP7_75t_L g5342 ( 
.A(n_5325),
.B(n_5314),
.Y(n_5342)
);

NOR2x1_ASAP7_75t_L g5343 ( 
.A(n_5324),
.B(n_5316),
.Y(n_5343)
);

INVxp67_ASAP7_75t_L g5344 ( 
.A(n_5329),
.Y(n_5344)
);

NOR2xp33_ASAP7_75t_L g5345 ( 
.A(n_5326),
.B(n_5311),
.Y(n_5345)
);

XNOR2xp5_ASAP7_75t_L g5346 ( 
.A(n_5328),
.B(n_418),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5337),
.Y(n_5347)
);

NOR2x1_ASAP7_75t_L g5348 ( 
.A(n_5330),
.B(n_421),
.Y(n_5348)
);

NOR2x1_ASAP7_75t_L g5349 ( 
.A(n_5327),
.B(n_423),
.Y(n_5349)
);

HB1xp67_ASAP7_75t_L g5350 ( 
.A(n_5333),
.Y(n_5350)
);

AND2x2_ASAP7_75t_L g5351 ( 
.A(n_5336),
.B(n_424),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_5332),
.B(n_425),
.Y(n_5352)
);

NAND2x1p5_ASAP7_75t_L g5353 ( 
.A(n_5335),
.B(n_425),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5339),
.B(n_426),
.Y(n_5354)
);

OR2x2_ASAP7_75t_L g5355 ( 
.A(n_5334),
.B(n_426),
.Y(n_5355)
);

NOR4xp25_ASAP7_75t_L g5356 ( 
.A(n_5344),
.B(n_5323),
.C(n_5338),
.D(n_5331),
.Y(n_5356)
);

NOR2xp67_ASAP7_75t_SL g5357 ( 
.A(n_5350),
.B(n_427),
.Y(n_5357)
);

NOR2xp67_ASAP7_75t_L g5358 ( 
.A(n_5346),
.B(n_428),
.Y(n_5358)
);

OR3x2_ASAP7_75t_L g5359 ( 
.A(n_5347),
.B(n_429),
.C(n_430),
.Y(n_5359)
);

INVxp67_ASAP7_75t_SL g5360 ( 
.A(n_5353),
.Y(n_5360)
);

NOR3xp33_ASAP7_75t_L g5361 ( 
.A(n_5340),
.B(n_429),
.C(n_431),
.Y(n_5361)
);

AND2x4_ASAP7_75t_L g5362 ( 
.A(n_5351),
.B(n_431),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_5352),
.Y(n_5363)
);

NOR2xp67_ASAP7_75t_SL g5364 ( 
.A(n_5354),
.B(n_432),
.Y(n_5364)
);

NAND3xp33_ASAP7_75t_SL g5365 ( 
.A(n_5355),
.B(n_433),
.C(n_434),
.Y(n_5365)
);

NOR3xp33_ASAP7_75t_SL g5366 ( 
.A(n_5345),
.B(n_433),
.C(n_434),
.Y(n_5366)
);

NAND4xp25_ASAP7_75t_L g5367 ( 
.A(n_5341),
.B(n_435),
.C(n_436),
.D(n_438),
.Y(n_5367)
);

NOR2x1_ASAP7_75t_L g5368 ( 
.A(n_5343),
.B(n_435),
.Y(n_5368)
);

NAND4xp25_ASAP7_75t_L g5369 ( 
.A(n_5342),
.B(n_439),
.C(n_440),
.D(n_441),
.Y(n_5369)
);

NOR2x1p5_ASAP7_75t_L g5370 ( 
.A(n_5348),
.B(n_439),
.Y(n_5370)
);

NAND4xp25_ASAP7_75t_L g5371 ( 
.A(n_5349),
.B(n_440),
.C(n_444),
.D(n_445),
.Y(n_5371)
);

NOR2x1_ASAP7_75t_L g5372 ( 
.A(n_5343),
.B(n_444),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_5357),
.Y(n_5373)
);

CKINVDCx16_ASAP7_75t_R g5374 ( 
.A(n_5356),
.Y(n_5374)
);

XOR2xp5_ASAP7_75t_L g5375 ( 
.A(n_5359),
.B(n_445),
.Y(n_5375)
);

NOR2xp33_ASAP7_75t_L g5376 ( 
.A(n_5371),
.B(n_447),
.Y(n_5376)
);

INVxp67_ASAP7_75t_L g5377 ( 
.A(n_5362),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5366),
.B(n_447),
.Y(n_5378)
);

AND2x2_ASAP7_75t_L g5379 ( 
.A(n_5370),
.B(n_449),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5368),
.Y(n_5380)
);

HB1xp67_ASAP7_75t_L g5381 ( 
.A(n_5372),
.Y(n_5381)
);

BUFx4f_ASAP7_75t_SL g5382 ( 
.A(n_5363),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_5364),
.Y(n_5383)
);

AOI221x1_ASAP7_75t_L g5384 ( 
.A1(n_5365),
.A2(n_449),
.B1(n_450),
.B2(n_452),
.C(n_453),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5362),
.Y(n_5385)
);

AOI32xp33_ASAP7_75t_L g5386 ( 
.A1(n_5378),
.A2(n_5360),
.A3(n_5361),
.B1(n_5358),
.B2(n_5369),
.Y(n_5386)
);

OAI22x1_ASAP7_75t_SL g5387 ( 
.A1(n_5385),
.A2(n_5367),
.B1(n_452),
.B2(n_455),
.Y(n_5387)
);

AOI221xp5_ASAP7_75t_L g5388 ( 
.A1(n_5376),
.A2(n_450),
.B1(n_455),
.B2(n_456),
.C(n_457),
.Y(n_5388)
);

INVx2_ASAP7_75t_L g5389 ( 
.A(n_5379),
.Y(n_5389)
);

BUFx4f_ASAP7_75t_SL g5390 ( 
.A(n_5373),
.Y(n_5390)
);

AOI322xp5_ASAP7_75t_L g5391 ( 
.A1(n_5374),
.A2(n_457),
.A3(n_459),
.B1(n_460),
.B2(n_461),
.C1(n_462),
.C2(n_463),
.Y(n_5391)
);

AOI322xp5_ASAP7_75t_L g5392 ( 
.A1(n_5383),
.A2(n_460),
.A3(n_462),
.B1(n_464),
.B2(n_466),
.C1(n_468),
.C2(n_469),
.Y(n_5392)
);

OAI22xp5_ASAP7_75t_L g5393 ( 
.A1(n_5390),
.A2(n_5375),
.B1(n_5377),
.B2(n_5382),
.Y(n_5393)
);

AOI22xp5_ASAP7_75t_L g5394 ( 
.A1(n_5387),
.A2(n_5389),
.B1(n_5380),
.B2(n_5381),
.Y(n_5394)
);

AOI22xp5_ASAP7_75t_L g5395 ( 
.A1(n_5388),
.A2(n_5384),
.B1(n_468),
.B2(n_525),
.Y(n_5395)
);

AOI22xp5_ASAP7_75t_L g5396 ( 
.A1(n_5386),
.A2(n_5391),
.B1(n_5392),
.B2(n_528),
.Y(n_5396)
);

AOI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5390),
.A2(n_523),
.B1(n_526),
.B2(n_529),
.Y(n_5397)
);

OAI22xp5_ASAP7_75t_L g5398 ( 
.A1(n_5390),
.A2(n_531),
.B1(n_532),
.B2(n_534),
.Y(n_5398)
);

AOI22xp5_ASAP7_75t_L g5399 ( 
.A1(n_5390),
.A2(n_535),
.B1(n_537),
.B2(n_538),
.Y(n_5399)
);

AOI22xp5_ASAP7_75t_L g5400 ( 
.A1(n_5393),
.A2(n_550),
.B1(n_552),
.B2(n_553),
.Y(n_5400)
);

OAI221xp5_ASAP7_75t_L g5401 ( 
.A1(n_5394),
.A2(n_5395),
.B1(n_5396),
.B2(n_5398),
.C(n_5397),
.Y(n_5401)
);

NOR3xp33_ASAP7_75t_L g5402 ( 
.A(n_5399),
.B(n_555),
.C(n_557),
.Y(n_5402)
);

NAND3xp33_ASAP7_75t_L g5403 ( 
.A(n_5394),
.B(n_563),
.C(n_565),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5395),
.B(n_566),
.Y(n_5404)
);

NAND2xp5_ASAP7_75t_SL g5405 ( 
.A(n_5394),
.B(n_567),
.Y(n_5405)
);

AOI22xp5_ASAP7_75t_L g5406 ( 
.A1(n_5402),
.A2(n_569),
.B1(n_570),
.B2(n_573),
.Y(n_5406)
);

AOI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_5404),
.A2(n_1764),
.B(n_579),
.Y(n_5407)
);

OAI211xp5_ASAP7_75t_SL g5408 ( 
.A1(n_5401),
.A2(n_578),
.B(n_581),
.C(n_586),
.Y(n_5408)
);

AOI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_5405),
.A2(n_587),
.B1(n_588),
.B2(n_591),
.Y(n_5409)
);

INVxp67_ASAP7_75t_L g5410 ( 
.A(n_5403),
.Y(n_5410)
);

AOI22xp5_ASAP7_75t_L g5411 ( 
.A1(n_5408),
.A2(n_5400),
.B1(n_598),
.B2(n_606),
.Y(n_5411)
);

OAI22xp5_ASAP7_75t_L g5412 ( 
.A1(n_5406),
.A2(n_593),
.B1(n_607),
.B2(n_613),
.Y(n_5412)
);

INVx1_ASAP7_75t_SL g5413 ( 
.A(n_5407),
.Y(n_5413)
);

OAI22xp5_ASAP7_75t_L g5414 ( 
.A1(n_5410),
.A2(n_617),
.B1(n_619),
.B2(n_621),
.Y(n_5414)
);

INVx3_ASAP7_75t_L g5415 ( 
.A(n_5413),
.Y(n_5415)
);

AOI21xp33_ASAP7_75t_L g5416 ( 
.A1(n_5411),
.A2(n_5409),
.B(n_625),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_L g5417 ( 
.A(n_5412),
.B(n_622),
.Y(n_5417)
);

AOI221xp5_ASAP7_75t_L g5418 ( 
.A1(n_5414),
.A2(n_627),
.B1(n_629),
.B2(n_636),
.C(n_637),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5411),
.Y(n_5419)
);

AOI21xp5_ASAP7_75t_L g5420 ( 
.A1(n_5419),
.A2(n_1764),
.B(n_1597),
.Y(n_5420)
);

OAI22xp33_ASAP7_75t_L g5421 ( 
.A1(n_5417),
.A2(n_639),
.B1(n_640),
.B2(n_642),
.Y(n_5421)
);

OAI21xp5_ASAP7_75t_SL g5422 ( 
.A1(n_5416),
.A2(n_649),
.B(n_652),
.Y(n_5422)
);

AOI21xp5_ASAP7_75t_L g5423 ( 
.A1(n_5415),
.A2(n_1764),
.B(n_1643),
.Y(n_5423)
);

AO21x1_ASAP7_75t_SL g5424 ( 
.A1(n_5418),
.A2(n_653),
.B(n_655),
.Y(n_5424)
);

OA21x2_ASAP7_75t_L g5425 ( 
.A1(n_5419),
.A2(n_658),
.B(n_1934),
.Y(n_5425)
);

AOI21xp5_ASAP7_75t_L g5426 ( 
.A1(n_5419),
.A2(n_1566),
.B(n_1580),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_L g5427 ( 
.A(n_5415),
.B(n_1566),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_5415),
.B(n_1566),
.Y(n_5428)
);

A2O1A1O1Ixp25_ASAP7_75t_L g5429 ( 
.A1(n_5416),
.A2(n_2513),
.B(n_1934),
.C(n_1927),
.D(n_1596),
.Y(n_5429)
);

AOI22xp33_ASAP7_75t_L g5430 ( 
.A1(n_5424),
.A2(n_1934),
.B1(n_1927),
.B2(n_2513),
.Y(n_5430)
);

AOI22xp33_ASAP7_75t_L g5431 ( 
.A1(n_5427),
.A2(n_1934),
.B1(n_1927),
.B2(n_2513),
.Y(n_5431)
);

AOI22xp5_ASAP7_75t_L g5432 ( 
.A1(n_5422),
.A2(n_1566),
.B1(n_1580),
.B2(n_1582),
.Y(n_5432)
);

OAI22xp5_ASAP7_75t_L g5433 ( 
.A1(n_5428),
.A2(n_1580),
.B1(n_1582),
.B2(n_1596),
.Y(n_5433)
);

OAI22xp5_ASAP7_75t_L g5434 ( 
.A1(n_5426),
.A2(n_1580),
.B1(n_1582),
.B2(n_1596),
.Y(n_5434)
);

AOI22xp5_ASAP7_75t_L g5435 ( 
.A1(n_5425),
.A2(n_1582),
.B1(n_1596),
.B2(n_1597),
.Y(n_5435)
);

OAI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_5429),
.A2(n_1597),
.B(n_1600),
.Y(n_5436)
);

AO22x2_ASAP7_75t_L g5437 ( 
.A1(n_5423),
.A2(n_1597),
.B1(n_1600),
.B2(n_1616),
.Y(n_5437)
);

AOI22xp5_ASAP7_75t_L g5438 ( 
.A1(n_5425),
.A2(n_1600),
.B1(n_1616),
.B2(n_1622),
.Y(n_5438)
);

AOI22xp5_ASAP7_75t_L g5439 ( 
.A1(n_5421),
.A2(n_1600),
.B1(n_1616),
.B2(n_1622),
.Y(n_5439)
);

INVxp67_ASAP7_75t_L g5440 ( 
.A(n_5432),
.Y(n_5440)
);

XOR2xp5_ASAP7_75t_L g5441 ( 
.A(n_5439),
.B(n_5420),
.Y(n_5441)
);

AO21x2_ASAP7_75t_L g5442 ( 
.A1(n_5436),
.A2(n_1616),
.B(n_1622),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_5434),
.A2(n_1622),
.B(n_1625),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_5435),
.B(n_1625),
.Y(n_5444)
);

AOI21xp33_ASAP7_75t_L g5445 ( 
.A1(n_5433),
.A2(n_1625),
.B(n_1643),
.Y(n_5445)
);

OAI22xp5_ASAP7_75t_L g5446 ( 
.A1(n_5438),
.A2(n_1625),
.B1(n_1643),
.B2(n_1650),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_5437),
.B(n_1643),
.Y(n_5447)
);

AOI22xp5_ASAP7_75t_SL g5448 ( 
.A1(n_5440),
.A2(n_5430),
.B1(n_5431),
.B2(n_1664),
.Y(n_5448)
);

HB1xp67_ASAP7_75t_L g5449 ( 
.A(n_5442),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5441),
.Y(n_5450)
);

OAI22xp33_ASAP7_75t_L g5451 ( 
.A1(n_5444),
.A2(n_5447),
.B1(n_5446),
.B2(n_5443),
.Y(n_5451)
);

AOI221x1_ASAP7_75t_L g5452 ( 
.A1(n_5450),
.A2(n_5445),
.B1(n_1661),
.B2(n_1664),
.C(n_1667),
.Y(n_5452)
);

AOI21xp5_ASAP7_75t_L g5453 ( 
.A1(n_5452),
.A2(n_5451),
.B(n_5449),
.Y(n_5453)
);

AOI211xp5_ASAP7_75t_L g5454 ( 
.A1(n_5453),
.A2(n_5448),
.B(n_1661),
.C(n_1664),
.Y(n_5454)
);


endmodule