module fake_jpeg_12665_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx6f_ASAP7_75t_SL g74 ( 
.A(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_82),
.B(n_69),
.Y(n_101)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_5),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_6),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_52),
.B1(n_77),
.B2(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_92),
.B1(n_102),
.B2(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_65),
.B1(n_54),
.B2(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_58),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_73),
.B(n_53),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_101),
.A2(n_6),
.B(n_7),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_77),
.B1(n_56),
.B2(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_55),
.Y(n_103)
);

CKINVDCx10_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_98),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_111),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_75),
.C(n_68),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_116),
.Y(n_148)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_81),
.B1(n_56),
.B2(n_49),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_10),
.B(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_122),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_60),
.C(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_27),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_25),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_126),
.B(n_59),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_63),
.B(n_62),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_9),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_66),
.B1(n_59),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_134),
.B1(n_140),
.B2(n_145),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_66),
.B1(n_51),
.B2(n_11),
.Y(n_134)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_9),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_139),
.C(n_42),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_12),
.B(n_13),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_22),
.B(n_24),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_35),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_157),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_148),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_162),
.B(n_163),
.Y(n_170)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_148),
.C(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_171),
.C(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_127),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_156),
.B(n_139),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_150),
.B1(n_164),
.B2(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_173),
.A2(n_174),
.B(n_141),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_170),
.C(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

AOI21x1_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_166),
.B(n_136),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_154),
.C(n_131),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_162),
.Y(n_182)
);


endmodule