module fake_jpeg_31889_n_243 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_243);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_243;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_37),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_34),
.C(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_65),
.C(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_23),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_18),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_15),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_20),
.B1(n_33),
.B2(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_20),
.B1(n_22),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_67),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_22),
.B1(n_17),
.B2(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_78),
.Y(n_109)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_21),
.B(n_31),
.C(n_29),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_95),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_99),
.B1(n_105),
.B2(n_63),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_15),
.B1(n_22),
.B2(n_28),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_96),
.B1(n_70),
.B2(n_71),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_50),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_22),
.B1(n_16),
.B2(n_28),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_31),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_106),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_30),
.B1(n_16),
.B2(n_22),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_14),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_100),
.B(n_13),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_68),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_2),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_111),
.B(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_67),
.B1(n_79),
.B2(n_63),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_133),
.B1(n_83),
.B2(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_97),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_128),
.Y(n_165)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_114),
.Y(n_158)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_110),
.B1(n_91),
.B2(n_83),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_3),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_52),
.B(n_5),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_129),
.B(n_9),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_4),
.B(n_5),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_11),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_4),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_7),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_8),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_9),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_9),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_142),
.B(n_144),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_110),
.B(n_91),
.C(n_105),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_165),
.B(n_145),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_152),
.B1(n_160),
.B2(n_164),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_131),
.C(n_120),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_91),
.B1(n_83),
.B2(n_81),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_94),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_82),
.B(n_87),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_135),
.B(n_121),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_133),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_89),
.B1(n_11),
.B2(n_10),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_87),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_113),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_139),
.B1(n_112),
.B2(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_119),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_180),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_149),
.B1(n_167),
.B2(n_171),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_127),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_130),
.C(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_171),
.B(n_173),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_129),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_174),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_125),
.B(n_126),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_114),
.C(n_115),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_116),
.C(n_121),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_152),
.B1(n_147),
.B2(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_192),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_150),
.B1(n_164),
.B2(n_160),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_172),
.B1(n_181),
.B2(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_198),
.B(n_190),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_203),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_183),
.B1(n_180),
.B2(n_159),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_191),
.B1(n_195),
.B2(n_187),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_170),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_209),
.Y(n_213)
);

OA21x2_ASAP7_75t_SL g207 ( 
.A1(n_189),
.A2(n_175),
.B(n_146),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_198),
.B(n_190),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_182),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_187),
.Y(n_216)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_212),
.A2(n_192),
.B1(n_194),
.B2(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_206),
.B1(n_208),
.B2(n_212),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_221),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_220),
.B1(n_206),
.B2(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_184),
.C(n_146),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_227),
.Y(n_231)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_205),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_188),
.B1(n_196),
.B2(n_157),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_228),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_218),
.C(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_188),
.B(n_213),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_224),
.B1(n_217),
.B2(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_213),
.B1(n_222),
.B2(n_176),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_233),
.B(n_222),
.C(n_174),
.Y(n_237)
);

NOR4xp25_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_234),
.C(n_236),
.D(n_141),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.C(n_151),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_143),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_241),
.A2(n_143),
.B1(n_161),
.B2(n_156),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_161),
.Y(n_243)
);


endmodule