module real_aes_11366_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_56;
wire n_34;
wire n_55;
wire n_12;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_54;
wire n_51;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g28 ( .A(n_1), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_2), .B(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_2), .Y(n_37) );
BUFx2_ASAP7_75t_L g45 ( .A(n_3), .Y(n_45) );
INVx1_ASAP7_75t_L g19 ( .A(n_4), .Y(n_19) );
INVx1_ASAP7_75t_L g40 ( .A(n_5), .Y(n_40) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_6), .Y(n_24) );
INVx2_ASAP7_75t_L g31 ( .A(n_7), .Y(n_31) );
BUFx10_ASAP7_75t_L g47 ( .A(n_8), .Y(n_47) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_15), .Y(n_14) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_20), .B1(n_32), .B2(n_46), .C(n_48), .Y(n_10) );
BUFx2_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_13), .B(n_17), .Y(n_12) );
HB1xp67_ASAP7_75t_L g55 ( .A(n_13), .Y(n_55) );
INVx1_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
HB1xp67_ASAP7_75t_L g38 ( .A(n_19), .Y(n_38) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_21), .B(n_25), .Y(n_20) );
INVxp67_ASAP7_75t_L g56 ( .A(n_21), .Y(n_56) );
INVxp67_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
CKINVDCx20_ASAP7_75t_R g49 ( .A(n_25), .Y(n_49) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_26), .B(n_29), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
INVx1_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
CKINVDCx16_ASAP7_75t_R g32 ( .A(n_33), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_34), .B(n_39), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_36), .B(n_38), .Y(n_35) );
HB1xp67_ASAP7_75t_L g50 ( .A(n_36), .Y(n_50) );
INVx1_ASAP7_75t_L g36 ( .A(n_37), .Y(n_36) );
INVx1_ASAP7_75t_SL g52 ( .A(n_38), .Y(n_52) );
OAI22xp33_ASAP7_75t_SL g53 ( .A1(n_39), .A2(n_50), .B1(n_54), .B2(n_55), .Y(n_53) );
NOR2xp33_ASAP7_75t_L g39 ( .A(n_40), .B(n_41), .Y(n_39) );
INVx5_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
BUFx8_ASAP7_75t_SL g42 ( .A(n_43), .Y(n_42) );
INVx2_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
BUFx2_ASAP7_75t_L g44 ( .A(n_45), .Y(n_44) );
BUFx12f_ASAP7_75t_L g46 ( .A(n_47), .Y(n_46) );
O2A1O1Ixp33_ASAP7_75t_SL g48 ( .A1(n_49), .A2(n_50), .B(n_51), .C(n_56), .Y(n_48) );
CKINVDCx20_ASAP7_75t_R g54 ( .A(n_50), .Y(n_54) );
NOR2xp33_ASAP7_75t_L g51 ( .A(n_52), .B(n_53), .Y(n_51) );
endmodule