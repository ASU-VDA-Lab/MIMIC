module fake_jpeg_21615_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_45),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_27),
.B1(n_24),
.B2(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_73),
.B1(n_26),
.B2(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_29),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_35),
.Y(n_55)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_60),
.CI(n_37),
.CON(n_98),
.SN(n_98)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_27),
.B1(n_16),
.B2(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_22),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_35),
.C(n_27),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_25),
.C(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_17),
.B1(n_43),
.B2(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_30),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_19),
.B(n_30),
.C(n_24),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_92),
.A3(n_108),
.B1(n_32),
.B2(n_40),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_59),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_78),
.Y(n_129)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_83),
.A2(n_23),
.B1(n_32),
.B2(n_17),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_87),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_20),
.B1(n_31),
.B2(n_21),
.Y(n_85)
);

OAI22x1_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_40),
.B1(n_34),
.B2(n_39),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_47),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_35),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_21),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_47),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_64),
.B(n_55),
.C(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_109),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_102),
.Y(n_140)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_101),
.Y(n_139)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_39),
.B1(n_20),
.B2(n_17),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_30),
.B(n_33),
.C(n_23),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_26),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_40),
.C(n_18),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_34),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_39),
.C(n_37),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_144),
.C(n_0),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_79),
.B1(n_91),
.B2(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_126),
.B1(n_130),
.B2(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_112),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_89),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_107),
.B1(n_88),
.B2(n_106),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_82),
.A2(n_71),
.B1(n_17),
.B2(n_42),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_71),
.B1(n_17),
.B2(n_42),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_77),
.A2(n_20),
.B1(n_32),
.B2(n_40),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_126),
.B1(n_130),
.B2(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_80),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_143),
.B1(n_76),
.B2(n_108),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_110),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_20),
.B1(n_40),
.B2(n_34),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_157),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_94),
.B1(n_89),
.B2(n_84),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_156),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_138),
.B1(n_140),
.B2(n_137),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_96),
.B(n_34),
.C(n_97),
.D(n_105),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_150),
.A2(n_155),
.B(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_96),
.B(n_94),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_161),
.B(n_129),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_34),
.B(n_28),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_84),
.B1(n_104),
.B2(n_102),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_160),
.B(n_167),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_34),
.B(n_28),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_103),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_81),
.B1(n_101),
.B2(n_103),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_132),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_171),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_29),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_34),
.B1(n_18),
.B2(n_28),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_18),
.B1(n_28),
.B2(n_110),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_18),
.B1(n_7),
.B2(n_9),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_127),
.B1(n_136),
.B2(n_139),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_125),
.B(n_6),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_177),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_172),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_132),
.B(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_15),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_178),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_143),
.C(n_115),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_182),
.C(n_188),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_192),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_135),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_206),
.B(n_161),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_115),
.C(n_136),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_209),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_139),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_157),
.B1(n_173),
.B2(n_155),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_145),
.B(n_128),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_210),
.C(n_166),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_0),
.B(n_1),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_12),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_146),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_11),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_149),
.B1(n_153),
.B2(n_150),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_228),
.B1(n_232),
.B2(n_193),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_182),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_225),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_174),
.B(n_170),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_170),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_152),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_162),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_10),
.B(n_3),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_183),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_2),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_191),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_239),
.B(n_253),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_246),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_179),
.C(n_188),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_249),
.C(n_254),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_256),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_195),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_184),
.C(n_210),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_194),
.C(n_180),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_183),
.B1(n_193),
.B2(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_180),
.C(n_192),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_237),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AO22x1_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_226),
.B1(n_227),
.B2(n_222),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_225),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_229),
.B(n_230),
.C(n_218),
.D(n_204),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_243),
.C(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_230),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_240),
.A2(n_201),
.B1(n_211),
.B2(n_228),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_276),
.B1(n_277),
.B2(n_231),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_272),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_SL g271 ( 
.A(n_243),
.B(n_244),
.C(n_238),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_274),
.B(n_275),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_248),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_252),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_220),
.B1(n_214),
.B2(n_219),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_242),
.C(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_281),
.C(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_5),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_SL g280 ( 
.A1(n_264),
.A2(n_223),
.A3(n_187),
.B1(n_249),
.B2(n_254),
.C1(n_190),
.C2(n_233),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_291),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_257),
.C(n_256),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_245),
.C(n_224),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_185),
.B1(n_186),
.B2(n_3),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_236),
.C(n_235),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_263),
.C(n_266),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_185),
.B1(n_223),
.B2(n_186),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_276),
.B1(n_275),
.B2(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_288),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_304),
.B1(n_292),
.B2(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_270),
.C(n_260),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_303),
.B(n_5),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_265),
.C(n_271),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_5),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_5),
.B1(n_289),
.B2(n_284),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_310),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_279),
.B(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_294),
.C(n_293),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_316),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_307),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_294),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_315),
.C(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.C(n_320),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_310),
.B(n_314),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_324),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_309),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);


endmodule