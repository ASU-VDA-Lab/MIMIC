module real_jpeg_24282_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_80),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_170),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_1),
.A2(n_65),
.B1(n_67),
.B2(n_170),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_1),
.A2(n_54),
.B1(n_60),
.B2(n_170),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_22),
.B1(n_27),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_3),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_65),
.B1(n_67),
.B2(n_95),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_30),
.B1(n_40),
.B2(n_95),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_3),
.A2(n_54),
.B1(n_60),
.B2(n_95),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_39),
.B1(n_65),
.B2(n_67),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_39),
.B1(n_54),
.B2(n_60),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_39),
.Y(n_137)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_9),
.A2(n_30),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_81),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_9),
.A2(n_65),
.B1(n_67),
.B2(n_81),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_54),
.B1(n_60),
.B2(n_81),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_31),
.B1(n_35),
.B2(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_22),
.B1(n_27),
.B2(n_85),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_65),
.B1(n_67),
.B2(n_85),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_10),
.A2(n_54),
.B1(n_60),
.B2(n_85),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_171),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_21),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_65),
.C(n_91),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_224),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_11),
.B(n_135),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_11),
.A2(n_65),
.B1(n_67),
.B2(n_224),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_54),
.C(n_70),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_11),
.A2(n_53),
.B(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_12),
.A2(n_31),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_12),
.A2(n_22),
.B1(n_27),
.B2(n_119),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_12),
.A2(n_65),
.B1(n_67),
.B2(n_119),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_12),
.A2(n_54),
.B1(n_60),
.B2(n_119),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_14),
.A2(n_34),
.B1(n_54),
.B2(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_34),
.B1(n_65),
.B2(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_14),
.A2(n_22),
.B1(n_27),
.B2(n_34),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_15),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_15),
.A2(n_64),
.B1(n_120),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_15),
.A2(n_54),
.B1(n_60),
.B2(n_64),
.Y(n_179)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_28),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_21),
.A2(n_28),
.B1(n_118),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_21),
.A2(n_28),
.B1(n_38),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_22),
.A2(n_27),
.B1(n_91),
.B2(n_92),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_22),
.B(n_26),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_22),
.B(n_249),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_27),
.A3(n_154),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_28),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_28),
.A2(n_123),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_30),
.Y(n_154)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_79),
.B(n_82),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_32),
.B(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_32),
.A2(n_79),
.B1(n_121),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_32),
.A2(n_121),
.B1(n_143),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_32),
.A2(n_82),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_37),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_37),
.B(n_355),
.Y(n_356)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_354),
.B(n_356),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_342),
.B(n_353),
.Y(n_46)
);

OAI31xp33_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_145),
.A3(n_160),
.B(n_339),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_124),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_49),
.B(n_124),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_86),
.C(n_102),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_50),
.A2(n_86),
.B1(n_87),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_50),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_75),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_51),
.A2(n_52),
.B(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_52),
.A2(n_61),
.B1(n_62),
.B2(n_76),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_53),
.A2(n_59),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_53),
.A2(n_56),
.B1(n_107),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_53),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_53),
.A2(n_198),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_53),
.B(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_53),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_60),
.B1(n_70),
.B2(n_71),
.Y(n_72)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_55),
.Y(n_201)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_55),
.Y(n_284)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_58),
.B(n_224),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_60),
.B(n_307),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_73),
.B2(n_74),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_68),
.B1(n_74),
.B2(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_67),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_65),
.B(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_68),
.A2(n_74),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_68),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_68),
.A2(n_74),
.B1(n_255),
.B2(n_257),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_72),
.A2(n_98),
.B1(n_113),
.B2(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_72),
.A2(n_181),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_72),
.A2(n_220),
.B(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_72),
.B(n_224),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_74),
.B(n_221),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_97),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_96),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_89),
.A2(n_90),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_89),
.A2(n_188),
.B(n_190),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_89),
.A2(n_190),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_90),
.A2(n_115),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_90),
.A2(n_174),
.B(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_98),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_98),
.A2(n_271),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_102),
.A2(n_103),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_114),
.C(n_116),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_104),
.A2(n_105),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_109),
.A2(n_196),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_114),
.B(n_116),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B(n_122),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_127),
.C(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_142),
.B2(n_144),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_139),
.C(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_134),
.A2(n_135),
.B1(n_189),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_134),
.A2(n_135),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_135),
.B(n_175),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_139),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_139),
.B(n_152),
.C(n_157),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_144),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_142),
.B(n_148),
.C(n_151),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_146),
.A2(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_159),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_147),
.B(n_159),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_153),
.Y(n_349)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_154),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_158),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_332),
.B(n_338),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_209),
.B(n_331),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_202),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_163),
.B(n_202),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_182),
.C(n_184),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_164),
.A2(n_165),
.B1(n_182),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_173),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_172),
.C(n_176),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_177),
.B(n_180),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_182),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_184),
.B(n_328),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_191),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_185),
.B(n_187),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_191),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_195),
.Y(n_226)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_199),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_337)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_241),
.B(n_325),
.C(n_330),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_235),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.C(n_227),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_212),
.A2(n_213),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.C(n_222),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_226),
.B(n_227),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_232),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_265),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_234),
.A2(n_296),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_319),
.B(n_324),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_272),
.B(n_318),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_261),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_246),
.B(n_261),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_254),
.C(n_258),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_247),
.B(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_254),
.A2(n_258),
.B1(n_259),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_312),
.B(n_317),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_292),
.B(n_311),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_286),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_286),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_300),
.B(n_310),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_298),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_305),
.B(n_309),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_337),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_344),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_346),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_348),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_350),
.C(n_352),
.Y(n_355)
);


endmodule