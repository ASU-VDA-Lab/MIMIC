module fake_jpeg_4299_n_68 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

HB1xp67_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_20),
.Y(n_22)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_17),
.Y(n_26)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_19),
.B(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_31),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_14),
.Y(n_37)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_14),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_28),
.Y(n_38)
);

A2O1A1O1Ixp25_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_42),
.B(n_25),
.C(n_10),
.D(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_28),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

AO221x1_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_24),
.B1(n_21),
.B2(n_16),
.C(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_9),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_25),
.B(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_12),
.B1(n_11),
.B2(n_24),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_11),
.C(n_15),
.Y(n_53)
);

FAx1_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_51),
.CI(n_53),
.CON(n_55),
.SN(n_55)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_44),
.B1(n_24),
.B2(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_16),
.B1(n_9),
.B2(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_3),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_3),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.Y(n_63)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_56),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_65),
.C(n_58),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_55),
.C(n_5),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_7),
.Y(n_68)
);


endmodule