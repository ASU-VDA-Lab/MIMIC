module real_aes_7292_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g449 ( .A(n_0), .Y(n_449) );
INVx1_ASAP7_75t_L g479 ( .A(n_1), .Y(n_479) );
INVx1_ASAP7_75t_L g193 ( .A(n_2), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_3), .A2(n_38), .B1(n_154), .B2(n_509), .Y(n_524) );
AOI21xp33_ASAP7_75t_L g161 ( .A1(n_4), .A2(n_135), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_5), .B(n_128), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_6), .A2(n_100), .B1(n_111), .B2(n_765), .Y(n_99) );
AND2x6_ASAP7_75t_L g140 ( .A(n_7), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_8), .A2(n_243), .B(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_9), .B(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g168 ( .A(n_10), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_11), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
INVx1_ASAP7_75t_L g473 ( .A(n_13), .Y(n_473) );
INVx1_ASAP7_75t_L g249 ( .A(n_14), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_15), .B(n_176), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_16), .B(n_129), .Y(n_550) );
AO32x2_ASAP7_75t_L g522 ( .A1(n_17), .A2(n_128), .A3(n_173), .B1(n_501), .B2(n_523), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_18), .A2(n_118), .B1(n_119), .B2(n_444), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_19), .B(n_154), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_20), .B(n_149), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_21), .B(n_129), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_22), .A2(n_50), .B1(n_154), .B2(n_509), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_23), .B(n_135), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_24), .A2(n_75), .B1(n_154), .B2(n_176), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_25), .B(n_154), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_26), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_27), .A2(n_247), .B(n_248), .C(n_250), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_28), .Y(n_452) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_29), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_30), .B(n_170), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_31), .B(n_166), .Y(n_195) );
INVx1_ASAP7_75t_L g182 ( .A(n_32), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_33), .B(n_170), .Y(n_539) );
INVx2_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_35), .B(n_154), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_36), .B(n_170), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_37), .A2(n_140), .B(n_144), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g180 ( .A(n_40), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_41), .B(n_166), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_42), .B(n_154), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_43), .A2(n_85), .B1(n_212), .B2(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_44), .B(n_154), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_45), .B(n_154), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_46), .Y(n_183) );
OAI222xp33_ASAP7_75t_L g454 ( .A1(n_47), .A2(n_455), .B1(n_752), .B2(n_753), .C1(n_758), .C2(n_762), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g752 ( .A(n_47), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_48), .B(n_478), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_49), .B(n_135), .Y(n_237) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_51), .A2(n_60), .B1(n_154), .B2(n_176), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_52), .A2(n_144), .B1(n_176), .B2(n_178), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_53), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_54), .B(n_154), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_55), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_56), .B(n_154), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_57), .A2(n_153), .B(n_165), .C(n_167), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_58), .Y(n_225) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_62), .B(n_154), .Y(n_480) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
AO32x2_ASAP7_75t_L g506 ( .A1(n_65), .A2(n_128), .A3(n_229), .B1(n_501), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g499 ( .A(n_66), .Y(n_499) );
INVx1_ASAP7_75t_L g534 ( .A(n_67), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_68), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_SL g148 ( .A1(n_69), .A2(n_149), .B(n_150), .C(n_153), .Y(n_148) );
INVxp67_ASAP7_75t_L g151 ( .A(n_70), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_71), .B(n_176), .Y(n_535) );
INVx1_ASAP7_75t_L g108 ( .A(n_72), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_73), .Y(n_186) );
INVx1_ASAP7_75t_L g218 ( .A(n_74), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_76), .A2(n_140), .B(n_144), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_77), .B(n_509), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_78), .B(n_176), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_79), .B(n_194), .Y(n_208) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_81), .B(n_149), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_82), .B(n_176), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_83), .A2(n_140), .B(n_144), .C(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g105 ( .A(n_84), .Y(n_105) );
OR2x2_ASAP7_75t_L g446 ( .A(n_84), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g457 ( .A(n_84), .B(n_448), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_86), .A2(n_98), .B1(n_176), .B2(n_177), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_87), .B(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_88), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_89), .A2(n_140), .B(n_144), .C(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_90), .Y(n_239) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_92), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_93), .B(n_194), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_94), .B(n_176), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_95), .B(n_128), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_97), .A2(n_135), .B(n_142), .Y(n_134) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_102), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_109), .Y(n_103) );
OR2x2_ASAP7_75t_L g460 ( .A(n_105), .B(n_448), .Y(n_460) );
NOR2x2_ASAP7_75t_L g761 ( .A(n_105), .B(n_447), .Y(n_761) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g448 ( .A(n_110), .B(n_449), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_453), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g764 ( .A(n_114), .Y(n_764) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_445), .B(n_450), .Y(n_116) );
INVx2_ASAP7_75t_L g444 ( .A(n_119), .Y(n_444) );
INVx1_ASAP7_75t_SL g458 ( .A(n_119), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_119), .A2(n_754), .B1(n_756), .B2(n_757), .Y(n_753) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND4x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_362), .C(n_409), .D(n_429), .Y(n_120) );
NOR3xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_292), .C(n_317), .Y(n_121) );
OAI211xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_200), .B(n_252), .C(n_282), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_171), .Y(n_124) );
INVx3_ASAP7_75t_SL g334 ( .A(n_125), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_125), .B(n_265), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_125), .B(n_187), .Y(n_415) );
AND2x2_ASAP7_75t_L g438 ( .A(n_125), .B(n_304), .Y(n_438) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_159), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g256 ( .A(n_127), .B(n_160), .Y(n_256) );
INVx3_ASAP7_75t_L g269 ( .A(n_127), .Y(n_269) );
AND2x2_ASAP7_75t_L g274 ( .A(n_127), .B(n_159), .Y(n_274) );
OR2x2_ASAP7_75t_L g325 ( .A(n_127), .B(n_266), .Y(n_325) );
BUFx2_ASAP7_75t_L g345 ( .A(n_127), .Y(n_345) );
AND2x2_ASAP7_75t_L g355 ( .A(n_127), .B(n_266), .Y(n_355) );
AND2x2_ASAP7_75t_L g361 ( .A(n_127), .B(n_172), .Y(n_361) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_156), .Y(n_127) );
INVx4_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_128), .A2(n_485), .B(n_492), .Y(n_484) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_130), .B(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g243 ( .A(n_135), .Y(n_243) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_136), .B(n_140), .Y(n_184) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g478 ( .A(n_137), .Y(n_478) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g145 ( .A(n_138), .Y(n_145) );
INVx1_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
INVx1_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
INVx1_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
INVx4_ASAP7_75t_SL g155 ( .A(n_140), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_140), .A2(n_472), .B(n_476), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_140), .A2(n_486), .B(n_489), .Y(n_485) );
BUFx3_ASAP7_75t_L g501 ( .A(n_140), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_140), .A2(n_514), .B(n_518), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_140), .A2(n_533), .B(n_536), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_148), .C(n_155), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_155), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_143), .A2(n_155), .B(n_245), .C(n_246), .Y(n_244) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_145), .Y(n_154) );
BUFx3_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
INVx1_ASAP7_75t_L g509 ( .A(n_145), .Y(n_509) );
INVx1_ASAP7_75t_L g517 ( .A(n_149), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_152), .B(n_168), .Y(n_167) );
INVx5_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g507 ( .A1(n_152), .A2(n_166), .B1(n_508), .B2(n_510), .Y(n_507) );
O2A1O1Ixp5_ASAP7_75t_SL g533 ( .A1(n_153), .A2(n_194), .B(n_534), .C(n_535), .Y(n_533) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_154), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_155), .A2(n_175), .B1(n_183), .B2(n_184), .Y(n_174) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_157), .A2(n_161), .B(n_169), .Y(n_160) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_158), .B(n_215), .Y(n_214) );
AO21x1_ASAP7_75t_L g545 ( .A1(n_158), .A2(n_546), .B(n_549), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_158), .B(n_501), .C(n_546), .Y(n_564) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_160), .B(n_266), .Y(n_280) );
INVx2_ASAP7_75t_L g290 ( .A(n_160), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_160), .B(n_269), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_160), .B(n_266), .Y(n_314) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_160), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g372 ( .A(n_160), .Y(n_372) );
AND2x2_ASAP7_75t_L g418 ( .A(n_160), .B(n_172), .Y(n_418) );
O2A1O1Ixp5_ASAP7_75t_L g498 ( .A1(n_165), .A2(n_477), .B(n_499), .C(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_165), .A2(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx4_ASAP7_75t_L g235 ( .A(n_166), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_166), .A2(n_481), .B1(n_524), .B2(n_525), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_166), .A2(n_481), .B1(n_547), .B2(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
INVx2_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_170), .A2(n_242), .B(n_251), .Y(n_241) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_170), .A2(n_513), .B(n_521), .Y(n_512) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_170), .A2(n_532), .B(n_539), .Y(n_531) );
INVx3_ASAP7_75t_SL g291 ( .A(n_171), .Y(n_291) );
OR2x2_ASAP7_75t_L g344 ( .A(n_171), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_187), .Y(n_171) );
INVx3_ASAP7_75t_L g266 ( .A(n_172), .Y(n_266) );
AND2x2_ASAP7_75t_L g333 ( .A(n_172), .B(n_188), .Y(n_333) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_172), .Y(n_401) );
AOI33xp33_ASAP7_75t_L g405 ( .A1(n_172), .A2(n_334), .A3(n_341), .B1(n_350), .B2(n_406), .B3(n_407), .Y(n_405) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_173), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_189), .B(n_197), .Y(n_188) );
INVx2_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
INVx2_ASAP7_75t_L g196 ( .A(n_176), .Y(n_196) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_181), .B2(n_182), .Y(n_178) );
INVx2_ASAP7_75t_L g181 ( .A(n_179), .Y(n_181) );
INVx4_ASAP7_75t_L g247 ( .A(n_179), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_184), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_187), .B(n_269), .Y(n_268) );
NOR3xp33_ASAP7_75t_L g328 ( .A(n_187), .B(n_329), .C(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g354 ( .A(n_187), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_187), .B(n_361), .Y(n_364) );
AND2x2_ASAP7_75t_L g417 ( .A(n_187), .B(n_418), .Y(n_417) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g273 ( .A(n_188), .Y(n_273) );
OR2x2_ASAP7_75t_L g367 ( .A(n_188), .B(n_266), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g481 ( .A(n_194), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_194), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_194), .A2(n_496), .B(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_196), .A2(n_473), .B(n_474), .C(n_475), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_199), .B(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_199), .B(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_226), .Y(n_200) );
AOI32xp33_ASAP7_75t_L g318 ( .A1(n_201), .A2(n_319), .A3(n_321), .B1(n_323), .B2(n_326), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_201), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g421 ( .A(n_201), .Y(n_421) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g353 ( .A(n_202), .B(n_337), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_202), .B(n_299), .Y(n_373) );
AND2x2_ASAP7_75t_L g441 ( .A(n_202), .B(n_359), .Y(n_441) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
INVx3_ASAP7_75t_L g262 ( .A(n_203), .Y(n_262) );
AND2x2_ASAP7_75t_L g276 ( .A(n_203), .B(n_260), .Y(n_276) );
OR2x2_ASAP7_75t_L g281 ( .A(n_203), .B(n_259), .Y(n_281) );
INVx1_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
AND2x2_ASAP7_75t_L g296 ( .A(n_203), .B(n_270), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_203), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g351 ( .A(n_203), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_203), .B(n_436), .Y(n_435) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_213), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g250 ( .A(n_212), .Y(n_250) );
INVx1_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_213), .A2(n_471), .B(n_482), .Y(n_470) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_213), .A2(n_494), .B(n_502), .Y(n_493) );
INVx2_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
AND2x2_ASAP7_75t_L g306 ( .A(n_216), .B(n_227), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_216), .B(n_241), .Y(n_316) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_223), .B(n_224), .Y(n_216) );
INVx2_ASAP7_75t_L g436 ( .A(n_226), .Y(n_436) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_227), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
AND2x2_ASAP7_75t_L g321 ( .A(n_227), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g337 ( .A(n_227), .B(n_300), .Y(n_337) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_228), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g350 ( .A(n_228), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_228), .B(n_260), .Y(n_382) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_238), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_237), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
AND2x2_ASAP7_75t_L g261 ( .A(n_240), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g322 ( .A(n_240), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_240), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g359 ( .A(n_240), .Y(n_359) );
INVx1_ASAP7_75t_L g392 ( .A(n_240), .Y(n_392) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_241), .B(n_260), .Y(n_270) );
INVx1_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_247), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g475 ( .A(n_247), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_247), .A2(n_537), .B(n_538), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_257), .B1(n_263), .B2(n_270), .C(n_271), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_254), .B(n_274), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_254), .B(n_337), .Y(n_414) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_256), .B(n_304), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_256), .B(n_265), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_256), .B(n_279), .Y(n_408) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g330 ( .A(n_260), .Y(n_330) );
AND2x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
AND2x2_ASAP7_75t_L g315 ( .A(n_262), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_262), .B(n_285), .Y(n_331) );
AND2x2_ASAP7_75t_L g395 ( .A(n_262), .B(n_321), .Y(n_395) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g304 ( .A(n_266), .B(n_273), .Y(n_304) );
AND2x2_ASAP7_75t_L g400 ( .A(n_267), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_269), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_270), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_270), .B(n_277), .Y(n_365) );
AND2x2_ASAP7_75t_L g385 ( .A(n_270), .B(n_285), .Y(n_385) );
AND2x2_ASAP7_75t_L g406 ( .A(n_270), .B(n_350), .Y(n_406) );
OAI32xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_275), .A3(n_277), .B1(n_278), .B2(n_281), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g279 ( .A(n_273), .Y(n_279) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_273), .B(n_303), .Y(n_320) );
OR2x2_ASAP7_75t_L g324 ( .A(n_273), .B(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_273), .B(n_372), .Y(n_425) );
INVx1_ASAP7_75t_L g293 ( .A(n_274), .Y(n_293) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_275), .A2(n_366), .B1(n_412), .B2(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g283 ( .A(n_276), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g326 ( .A(n_276), .B(n_299), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_276), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g404 ( .A(n_276), .B(n_337), .Y(n_404) );
INVxp67_ASAP7_75t_L g340 ( .A(n_277), .Y(n_340) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g410 ( .A(n_279), .B(n_397), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_279), .B(n_360), .Y(n_433) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_281), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g426 ( .A(n_281), .B(n_427), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_286), .B(n_289), .Y(n_282) );
AND2x2_ASAP7_75t_L g295 ( .A(n_284), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g379 ( .A(n_288), .B(n_299), .Y(n_379) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g397 ( .A(n_290), .B(n_355), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_290), .B(n_354), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_291), .B(n_303), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_297), .C(n_307), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_293), .A2(n_328), .B1(n_332), .B2(n_335), .C(n_338), .Y(n_327) );
AOI31xp33_ASAP7_75t_L g422 ( .A1(n_293), .A2(n_423), .A3(n_424), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_303), .B2(n_305), .Y(n_297) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g423 ( .A(n_303), .Y(n_423) );
INVx1_ASAP7_75t_L g386 ( .A(n_304), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_306), .A2(n_430), .B(n_432), .C(n_434), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_311), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_312), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_314), .A2(n_348), .B1(n_367), .B2(n_403), .C(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g398 ( .A(n_315), .Y(n_398) );
INVx1_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g317 ( .A(n_318), .B(n_327), .C(n_342), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_319), .A2(n_369), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_321), .B(n_421), .Y(n_420) );
INVxp67_ASAP7_75t_L g428 ( .A(n_322), .Y(n_428) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_349), .Y(n_366) );
INVx1_ASAP7_75t_L g341 ( .A(n_330), .Y(n_341) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g339 ( .A(n_333), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_333), .B(n_371), .Y(n_370) );
NOR4xp25_ASAP7_75t_L g338 ( .A(n_334), .B(n_339), .C(n_340), .D(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .B1(n_353), .B2(n_354), .C1(n_356), .C2(n_360), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g440 ( .A(n_344), .Y(n_440) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_356), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_361), .A2(n_417), .B(n_419), .Y(n_416) );
NOR4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_374), .C(n_387), .D(n_402), .Y(n_362) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B1(n_366), .B2(n_367), .C(n_368), .Y(n_363) );
INVx1_ASAP7_75t_L g443 ( .A(n_364), .Y(n_443) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_371), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_380), .B2(n_381), .C1(n_384), .C2(n_386), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g409 ( .A1(n_379), .A2(n_410), .B(n_411), .C(n_422), .Y(n_409) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B1(n_394), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_407), .B1(n_440), .B2(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_437), .B(n_439), .C(n_442), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_446), .Y(n_451) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_450), .A2(n_454), .B(n_763), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B1(n_459), .B2(n_461), .Y(n_455) );
INVx2_ASAP7_75t_L g755 ( .A(n_456), .Y(n_755) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g756 ( .A(n_460), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_461), .Y(n_757) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_462), .B(n_718), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_622), .C(n_706), .Y(n_462) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_565), .C(n_587), .D(n_603), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_503), .B1(n_526), .B2(n_544), .C(n_551), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_483), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_467), .B(n_544), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g617 ( .A(n_467), .B(n_605), .C(n_618), .D(n_620), .Y(n_617) );
INVxp67_ASAP7_75t_L g734 ( .A(n_467), .Y(n_734) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g616 ( .A(n_468), .B(n_554), .Y(n_616) );
AND2x2_ASAP7_75t_L g640 ( .A(n_468), .B(n_483), .Y(n_640) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g607 ( .A(n_469), .B(n_543), .Y(n_607) );
AND2x2_ASAP7_75t_L g647 ( .A(n_469), .B(n_628), .Y(n_647) );
AND2x2_ASAP7_75t_L g664 ( .A(n_469), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_469), .B(n_484), .Y(n_688) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g542 ( .A(n_470), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g559 ( .A(n_470), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g571 ( .A(n_470), .B(n_484), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_470), .B(n_493), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_479), .B(n_480), .C(n_481), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_481), .A2(n_490), .B(n_491), .Y(n_489) );
AND2x2_ASAP7_75t_L g574 ( .A(n_483), .B(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_483), .A2(n_624), .B1(n_627), .B2(n_629), .C(n_633), .Y(n_623) );
AND2x2_ASAP7_75t_L g682 ( .A(n_483), .B(n_647), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_483), .B(n_664), .Y(n_716) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
INVx3_ASAP7_75t_L g543 ( .A(n_484), .Y(n_543) );
AND2x2_ASAP7_75t_L g591 ( .A(n_484), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g645 ( .A(n_484), .B(n_560), .Y(n_645) );
AND2x2_ASAP7_75t_L g703 ( .A(n_484), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g544 ( .A(n_493), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g560 ( .A(n_493), .Y(n_560) );
INVx1_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_493), .Y(n_621) );
AND2x2_ASAP7_75t_L g666 ( .A(n_493), .B(n_543), .Y(n_666) );
OR2x2_ASAP7_75t_L g705 ( .A(n_493), .B(n_545), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B(n_501), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_503), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_511), .Y(n_503) );
AND2x2_ASAP7_75t_L g701 ( .A(n_504), .B(n_698), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_504), .B(n_683), .Y(n_733) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g632 ( .A(n_505), .B(n_556), .Y(n_632) );
AND2x2_ASAP7_75t_L g681 ( .A(n_505), .B(n_529), .Y(n_681) );
INVx1_ASAP7_75t_L g727 ( .A(n_505), .Y(n_727) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
AND2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_556), .Y(n_582) );
INVx1_ASAP7_75t_L g599 ( .A(n_506), .Y(n_599) );
AND2x2_ASAP7_75t_L g605 ( .A(n_506), .B(n_522), .Y(n_605) );
AND2x2_ASAP7_75t_L g673 ( .A(n_511), .B(n_581), .Y(n_673) );
INVx2_ASAP7_75t_L g738 ( .A(n_511), .Y(n_738) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
AND2x2_ASAP7_75t_L g555 ( .A(n_512), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g568 ( .A(n_512), .B(n_530), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_512), .B(n_529), .Y(n_596) );
INVx1_ASAP7_75t_L g602 ( .A(n_512), .Y(n_602) );
INVx1_ASAP7_75t_L g619 ( .A(n_512), .Y(n_619) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_512), .Y(n_631) );
INVx2_ASAP7_75t_L g699 ( .A(n_512), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
INVx2_ASAP7_75t_L g556 ( .A(n_522), .Y(n_556) );
BUFx2_ASAP7_75t_L g653 ( .A(n_522), .Y(n_653) );
AND2x2_ASAP7_75t_L g698 ( .A(n_522), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_540), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_528), .B(n_635), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_528), .A2(n_697), .B(n_711), .Y(n_721) );
AND2x2_ASAP7_75t_L g746 ( .A(n_528), .B(n_632), .Y(n_746) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g668 ( .A(n_530), .Y(n_668) );
AND2x2_ASAP7_75t_L g697 ( .A(n_530), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_531), .Y(n_581) );
INVx2_ASAP7_75t_L g600 ( .A(n_531), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_531), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g554 ( .A(n_541), .Y(n_554) );
OR2x2_ASAP7_75t_L g567 ( .A(n_541), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g635 ( .A(n_541), .B(n_631), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_541), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g736 ( .A(n_541), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_541), .B(n_673), .Y(n_748) );
AND2x2_ASAP7_75t_L g627 ( .A(n_542), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g650 ( .A(n_542), .B(n_544), .Y(n_650) );
INVx2_ASAP7_75t_L g562 ( .A(n_543), .Y(n_562) );
AND2x2_ASAP7_75t_L g590 ( .A(n_543), .B(n_563), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_543), .B(n_615), .Y(n_671) );
AND2x2_ASAP7_75t_L g585 ( .A(n_544), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g732 ( .A(n_544), .Y(n_732) );
AND2x2_ASAP7_75t_L g744 ( .A(n_544), .B(n_607), .Y(n_744) );
AND2x2_ASAP7_75t_L g570 ( .A(n_545), .B(n_560), .Y(n_570) );
INVx1_ASAP7_75t_L g665 ( .A(n_545), .Y(n_665) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g563 ( .A(n_550), .B(n_564), .Y(n_563) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_554), .B(n_601), .Y(n_610) );
OR2x2_ASAP7_75t_L g742 ( .A(n_554), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g659 ( .A(n_555), .B(n_600), .Y(n_659) );
AND2x2_ASAP7_75t_L g667 ( .A(n_555), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g726 ( .A(n_555), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g750 ( .A(n_555), .B(n_597), .Y(n_750) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_556), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g737 ( .A(n_556), .B(n_600), .Y(n_737) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g589 ( .A(n_559), .B(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g751 ( .A(n_559), .Y(n_751) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
AND2x2_ASAP7_75t_L g637 ( .A(n_562), .B(n_570), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_562), .B(n_705), .Y(n_731) );
INVx2_ASAP7_75t_L g576 ( .A(n_563), .Y(n_576) );
INVx3_ASAP7_75t_L g628 ( .A(n_563), .Y(n_628) );
OR2x2_ASAP7_75t_L g656 ( .A(n_563), .B(n_657), .Y(n_656) );
AOI311xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .A3(n_571), .B(n_572), .C(n_583), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g603 ( .A1(n_566), .A2(n_604), .B(n_606), .C(n_608), .Y(n_603) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_SL g588 ( .A(n_568), .Y(n_588) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g606 ( .A(n_570), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_570), .B(n_586), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_570), .B(n_571), .Y(n_739) );
AND2x2_ASAP7_75t_L g661 ( .A(n_571), .B(n_575), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_577), .B(n_578), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g719 ( .A(n_575), .B(n_607), .Y(n_719) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_576), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g613 ( .A(n_576), .Y(n_613) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AND2x2_ASAP7_75t_L g604 ( .A(n_580), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
AND2x4_ASAP7_75t_L g711 ( .A(n_582), .B(n_680), .Y(n_711) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g662 ( .A1(n_585), .A2(n_651), .B1(n_663), .B2(n_667), .C1(n_669), .C2(n_673), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B(n_591), .C(n_594), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_588), .B(n_632), .Y(n_655) );
INVx1_ASAP7_75t_L g677 ( .A(n_590), .Y(n_677) );
INVx1_ASAP7_75t_L g611 ( .A(n_592), .Y(n_611) );
OR2x2_ASAP7_75t_L g676 ( .A(n_593), .B(n_677), .Y(n_676) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_597), .B(n_601), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_595), .B(n_613), .C(n_614), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_595), .A2(n_632), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_599), .Y(n_652) );
AND2x2_ASAP7_75t_SL g618 ( .A(n_600), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g709 ( .A(n_600), .Y(n_709) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_600), .Y(n_725) );
INVx2_ASAP7_75t_L g683 ( .A(n_601), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_605), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g657 ( .A(n_607), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B1(n_612), .B2(n_616), .C(n_617), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_611), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g745 ( .A(n_611), .Y(n_745) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g626 ( .A(n_618), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_618), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g684 ( .A(n_618), .B(n_632), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_618), .B(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g717 ( .A(n_618), .B(n_652), .Y(n_717) );
BUFx3_ASAP7_75t_L g680 ( .A(n_619), .Y(n_680) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND5xp2_ASAP7_75t_L g622 ( .A(n_623), .B(n_641), .C(n_662), .D(n_674), .E(n_689), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AOI32xp33_ASAP7_75t_L g714 ( .A1(n_626), .A2(n_653), .A3(n_669), .B1(n_715), .B2(n_717), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_628), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g638 ( .A(n_632), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B1(n_638), .B2(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_648), .B1(n_650), .B2(n_651), .C(n_654), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g713 ( .A(n_645), .B(n_664), .Y(n_713) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_650), .A2(n_711), .B1(n_729), .B2(n_734), .C(n_735), .Y(n_728) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_L g694 ( .A(n_653), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_658), .B2(n_660), .Y(n_654) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g672 ( .A(n_664), .Y(n_672) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B1(n_682), .B2(n_683), .C1(n_684), .C2(n_685), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g729 ( .A1(n_683), .A2(n_730), .B1(n_732), .B2(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_692), .B(n_695), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_700), .B(n_702), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g743 ( .A(n_698), .Y(n_743) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
A2O1A1Ixp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B(n_712), .C(n_714), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B(n_722), .C(n_747), .Y(n_718) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_719), .Y(n_723) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_728), .C(n_740), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B(n_739), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
endmodule