module fake_jpeg_29743_n_20 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_20;

wire n_13;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

INVx11_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_SL g11 ( 
.A1(n_8),
.A2(n_4),
.B1(n_3),
.B2(n_5),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_2),
.A2(n_5),
.B1(n_4),
.B2(n_7),
.Y(n_12)
);

OA22x2_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_15),
.B1(n_9),
.B2(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_19)
);

AOI322xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_13),
.A3(n_16),
.B1(n_15),
.B2(n_0),
.C1(n_6),
.C2(n_1),
.Y(n_20)
);


endmodule