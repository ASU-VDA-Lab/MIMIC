module fake_jpeg_20658_n_184 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_17),
.B1(n_21),
.B2(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_19),
.B1(n_13),
.B2(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_25),
.B1(n_22),
.B2(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_51),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_25),
.B(n_23),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_37),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_39),
.C(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_36),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_50),
.B(n_51),
.C(n_41),
.Y(n_69)
);

OR2x4_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_63),
.B(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_50),
.B1(n_63),
.B2(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_32),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_76),
.B(n_81),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_46),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_49),
.B(n_51),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_60),
.B(n_35),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_48),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_57),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_8),
.B(n_9),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_77),
.B1(n_58),
.B2(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_95),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_59),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_91),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_67),
.B1(n_55),
.B2(n_31),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_66),
.B(n_68),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_43),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_94),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_80),
.B1(n_71),
.B2(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_60),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_42),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_16),
.B1(n_18),
.B2(n_15),
.C(n_20),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_96),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_16),
.B(n_19),
.C(n_9),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_0),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_112),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_28),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_111),
.C(n_113),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_33),
.C(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_28),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_92),
.C(n_82),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.C(n_124),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_95),
.C(n_87),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_33),
.C(n_47),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_125),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_31),
.C(n_24),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_127),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_13),
.B1(n_24),
.B2(n_11),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_131),
.B(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_65),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_65),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_111),
.B1(n_115),
.B2(n_112),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_115),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_108),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_137),
.B(n_138),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_108),
.B(n_1),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_118),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_23),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_124),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_141),
.B(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_136),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_139),
.B1(n_135),
.B2(n_24),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_13),
.C(n_24),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_160),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_52),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2x1_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_52),
.Y(n_159)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_32),
.B(n_1),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_23),
.C(n_19),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_150),
.C(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_168),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_163),
.C(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_174),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_159),
.B(n_32),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_173),
.B(n_3),
.C(n_4),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_2),
.C(n_3),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_3),
.B(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

OAI321xp33_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_176),
.C(n_178),
.Y(n_179)
);

AO21x1_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_181),
.B(n_5),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_178),
.A2(n_7),
.B(n_5),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_6),
.C(n_7),
.Y(n_183)
);


endmodule