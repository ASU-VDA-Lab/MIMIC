module fake_jpeg_26181_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_1),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_2),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_7),
.C(n_12),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_17),
.B1(n_23),
.B2(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_36)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_13),
.B(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_14),
.B1(n_10),
.B2(n_19),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_37),
.B1(n_15),
.B2(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_25),
.B1(n_30),
.B2(n_10),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_26),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.C(n_38),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_38),
.B(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_43),
.C(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_8),
.B1(n_21),
.B2(n_44),
.Y(n_46)
);


endmodule