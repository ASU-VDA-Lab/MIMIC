module real_aes_943_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_0), .B(n_116), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_1), .A2(n_125), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_2), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_3), .B(n_116), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_4), .B(n_132), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_5), .B(n_132), .Y(n_491) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_7), .B(n_132), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_8), .Y(n_756) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_9), .B(n_134), .Y(n_480) );
AND2x2_ASAP7_75t_L g181 ( .A(n_10), .B(n_166), .Y(n_181) );
AND2x2_ASAP7_75t_L g189 ( .A(n_11), .B(n_110), .Y(n_189) );
INVx2_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_13), .A2(n_24), .B1(n_116), .B2(n_125), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_14), .B(n_132), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_15), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_16), .B(n_116), .Y(n_476) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_17), .A2(n_166), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_18), .B(n_151), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_19), .B(n_132), .Y(n_468) );
AO21x1_ASAP7_75t_L g486 ( .A1(n_20), .A2(n_116), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_21), .B(n_116), .Y(n_160) );
INVx1_ASAP7_75t_L g444 ( .A(n_22), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_23), .A2(n_87), .B1(n_116), .B2(n_197), .Y(n_196) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_25), .B(n_132), .Y(n_499) );
NAND2x1_ASAP7_75t_L g517 ( .A(n_26), .B(n_134), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_27), .A2(n_741), .B1(n_743), .B2(n_747), .Y(n_742) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_28), .A2(n_84), .B(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g137 ( .A(n_28), .B(n_84), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_29), .B(n_134), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_30), .B(n_132), .Y(n_479) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_31), .A2(n_110), .B(n_114), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_32), .B(n_134), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_33), .A2(n_125), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_34), .B(n_132), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_35), .A2(n_125), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g122 ( .A(n_36), .B(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g126 ( .A(n_36), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g205 ( .A(n_36), .Y(n_205) );
OR2x6_ASAP7_75t_L g442 ( .A(n_37), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_38), .B(n_116), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_39), .B(n_116), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_40), .B(n_132), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_41), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_42), .B(n_134), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_43), .B(n_116), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_44), .A2(n_125), .B(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_45), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_46), .A2(n_125), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_47), .B(n_134), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_48), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_49), .B(n_134), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_50), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g119 ( .A(n_51), .Y(n_119) );
INVx1_ASAP7_75t_L g129 ( .A(n_51), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_52), .B(n_132), .Y(n_187) );
AND2x2_ASAP7_75t_L g150 ( .A(n_53), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_54), .B(n_134), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_55), .B(n_132), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_56), .B(n_134), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_57), .A2(n_125), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_58), .B(n_116), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_59), .B(n_116), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_60), .A2(n_125), .B(n_142), .Y(n_141) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_61), .A2(n_99), .B1(n_749), .B2(n_760), .C1(n_773), .C2(n_777), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g762 ( .A1(n_61), .A2(n_102), .B1(n_103), .B2(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_61), .Y(n_763) );
AND2x2_ASAP7_75t_L g167 ( .A(n_62), .B(n_147), .Y(n_167) );
AO21x1_ASAP7_75t_L g488 ( .A1(n_63), .A2(n_125), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_64), .B(n_116), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_65), .B(n_134), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_66), .B(n_116), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_67), .B(n_134), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_68), .A2(n_92), .B1(n_125), .B2(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_69), .B(n_132), .Y(n_163) );
AND2x2_ASAP7_75t_L g510 ( .A(n_70), .B(n_147), .Y(n_510) );
INVx1_ASAP7_75t_L g121 ( .A(n_71), .Y(n_121) );
INVx1_ASAP7_75t_L g127 ( .A(n_71), .Y(n_127) );
AND2x2_ASAP7_75t_L g520 ( .A(n_72), .B(n_110), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_73), .B(n_134), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_74), .A2(n_125), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_75), .A2(n_125), .B(n_226), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_76), .A2(n_125), .B(n_130), .Y(n_124) );
AND2x2_ASAP7_75t_L g146 ( .A(n_77), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_78), .B(n_151), .Y(n_194) );
INVx1_ASAP7_75t_L g445 ( .A(n_79), .Y(n_445) );
AND2x2_ASAP7_75t_L g455 ( .A(n_80), .B(n_110), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_81), .B(n_116), .Y(n_470) );
AND2x2_ASAP7_75t_L g229 ( .A(n_82), .B(n_166), .Y(n_229) );
AND2x2_ASAP7_75t_L g487 ( .A(n_83), .B(n_136), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_85), .B(n_134), .Y(n_469) );
AND2x2_ASAP7_75t_L g502 ( .A(n_86), .B(n_110), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_88), .B(n_132), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_89), .A2(n_125), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_90), .B(n_134), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_91), .A2(n_125), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_93), .B(n_132), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_94), .B(n_132), .Y(n_460) );
BUFx2_ASAP7_75t_L g165 ( .A(n_95), .Y(n_165) );
BUFx2_ASAP7_75t_L g757 ( .A(n_96), .Y(n_757) );
BUFx2_ASAP7_75t_SL g781 ( .A(n_96), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_97), .A2(n_125), .B(n_478), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_741), .B(n_742), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_439), .B1(n_446), .B2(n_737), .Y(n_101) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_103), .A2(n_447), .B1(n_744), .B2(n_745), .Y(n_743) );
AND3x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_317), .C(n_413), .Y(n_103) );
NOR3xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_259), .C(n_286), .Y(n_104) );
OAI211xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_168), .B(n_208), .C(n_232), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_148), .Y(n_106) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_107), .A2(n_210), .B(n_214), .C(n_220), .Y(n_209) );
OR2x2_ASAP7_75t_L g332 ( .A(n_107), .B(n_269), .Y(n_332) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g299 ( .A(n_108), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_108), .B(n_270), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_108), .B(n_415), .Y(n_430) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_138), .Y(n_108) );
AND2x2_ASAP7_75t_L g216 ( .A(n_109), .B(n_149), .Y(n_216) );
INVx1_ASAP7_75t_L g236 ( .A(n_109), .Y(n_236) );
OR2x2_ASAP7_75t_L g251 ( .A(n_109), .B(n_158), .Y(n_251) );
INVx2_ASAP7_75t_L g257 ( .A(n_109), .Y(n_257) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_109), .Y(n_312) );
INVx1_ASAP7_75t_L g389 ( .A(n_109), .Y(n_389) );
INVx3_ASAP7_75t_L g139 ( .A(n_110), .Y(n_139) );
INVx4_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_111), .A2(n_183), .B(n_189), .Y(n_182) );
INVx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx4f_ASAP7_75t_L g166 ( .A(n_112), .Y(n_166) );
AND2x4_ASAP7_75t_L g136 ( .A(n_113), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_113), .B(n_137), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_124), .B(n_136), .Y(n_114) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_122), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
AND2x6_ASAP7_75t_L g134 ( .A(n_118), .B(n_127), .Y(n_134) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g132 ( .A(n_120), .B(n_129), .Y(n_132) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx5_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
AND2x2_ASAP7_75t_L g128 ( .A(n_123), .B(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_123), .Y(n_200) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
BUFx3_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
INVx2_ASAP7_75t_L g207 ( .A(n_127), .Y(n_207) );
AND2x4_ASAP7_75t_L g203 ( .A(n_128), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g199 ( .A(n_129), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_133), .B(n_135), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_134), .B(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_135), .A2(n_143), .B(n_144), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_135), .A2(n_156), .B(n_157), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_135), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_135), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_135), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_135), .A2(n_227), .B(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_135), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_135), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_135), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_135), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_135), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_135), .A2(n_507), .B(n_508), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_135), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_135), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_136), .A2(n_153), .B(n_154), .Y(n_152) );
INVx1_ASAP7_75t_SL g464 ( .A(n_136), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_136), .A2(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_136), .B(n_493), .Y(n_492) );
NOR2x1_ASAP7_75t_SL g238 ( .A(n_138), .B(n_158), .Y(n_238) );
AND2x2_ASAP7_75t_L g268 ( .A(n_138), .B(n_257), .Y(n_268) );
AO21x1_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_140), .B(n_146), .Y(n_138) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_139), .A2(n_140), .B(n_146), .Y(n_219) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_139), .A2(n_496), .B(n_502), .Y(n_495) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_139), .A2(n_504), .B(n_510), .Y(n_503) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_139), .A2(n_496), .B(n_502), .Y(n_531) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_139), .A2(n_504), .B(n_510), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_147), .Y(n_151) );
OR2x2_ASAP7_75t_L g262 ( .A(n_148), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_148), .B(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g390 ( .A(n_148), .Y(n_390) );
NAND2x1_ASAP7_75t_L g148 ( .A(n_149), .B(n_158), .Y(n_148) );
OR2x2_ASAP7_75t_SL g250 ( .A(n_149), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g254 ( .A(n_149), .Y(n_254) );
INVx4_ASAP7_75t_L g270 ( .A(n_149), .Y(n_270) );
OR2x2_ASAP7_75t_L g285 ( .A(n_149), .B(n_218), .Y(n_285) );
AND2x2_ASAP7_75t_L g324 ( .A(n_149), .B(n_238), .Y(n_324) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_149), .Y(n_336) );
OR2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_151), .Y(n_174) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_151), .A2(n_196), .B(n_202), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_151), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_151), .A2(n_457), .B(n_458), .Y(n_456) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_151), .A2(n_524), .B(n_528), .Y(n_523) );
OA21x2_ASAP7_75t_L g563 ( .A1(n_151), .A2(n_524), .B(n_528), .Y(n_563) );
AND2x2_ASAP7_75t_L g217 ( .A(n_158), .B(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g269 ( .A(n_158), .B(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g284 ( .A(n_158), .Y(n_284) );
AND2x2_ASAP7_75t_L g300 ( .A(n_158), .B(n_270), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_158), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g345 ( .A(n_158), .B(n_257), .Y(n_345) );
INVx2_ASAP7_75t_SL g415 ( .A(n_158), .Y(n_415) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_167), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_166), .Y(n_159) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp67_ASAP7_75t_L g169 ( .A(n_170), .B(n_190), .Y(n_169) );
OAI211xp5_ASAP7_75t_L g286 ( .A1(n_170), .A2(n_287), .B(n_291), .C(n_307), .Y(n_286) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g382 ( .A(n_171), .B(n_221), .Y(n_382) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_182), .Y(n_171) );
INVx2_ASAP7_75t_L g231 ( .A(n_172), .Y(n_231) );
AND2x4_ASAP7_75t_SL g242 ( .A(n_172), .B(n_222), .Y(n_242) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
AND2x2_ASAP7_75t_L g304 ( .A(n_172), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g378 ( .A(n_172), .Y(n_378) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
AND2x2_ASAP7_75t_L g323 ( .A(n_173), .B(n_182), .Y(n_323) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_181), .Y(n_173) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_174), .A2(n_514), .B(n_520), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_180), .Y(n_175) );
INVx2_ASAP7_75t_L g213 ( .A(n_182), .Y(n_213) );
AND2x2_ASAP7_75t_L g273 ( .A(n_182), .B(n_222), .Y(n_273) );
INVx2_ASAP7_75t_L g305 ( .A(n_182), .Y(n_305) );
OR2x2_ASAP7_75t_L g328 ( .A(n_182), .B(n_193), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_190), .B(n_245), .Y(n_352) );
AND2x2_ASAP7_75t_L g386 ( .A(n_190), .B(n_322), .Y(n_386) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI31xp33_ASAP7_75t_SL g307 ( .A1(n_191), .A2(n_288), .A3(n_308), .B(n_315), .Y(n_307) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_192), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx3_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
AND2x2_ASAP7_75t_L g258 ( .A(n_193), .B(n_221), .Y(n_258) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AND2x4_ASAP7_75t_L g248 ( .A(n_194), .B(n_195), .Y(n_248) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_201), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2x1p5_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx3_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g393 ( .A(n_211), .Y(n_393) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_213), .B(n_222), .Y(n_275) );
AND2x2_ASAP7_75t_L g316 ( .A(n_213), .B(n_231), .Y(n_316) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g296 ( .A(n_217), .B(n_254), .Y(n_296) );
AND2x2_ASAP7_75t_L g255 ( .A(n_218), .B(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_218), .Y(n_264) );
INVx2_ASAP7_75t_L g314 ( .A(n_218), .Y(n_314) );
AND2x2_ASAP7_75t_L g404 ( .A(n_218), .B(n_389), .Y(n_404) );
INVx3_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g410 ( .A(n_220), .Y(n_410) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_221), .B(n_280), .Y(n_349) );
AND2x2_ASAP7_75t_L g397 ( .A(n_221), .B(n_323), .Y(n_397) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g306 ( .A(n_222), .B(n_278), .Y(n_306) );
AND2x2_ASAP7_75t_L g315 ( .A(n_222), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g327 ( .A(n_222), .Y(n_327) );
BUFx2_ASAP7_75t_L g343 ( .A(n_222), .Y(n_343) );
AND2x4_ASAP7_75t_L g377 ( .A(n_222), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g422 ( .A(n_222), .B(n_323), .Y(n_422) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AOI222xp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_239), .B1(n_243), .B2(n_249), .C1(n_252), .C2(n_258), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_234), .A2(n_298), .B1(n_301), .B2(n_306), .Y(n_297) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g281 ( .A(n_235), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_SL g295 ( .A(n_235), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_235), .B(n_300), .Y(n_433) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g394 ( .A(n_236), .B(n_300), .Y(n_394) );
OR2x2_ASAP7_75t_L g371 ( .A(n_237), .B(n_253), .Y(n_371) );
OR2x2_ASAP7_75t_L g379 ( .A(n_237), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g363 ( .A(n_238), .B(n_256), .Y(n_363) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OR2x2_ASAP7_75t_L g271 ( .A(n_241), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g421 ( .A(n_241), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g372 ( .A(n_242), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_242), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g407 ( .A(n_242), .Y(n_407) );
INVxp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
INVx2_ASAP7_75t_L g392 ( .A(n_245), .Y(n_392) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g294 ( .A(n_246), .B(n_273), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_247), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g293 ( .A(n_247), .Y(n_293) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_247), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g396 ( .A(n_247), .B(n_268), .Y(n_396) );
INVx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g330 ( .A(n_248), .B(n_316), .Y(n_330) );
AND2x2_ASAP7_75t_L g373 ( .A(n_248), .B(n_305), .Y(n_373) );
AND2x4_ASAP7_75t_L g288 ( .A(n_249), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g429 ( .A(n_251), .B(n_285), .Y(n_429) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_253), .B(n_268), .Y(n_412) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_254), .B(n_268), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_254), .A2(n_295), .B(n_396), .C(n_397), .Y(n_395) );
AND2x2_ASAP7_75t_L g426 ( .A(n_254), .B(n_404), .Y(n_426) );
INVx1_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_258), .B(n_322), .Y(n_321) );
OAI21xp33_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_271), .B(n_274), .Y(n_259) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_262), .A2(n_415), .B1(n_416), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_270), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g362 ( .A(n_270), .Y(n_362) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B(n_281), .Y(n_274) );
INVx1_ASAP7_75t_L g353 ( .A(n_275), .Y(n_353) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g338 ( .A(n_293), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g375 ( .A(n_293), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_293), .B(n_323), .Y(n_411) );
INVx1_ASAP7_75t_L g431 ( .A(n_294), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_296), .A2(n_399), .B1(n_402), .B2(n_405), .C(n_408), .Y(n_398) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI321xp33_ASAP7_75t_L g419 ( .A1(n_301), .A2(n_336), .A3(n_420), .B1(n_423), .B2(n_425), .C(n_427), .Y(n_419) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g360 ( .A(n_305), .Y(n_360) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g380 ( .A(n_311), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_313), .A2(n_341), .B1(n_345), .B2(n_346), .C(n_351), .Y(n_340) );
INVxp67_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
INVx1_ASAP7_75t_L g339 ( .A(n_316), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_318), .B(n_364), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_340), .C(n_355), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_324), .B1(n_325), .B2(n_331), .C(n_333), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g438 ( .A(n_323), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_326), .B(n_329), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_327), .B(n_373), .Y(n_418) );
INVx2_ASAP7_75t_SL g350 ( .A(n_328), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_329), .A2(n_334), .B1(n_335), .B2(n_338), .Y(n_333) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_337), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_338), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g344 ( .A(n_339), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_341), .A2(n_384), .B1(n_386), .B2(n_387), .C1(n_391), .C2(n_394), .Y(n_383) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_342), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g417 ( .A(n_342), .B(n_396), .Y(n_417) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_350), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_350), .B(n_410), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_354), .Y(n_351) );
NAND2xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_361), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
NAND4xp25_ASAP7_75t_SL g364 ( .A(n_365), .B(n_383), .C(n_395), .D(n_398), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B(n_372), .C(n_374), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_371), .A2(n_375), .B1(n_379), .B2(n_381), .Y(n_374) );
INVx1_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_390), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_407), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B(n_412), .Y(n_408) );
NOR4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .C(n_432), .D(n_434), .Y(n_413) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx3_ASAP7_75t_SL g746 ( .A(n_439), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
AND2x6_ASAP7_75t_SL g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OR2x6_ASAP7_75t_SL g739 ( .A(n_441), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g748 ( .A(n_441), .B(n_442), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_441), .B(n_740), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_442), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x4_ASAP7_75t_L g447 ( .A(n_448), .B(n_646), .Y(n_447) );
NOR4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_564), .C(n_590), .D(n_630), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_481), .B(n_511), .C(n_550), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_462), .Y(n_451) );
AND2x2_ASAP7_75t_L g717 ( .A(n_452), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_453), .B(n_462), .Y(n_584) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g512 ( .A(n_454), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_454), .B(n_537), .Y(n_536) );
INVx5_ASAP7_75t_L g570 ( .A(n_454), .Y(n_570) );
NOR2x1_ASAP7_75t_SL g612 ( .A(n_454), .B(n_463), .Y(n_612) );
AND2x2_ASAP7_75t_L g668 ( .A(n_454), .B(n_474), .Y(n_668) );
OR2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_463), .B(n_474), .Y(n_540) );
AND2x2_ASAP7_75t_L g601 ( .A(n_463), .B(n_570), .Y(n_601) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_471), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_464), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_464), .A2(n_465), .B(n_471), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
AND2x2_ASAP7_75t_L g613 ( .A(n_473), .B(n_537), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_473), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g657 ( .A(n_473), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g690 ( .A(n_473), .B(n_512), .Y(n_690) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g534 ( .A(n_474), .Y(n_534) );
AND2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g602 ( .A(n_474), .Y(n_602) );
OR2x2_ASAP7_75t_L g678 ( .A(n_474), .B(n_537), .Y(n_678) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
AOI211x1_ASAP7_75t_SL g607 ( .A1(n_483), .A2(n_599), .B(n_608), .C(n_610), .Y(n_607) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_483), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_483), .B(n_650), .Y(n_697) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g547 ( .A(n_484), .Y(n_547) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
OAI21x1_ASAP7_75t_SL g485 ( .A1(n_486), .A2(n_488), .B(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g493 ( .A(n_487), .Y(n_493) );
AOI322xp5_ASAP7_75t_L g511 ( .A1(n_494), .A2(n_512), .A3(n_521), .B1(n_529), .B2(n_532), .C1(n_538), .C2(n_541), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_494), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_503), .Y(n_494) );
INVx2_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
INVxp67_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
BUFx3_ASAP7_75t_L g651 ( .A(n_495), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
INVx2_ASAP7_75t_L g560 ( .A(n_503), .Y(n_560) );
AND2x2_ASAP7_75t_L g609 ( .A(n_503), .B(n_523), .Y(n_609) );
AND2x2_ASAP7_75t_L g653 ( .A(n_503), .B(n_562), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_509), .Y(n_504) );
AND2x2_ASAP7_75t_L g538 ( .A(n_512), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_512), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_SL g732 ( .A(n_512), .B(n_567), .Y(n_732) );
INVx4_ASAP7_75t_L g537 ( .A(n_513), .Y(n_537) );
AND2x2_ASAP7_75t_L g569 ( .A(n_513), .B(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_513), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_521), .B(n_606), .Y(n_631) );
INVx1_ASAP7_75t_SL g670 ( .A(n_521), .Y(n_670) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AND2x4_ASAP7_75t_L g561 ( .A(n_522), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_522), .B(n_560), .Y(n_629) );
AND2x2_ASAP7_75t_L g681 ( .A(n_522), .B(n_531), .Y(n_681) );
OR2x2_ASAP7_75t_L g705 ( .A(n_522), .B(n_523), .Y(n_705) );
AND2x2_ASAP7_75t_L g529 ( .A(n_523), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g579 ( .A(n_523), .B(n_560), .Y(n_579) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_523), .B(n_547), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_529), .B(n_642), .Y(n_659) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g594 ( .A(n_531), .Y(n_594) );
AND2x4_ASAP7_75t_SL g634 ( .A(n_531), .B(n_548), .Y(n_634) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
OR2x2_ASAP7_75t_L g582 ( .A(n_533), .B(n_536), .Y(n_582) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g551 ( .A(n_534), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g699 ( .A(n_534), .B(n_612), .Y(n_699) );
AND2x2_ASAP7_75t_L g715 ( .A(n_534), .B(n_569), .Y(n_715) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI311xp33_ASAP7_75t_L g685 ( .A1(n_536), .A2(n_624), .A3(n_686), .B(n_688), .C(n_695), .Y(n_685) );
AND2x4_ASAP7_75t_L g552 ( .A(n_537), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g556 ( .A(n_537), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g626 ( .A(n_537), .B(n_570), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_537), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g669 ( .A(n_537), .B(n_656), .Y(n_669) );
AND2x2_ASAP7_75t_L g555 ( .A(n_539), .B(n_556), .Y(n_555) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_540), .Y(n_573) );
OR2x2_ASAP7_75t_L g662 ( .A(n_540), .B(n_626), .Y(n_662) );
INVx1_ASAP7_75t_L g718 ( .A(n_540), .Y(n_718) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g627 ( .A(n_544), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_544), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g716 ( .A(n_544), .B(n_589), .Y(n_716) );
BUFx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g559 ( .A(n_545), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g578 ( .A(n_545), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g640 ( .A(n_546), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_546), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g589 ( .A(n_547), .B(n_560), .Y(n_589) );
AND2x4_ASAP7_75t_L g642 ( .A(n_547), .B(n_549), .Y(n_642) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OAI21xp33_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_555), .B(n_557), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_551), .A2(n_637), .B1(n_641), .B2(n_643), .Y(n_636) );
AND2x2_ASAP7_75t_SL g596 ( .A(n_552), .B(n_570), .Y(n_596) );
INVx2_ASAP7_75t_L g658 ( .A(n_552), .Y(n_658) );
AND2x2_ASAP7_75t_L g672 ( .A(n_552), .B(n_668), .Y(n_672) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g568 ( .A(n_554), .Y(n_568) );
INVx1_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
INVx1_ASAP7_75t_L g572 ( .A(n_556), .Y(n_572) );
AND3x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_601), .C(n_602), .Y(n_600) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g664 ( .A(n_559), .Y(n_664) );
AND2x2_ASAP7_75t_L g592 ( .A(n_561), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g663 ( .A(n_561), .B(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_561), .A2(n_675), .B1(n_679), .B2(n_682), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_561), .B(n_709), .Y(n_713) );
BUFx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g575 ( .A(n_563), .Y(n_575) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_563), .Y(n_694) );
OAI221xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_574), .B1(n_576), .B2(n_577), .C(n_580), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_571), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g656 ( .A(n_568), .Y(n_656) );
INVx2_ASAP7_75t_SL g645 ( .A(n_569), .Y(n_645) );
AND2x2_ASAP7_75t_L g727 ( .A(n_569), .B(n_594), .Y(n_727) );
INVx4_ASAP7_75t_L g618 ( .A(n_570), .Y(n_618) );
INVx1_ASAP7_75t_L g576 ( .A(n_571), .Y(n_576) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x4_ASAP7_75t_L g687 ( .A(n_575), .B(n_642), .Y(n_687) );
INVx1_ASAP7_75t_SL g726 ( .A(n_575), .Y(n_726) );
AND2x2_ASAP7_75t_L g731 ( .A(n_575), .B(n_634), .Y(n_731) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g673 ( .A(n_579), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_583), .B(n_585), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g606 ( .A(n_587), .Y(n_606) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g603 ( .A(n_589), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g693 ( .A(n_589), .B(n_694), .Y(n_693) );
OAI211xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_595), .B(n_597), .C(n_614), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g686 ( .A(n_593), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_594), .B(n_609), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_594), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g719 ( .A(n_594), .B(n_642), .Y(n_719) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_595), .A2(n_619), .B1(n_631), .B2(n_632), .C(n_636), .Y(n_630) );
INVx3_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g701 ( .A(n_596), .B(n_602), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_603), .A3(n_605), .B1(n_607), .B2(n_611), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_601), .Y(n_691) );
INVx2_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g733 ( .A1(n_602), .A2(n_654), .B(n_734), .C(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g639 ( .A(n_604), .Y(n_639) );
OR2x2_ASAP7_75t_L g735 ( .A(n_604), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_608), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g696 ( .A(n_611), .Y(n_696) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g677 ( .A(n_612), .Y(n_677) );
OAI21xp33_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_623), .B(n_627), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
OR2x2_ASAP7_75t_L g654 ( .A(n_617), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_618), .B(n_621), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_620), .A2(n_652), .B1(n_721), .B2(n_724), .C(n_728), .Y(n_720) );
INVx2_ASAP7_75t_L g723 ( .A(n_620), .Y(n_723) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
OR2x2_ASAP7_75t_L g644 ( .A(n_624), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g711 ( .A(n_624), .B(n_669), .Y(n_711) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g709 ( .A(n_634), .Y(n_709) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_642), .B(n_672), .Y(n_729) );
INVx2_ASAP7_75t_L g736 ( .A(n_642), .Y(n_736) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_644), .A2(n_707), .B1(n_710), .B2(n_712), .C(n_714), .Y(n_706) );
AND5x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_685), .C(n_700), .D(n_720), .E(n_730), .Y(n_646) );
NOR2xp33_ASAP7_75t_SL g647 ( .A(n_648), .B(n_665), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_654), .B1(n_657), .B2(n_659), .C(n_660), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_670), .B1(n_671), .B2(n_673), .C(n_674), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_670), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
OR2x2_ASAP7_75t_L g683 ( .A(n_678), .B(n_684), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_719), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g730 ( .A1(n_716), .A2(n_731), .B(n_732), .C(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g734 ( .A(n_727), .Y(n_734) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g744 ( .A(n_738), .Y(n_744) );
CKINVDCx11_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx4_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_758), .Y(n_751) );
INVxp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_754), .B(n_757), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_SL g776 ( .A(n_755), .B(n_757), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g778 ( .A1(n_755), .A2(n_779), .B(n_782), .Y(n_778) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_R g766 ( .A(n_759), .Y(n_766) );
BUFx3_ASAP7_75t_L g771 ( .A(n_759), .Y(n_771) );
BUFx2_ASAP7_75t_L g783 ( .A(n_759), .Y(n_783) );
INVxp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B(n_767), .Y(n_761) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
NOR2xp33_ASAP7_75t_SL g767 ( .A(n_768), .B(n_772), .Y(n_767) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx9p33_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
CKINVDCx11_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
CKINVDCx8_ASAP7_75t_R g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
endmodule