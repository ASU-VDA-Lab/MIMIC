module fake_netlist_1_7608_n_753 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_753);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_753;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_216;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g82 ( .A(n_6), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_57), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_0), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_52), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_11), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_48), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_1), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_23), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_25), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_7), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_53), .Y(n_93) );
INVx1_ASAP7_75t_SL g94 ( .A(n_37), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_45), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_62), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_15), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_70), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_43), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_38), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_76), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_2), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_55), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_22), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_14), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_81), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_58), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_30), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_8), .Y(n_113) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_18), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_61), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_69), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_8), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_60), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_31), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_13), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_24), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_34), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_39), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_27), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_2), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_16), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_18), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_115), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_83), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_119), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
AND3x2_ASAP7_75t_L g136 ( .A(n_92), .B(n_0), .C(n_1), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_86), .B(n_3), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_114), .B(n_4), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_89), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_114), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_105), .Y(n_142) );
NAND2xp33_ASAP7_75t_SL g143 ( .A(n_120), .B(n_4), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_117), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_90), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_114), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_124), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_114), .Y(n_150) );
OAI21x1_ASAP7_75t_L g151 ( .A1(n_95), .A2(n_41), .B(n_78), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
NAND2xp33_ASAP7_75t_R g153 ( .A(n_84), .B(n_40), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_87), .A2(n_42), .B(n_75), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_93), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_88), .B(n_5), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_88), .B(n_6), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_100), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_131), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_100), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_94), .Y(n_163) );
NOR2xp67_ASAP7_75t_L g164 ( .A(n_96), .B(n_7), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_123), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_97), .B(n_9), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_98), .Y(n_170) );
BUFx8_ASAP7_75t_L g171 ( .A(n_106), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_101), .B(n_9), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_97), .B(n_10), .Y(n_173) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_101), .B(n_46), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_109), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_99), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_174), .A2(n_125), .B1(n_108), .B2(n_110), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_176), .B(n_130), .Y(n_179) );
AO22x2_ASAP7_75t_L g180 ( .A1(n_173), .A2(n_104), .B1(n_111), .B2(n_128), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_137), .B(n_116), .Y(n_181) );
INVx4_ASAP7_75t_SL g182 ( .A(n_173), .Y(n_182) );
INVx8_ASAP7_75t_L g183 ( .A(n_173), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_176), .B(n_130), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_173), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_144), .B(n_112), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_158), .B(n_129), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_137), .B(n_112), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_140), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_174), .B(n_121), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_145), .B(n_111), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_169), .Y(n_203) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_151), .A2(n_116), .B(n_128), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_159), .Y(n_206) );
AND2x6_ASAP7_75t_L g207 ( .A(n_167), .B(n_102), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_148), .B(n_129), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_145), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_135), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_132), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_171), .B(n_127), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_142), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_152), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_133), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_156), .B(n_103), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_156), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_135), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_171), .B(n_127), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_161), .B(n_107), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_171), .Y(n_224) );
OR2x2_ASAP7_75t_SL g225 ( .A(n_157), .B(n_99), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_161), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_166), .B(n_126), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_162), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_166), .B(n_126), .Y(n_229) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_174), .A2(n_104), .B1(n_102), .B2(n_122), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
INVx6_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_175), .B(n_122), .Y(n_233) );
AOI22xp33_ASAP7_75t_SL g234 ( .A1(n_138), .A2(n_113), .B1(n_91), .B2(n_82), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_170), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_162), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_135), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_170), .Y(n_239) );
AND2x6_ASAP7_75t_L g240 ( .A(n_157), .B(n_118), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_162), .Y(n_242) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_134), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_141), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_141), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_212), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_165), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_183), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_232), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_179), .B(n_149), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_208), .A2(n_172), .B(n_139), .C(n_103), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_224), .B(n_164), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_212), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_221), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_221), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_177), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_179), .B(n_164), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_243), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_238), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_224), .B(n_151), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_198), .A2(n_153), .B1(n_143), .B2(n_107), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_207), .B(n_118), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_238), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_194), .B(n_151), .Y(n_267) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_241), .Y(n_268) );
CKINVDCx11_ASAP7_75t_R g269 ( .A(n_213), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_207), .B(n_136), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_191), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_245), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_241), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_218), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_207), .B(n_154), .Y(n_275) );
NAND2xp33_ASAP7_75t_SL g276 ( .A(n_196), .B(n_160), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_207), .B(n_154), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_245), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_232), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_207), .B(n_154), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_182), .B(n_150), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_217), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_197), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_197), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_194), .B(n_10), .Y(n_286) );
CKINVDCx16_ASAP7_75t_R g287 ( .A(n_200), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_207), .B(n_147), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_207), .B(n_147), .Y(n_289) );
NOR2xp33_ASAP7_75t_R g290 ( .A(n_196), .B(n_49), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_230), .A2(n_147), .B1(n_141), .B2(n_150), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_187), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_194), .B(n_12), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_184), .B(n_150), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_232), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_183), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_194), .B(n_12), .Y(n_298) );
CKINVDCx11_ASAP7_75t_R g299 ( .A(n_218), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_199), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_183), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_184), .B(n_13), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_240), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_192), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_187), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_199), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_182), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_208), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_188), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_188), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_182), .B(n_14), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_189), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_192), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_246), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_182), .B(n_16), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_186), .B(n_150), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_210), .B(n_150), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_209), .B(n_17), .Y(n_319) );
NOR2xp33_ASAP7_75t_R g320 ( .A(n_215), .B(n_50), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_203), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_309), .B(n_178), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_275), .A2(n_246), .B(n_185), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_304), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g326 ( .A1(n_286), .A2(n_230), .B1(n_240), .B2(n_180), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_301), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_214), .B(n_222), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_297), .B(n_223), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_302), .B(n_240), .Y(n_331) );
CKINVDCx11_ASAP7_75t_R g332 ( .A(n_269), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_257), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_281), .A2(n_204), .B(n_228), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_286), .B(n_230), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_257), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_304), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_286), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_259), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_302), .B(n_240), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_259), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_293), .A2(n_230), .B1(n_180), .B2(n_225), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_283), .A2(n_180), .B(n_181), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_293), .B(n_223), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_260), .B(n_240), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_273), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_293), .A2(n_240), .B1(n_180), .B2(n_233), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_251), .B(n_248), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_293), .B(n_219), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_298), .A2(n_240), .B1(n_234), .B2(n_190), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_315), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_298), .A2(n_225), .B1(n_226), .B2(n_239), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_258), .B(n_219), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_298), .A2(n_226), .B1(n_217), .B2(n_239), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_268), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_271), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_271), .Y(n_363) );
AND3x1_ASAP7_75t_SL g364 ( .A(n_287), .B(n_215), .C(n_203), .Y(n_364) );
NAND2xp33_ASAP7_75t_L g365 ( .A(n_250), .B(n_235), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_297), .B(n_220), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_258), .B(n_220), .Y(n_367) );
BUFx2_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_297), .B(n_231), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_319), .A2(n_231), .B1(n_235), .B2(n_236), .Y(n_370) );
INVx5_ASAP7_75t_L g371 ( .A(n_301), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_249), .B(n_236), .Y(n_372) );
INVx3_ASAP7_75t_SL g373 ( .A(n_312), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_278), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_312), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_319), .A2(n_211), .B1(n_195), .B2(n_229), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_312), .B(n_201), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_264), .B(n_291), .C(n_267), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_287), .B1(n_274), .B2(n_264), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_360), .A2(n_319), .B1(n_316), .B2(n_312), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_368), .A2(n_274), .B1(n_320), .B2(n_290), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_332), .Y(n_384) );
AOI222xp33_ASAP7_75t_L g385 ( .A1(n_323), .A2(n_276), .B1(n_299), .B2(n_319), .C1(n_227), .C2(n_267), .Y(n_385) );
NAND2xp33_ASAP7_75t_R g386 ( .A(n_368), .B(n_261), .Y(n_386) );
NAND2xp33_ASAP7_75t_SL g387 ( .A(n_373), .B(n_316), .Y(n_387) );
AOI21xp5_ASAP7_75t_SL g388 ( .A1(n_370), .A2(n_316), .B(n_280), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_352), .A2(n_316), .B1(n_321), .B2(n_278), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_354), .B(n_284), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_336), .B(n_284), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_326), .A2(n_321), .B1(n_285), .B2(n_307), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_351), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_329), .B(n_270), .Y(n_396) );
AO31x2_ASAP7_75t_L g397 ( .A1(n_334), .A2(n_189), .A3(n_202), .B(n_205), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_371), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_371), .B(n_303), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_333), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_SL g401 ( .A1(n_333), .A2(n_307), .B(n_300), .C(n_285), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_361), .B(n_261), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_353), .B(n_303), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_329), .B(n_300), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_339), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_324), .A2(n_315), .B(n_263), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_339), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_377), .A2(n_303), .B1(n_265), .B2(n_249), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_364), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_342), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_329), .B(n_252), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_341), .A2(n_249), .B1(n_295), .B2(n_308), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_393), .B(n_336), .Y(n_415) );
OA21x2_ASAP7_75t_L g416 ( .A1(n_407), .A2(n_348), .B(n_328), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_381), .A2(n_346), .B1(n_341), .B2(n_348), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_388), .B(n_358), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_380), .A2(n_356), .B1(n_329), .B2(n_363), .C(n_375), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_400), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_389), .A2(n_263), .B(n_330), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_385), .A2(n_383), .B1(n_390), .B2(n_391), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_408), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_392), .A2(n_378), .B1(n_342), .B2(n_375), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_410), .A2(n_338), .B1(n_376), .B2(n_378), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_406), .B(n_344), .Y(n_427) );
AOI33xp33_ASAP7_75t_L g428 ( .A1(n_392), .A2(n_363), .A3(n_344), .B1(n_362), .B2(n_378), .B3(n_366), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_408), .B(n_362), .Y(n_429) );
AO22x1_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_373), .B1(n_376), .B2(n_378), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_411), .A2(n_379), .B1(n_359), .B2(n_343), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_393), .A2(n_379), .B1(n_331), .B2(n_350), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_387), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_411), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_405), .A2(n_367), .B1(n_263), .B2(n_372), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_397), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_412), .A2(n_369), .B1(n_366), .B2(n_192), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_204), .B(n_374), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_410), .A2(n_369), .B1(n_366), .B2(n_253), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_396), .B(n_366), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_397), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_394), .A2(n_374), .B(n_357), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_405), .A2(n_369), .B1(n_204), .B2(n_347), .Y(n_444) );
NAND3xp33_ASAP7_75t_SL g445 ( .A(n_422), .B(n_395), .C(n_384), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_436), .A2(n_387), .B(n_365), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_422), .B(n_395), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_424), .Y(n_448) );
NAND2xp33_ASAP7_75t_R g449 ( .A(n_433), .B(n_402), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_424), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_420), .B(n_398), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_436), .A2(n_404), .B1(n_382), .B2(n_403), .Y(n_452) );
OAI33xp33_ASAP7_75t_L g453 ( .A1(n_431), .A2(n_402), .A3(n_409), .B1(n_317), .B2(n_414), .B3(n_244), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_433), .A2(n_386), .B1(n_403), .B2(n_413), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
AOI21xp33_ASAP7_75t_SL g456 ( .A1(n_430), .A2(n_426), .B(n_417), .Y(n_456) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_431), .A2(n_345), .B(n_325), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_437), .A2(n_345), .B(n_325), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_425), .A2(n_433), .B1(n_418), .B2(n_417), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
OA332x1_ASAP7_75t_L g462 ( .A1(n_428), .A2(n_17), .A3(n_19), .B1(n_20), .B2(n_21), .B3(n_22), .C1(n_397), .C2(n_28), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_435), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_419), .A2(n_369), .B1(n_403), .B2(n_335), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_418), .A2(n_330), .B(n_322), .Y(n_465) );
OAI33xp33_ASAP7_75t_L g466 ( .A1(n_423), .A2(n_244), .A3(n_288), .B1(n_289), .B2(n_318), .B3(n_205), .Y(n_466) );
OAI22xp33_ASAP7_75t_SL g467 ( .A1(n_418), .A2(n_371), .B1(n_399), .B2(n_335), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_415), .B(n_371), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_419), .A2(n_335), .B1(n_399), .B2(n_327), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_435), .Y(n_470) );
OAI33xp33_ASAP7_75t_L g471 ( .A1(n_423), .A2(n_206), .A3(n_202), .B1(n_21), .B2(n_20), .B3(n_19), .Y(n_471) );
AND2x6_ASAP7_75t_L g472 ( .A(n_435), .B(n_399), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_429), .B(n_397), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_415), .B(n_357), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_418), .B(n_337), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_434), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_415), .B(n_371), .Y(n_477) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_421), .A2(n_206), .B(n_355), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_429), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_418), .A2(n_421), .B(n_442), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_429), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_425), .A2(n_340), .B1(n_322), .B2(n_355), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_476), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_445), .A2(n_440), .B(n_426), .C(n_438), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_455), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_475), .B(n_418), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_463), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_447), .B(n_456), .C(n_440), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_460), .A2(n_441), .B1(n_438), .B2(n_432), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_446), .A2(n_421), .B(n_442), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_473), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_473), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_479), .B(n_437), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_479), .B(n_442), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_452), .A2(n_441), .B1(n_432), .B2(n_434), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_481), .B(n_437), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_481), .B(n_443), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_464), .A2(n_444), .B1(n_427), .B2(n_434), .C(n_314), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_470), .B(n_443), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_475), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_470), .B(n_443), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_472), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_450), .B(n_443), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
AOI221x1_ASAP7_75t_L g508 ( .A1(n_465), .A2(n_427), .B1(n_340), .B2(n_315), .C(n_428), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_476), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_474), .B(n_444), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_459), .B(n_443), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_469), .A2(n_416), .B(n_327), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_451), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_461), .B(n_430), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_461), .B(n_416), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_474), .B(n_439), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_468), .B(n_327), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_458), .B(n_416), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_458), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_475), .B(n_416), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g525 ( .A1(n_462), .A2(n_314), .B1(n_305), .B2(n_347), .C1(n_282), .C2(n_337), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_457), .B(n_416), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_478), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_477), .Y(n_528) );
AO221x2_ASAP7_75t_L g529 ( .A1(n_462), .A2(n_439), .B1(n_29), .B2(n_32), .C(n_33), .Y(n_529) );
BUFx2_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
OAI221xp5_ASAP7_75t_SL g531 ( .A1(n_454), .A2(n_314), .B1(n_305), .B2(n_308), .C(n_311), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_472), .Y(n_532) );
INVx5_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
OAI33xp33_ASAP7_75t_L g534 ( .A1(n_467), .A2(n_292), .A3(n_313), .B1(n_311), .B2(n_310), .B3(n_306), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_476), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_511), .B(n_472), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_515), .B(n_472), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_489), .A2(n_482), .B(n_480), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_533), .B(n_476), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_496), .B(n_476), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_485), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_533), .Y(n_544) );
NOR4xp25_ASAP7_75t_SL g545 ( .A(n_531), .B(n_471), .C(n_453), .D(n_466), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_528), .B(n_457), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_530), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_493), .B(n_457), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_519), .B(n_478), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_498), .B(n_439), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_529), .B(n_193), .C(n_337), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_495), .B(n_439), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_498), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_484), .B(n_305), .C(n_313), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_499), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_499), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_533), .B(n_337), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_494), .B(n_439), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_506), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_495), .B(n_26), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_494), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_502), .B(n_36), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_521), .B(n_44), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_488), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_488), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_502), .B(n_47), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_504), .B(n_51), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_529), .B(n_305), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_504), .B(n_54), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_506), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_529), .B(n_337), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g577 ( .A(n_525), .B(n_306), .C(n_292), .D(n_310), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_486), .B(n_56), .Y(n_579) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_534), .B(n_256), .C(n_247), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_486), .B(n_59), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_486), .B(n_63), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_533), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_507), .Y(n_584) );
NAND4xp75_ASAP7_75t_L g585 ( .A(n_508), .B(n_64), .C(n_65), .D(n_67), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_497), .A2(n_256), .B1(n_255), .B2(n_279), .C(n_272), .Y(n_586) );
NOR3xp33_ASAP7_75t_L g587 ( .A(n_501), .B(n_247), .C(n_255), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_530), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_68), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_513), .B(n_72), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_532), .B(n_73), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_483), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_529), .B(n_74), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_490), .B(n_80), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_512), .B(n_517), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_507), .B(n_262), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_508), .B(n_193), .C(n_262), .Y(n_597) );
AO21x1_ASAP7_75t_L g598 ( .A1(n_505), .A2(n_254), .B(n_279), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_559), .B(n_503), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_599), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_559), .B(n_503), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_595), .B(n_517), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_542), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_556), .B(n_524), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g607 ( .A1(n_595), .A2(n_518), .B1(n_509), .B2(n_524), .C(n_526), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_560), .B(n_509), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_544), .A2(n_533), .B1(n_505), .B2(n_536), .Y(n_609) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_544), .A2(n_505), .B(n_535), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_556), .B(n_526), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_546), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_560), .B(n_518), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_548), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_547), .B(n_523), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_565), .B(n_510), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_549), .B(n_523), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_557), .B(n_510), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_592), .Y(n_619) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_541), .A2(n_522), .B(n_520), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_555), .B(n_522), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_563), .B(n_535), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_539), .B(n_491), .C(n_514), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_583), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_563), .B(n_527), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_575), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_577), .A2(n_527), .B1(n_296), .B2(n_250), .Y(n_627) );
OAI22xp5_ASAP7_75t_SL g628 ( .A1(n_583), .A2(n_296), .B1(n_250), .B2(n_280), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_575), .B(n_193), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_554), .A2(n_294), .B1(n_280), .B2(n_296), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_551), .B(n_272), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_551), .B(n_266), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_568), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_579), .A2(n_193), .B1(n_266), .B2(n_254), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_573), .Y(n_636) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_593), .A2(n_193), .B(n_294), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_562), .B(n_216), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_558), .B(n_296), .C(n_250), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_579), .A2(n_294), .B1(n_250), .B2(n_296), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_537), .A2(n_216), .B1(n_228), .B2(n_237), .C(n_242), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_584), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_562), .B(n_216), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_553), .B(n_228), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_594), .A2(n_237), .B1(n_250), .B2(n_296), .C(n_242), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_553), .B(n_237), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_581), .A2(n_582), .B1(n_588), .B2(n_550), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_584), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_538), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_599), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_561), .A2(n_540), .B(n_598), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_566), .B(n_570), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_566), .B(n_570), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_571), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_604), .B(n_552), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_611), .B(n_552), .Y(n_657) );
NOR2x1_ASAP7_75t_SL g658 ( .A(n_648), .B(n_540), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_611), .B(n_571), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_602), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_604), .B(n_574), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_600), .B(n_574), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_606), .B(n_590), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_602), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_619), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
AND2x4_ASAP7_75t_SL g667 ( .A(n_600), .B(n_582), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_607), .A2(n_572), .B1(n_581), .B2(n_589), .C(n_590), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_653), .A2(n_576), .B1(n_585), .B2(n_589), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_614), .B(n_545), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_614), .B(n_564), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_606), .B(n_564), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_610), .B(n_598), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_650), .B(n_597), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_626), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_605), .B(n_587), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_601), .B(n_591), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_612), .B(n_567), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_603), .B(n_596), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_608), .B(n_580), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_651), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_613), .B(n_561), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_649), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_624), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_624), .B(n_586), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_643), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_633), .B(n_585), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_634), .B(n_636), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_639), .B(n_625), .Y(n_689) );
INVxp67_ASAP7_75t_SL g690 ( .A(n_643), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_616), .B(n_618), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_615), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_629), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_617), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_670), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_666), .B(n_638), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_692), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_666), .B(n_638), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_673), .A2(n_627), .B(n_620), .C(n_623), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_691), .B(n_655), .Y(n_700) );
AND3x4_ASAP7_75t_L g701 ( .A(n_658), .B(n_627), .C(n_654), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_684), .B(n_665), .Y(n_702) );
XOR2x2_ASAP7_75t_L g703 ( .A(n_658), .B(n_609), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_691), .B(n_644), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_694), .B(n_644), .Y(n_705) );
BUFx3_ASAP7_75t_L g706 ( .A(n_686), .Y(n_706) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_690), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_665), .B(n_640), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_694), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_684), .B(n_622), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_688), .Y(n_711) );
INVxp67_ASAP7_75t_L g712 ( .A(n_687), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_667), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_689), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g715 ( .A(n_685), .B(n_652), .C(n_632), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_668), .A2(n_635), .B1(n_645), .B2(n_647), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_L g717 ( .A1(n_676), .A2(n_631), .B(n_646), .C(n_637), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_701), .A2(n_667), .B1(n_657), .B2(n_662), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_706), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_695), .A2(n_656), .B1(n_680), .B2(n_671), .C1(n_661), .C2(n_659), .Y(n_720) );
OA22x2_ASAP7_75t_L g721 ( .A1(n_701), .A2(n_669), .B1(n_659), .B2(n_663), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_703), .B(n_662), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_712), .B(n_657), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_697), .Y(n_724) );
NAND2xp33_ASAP7_75t_SL g725 ( .A(n_713), .B(n_663), .Y(n_725) );
AOI321xp33_ASAP7_75t_L g726 ( .A1(n_699), .A2(n_678), .A3(n_677), .B1(n_672), .B2(n_679), .C(n_682), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_707), .A2(n_672), .B(n_693), .Y(n_727) );
NAND2xp33_ASAP7_75t_R g728 ( .A(n_713), .B(n_674), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_712), .B(n_675), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_706), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_707), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_695), .A2(n_715), .B1(n_708), .B2(n_716), .Y(n_732) );
AND4x1_ASAP7_75t_L g733 ( .A(n_717), .B(n_674), .C(n_642), .D(n_675), .Y(n_733) );
OAI321xp33_ASAP7_75t_L g734 ( .A1(n_702), .A2(n_683), .A3(n_681), .B1(n_660), .B2(n_664), .C(n_641), .Y(n_734) );
OAI31xp33_ASAP7_75t_L g735 ( .A1(n_702), .A2(n_693), .A3(n_683), .B(n_681), .Y(n_735) );
AOI211xp5_ASAP7_75t_L g736 ( .A1(n_710), .A2(n_693), .B(n_630), .C(n_660), .Y(n_736) );
OAI322xp33_ASAP7_75t_L g737 ( .A1(n_714), .A2(n_628), .A3(n_629), .B1(n_664), .B2(n_711), .C1(n_698), .C2(n_696), .Y(n_737) );
NAND4xp25_ASAP7_75t_SL g738 ( .A(n_704), .B(n_700), .C(n_705), .D(n_709), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_710), .B(n_695), .Y(n_739) );
XNOR2xp5_ASAP7_75t_L g740 ( .A(n_733), .B(n_732), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_731), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_722), .B(n_739), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_729), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_722), .B(n_734), .C(n_737), .Y(n_744) );
AO22x2_ASAP7_75t_L g745 ( .A1(n_744), .A2(n_719), .B1(n_718), .B2(n_730), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_740), .B(n_721), .Y(n_746) );
OR4x2_ASAP7_75t_L g747 ( .A(n_740), .B(n_721), .C(n_728), .D(n_726), .Y(n_747) );
AO22x1_ASAP7_75t_L g748 ( .A1(n_747), .A2(n_742), .B1(n_741), .B2(n_743), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_746), .A2(n_725), .B1(n_738), .B2(n_735), .Y(n_749) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_745), .B1(n_728), .B2(n_720), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_749), .Y(n_751) );
AOI22xp5_ASAP7_75t_SL g752 ( .A1(n_751), .A2(n_723), .B1(n_727), .B2(n_724), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_752), .A2(n_750), .B(n_736), .Y(n_753) );
endmodule