module fake_netlist_1_2359_n_1407 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1407);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1407;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1390;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
BUFx2_ASAP7_75t_L g300 ( .A(n_48), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_143), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_196), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_9), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_169), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_125), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_41), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_6), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_134), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_257), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_213), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_222), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_78), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_179), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_232), .Y(n_314) );
INVxp67_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_120), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_31), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_299), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_256), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_220), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_117), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_267), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_156), .Y(n_324) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_178), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_199), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_227), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_202), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_180), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_51), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_123), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_20), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_25), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_204), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_60), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_25), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_30), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_211), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_144), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_253), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_41), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_298), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_255), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_264), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_176), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_168), .Y(n_349) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_250), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_53), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_186), .Y(n_352) );
INVxp33_ASAP7_75t_SL g353 ( .A(n_189), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_163), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_22), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_240), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_85), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_109), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_81), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_35), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_193), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_126), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_166), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_76), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_268), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_121), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_45), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_5), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_261), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_216), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_86), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_16), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_132), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_43), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_195), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_130), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_140), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_161), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_138), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_158), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_20), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_157), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_290), .Y(n_383) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_79), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_131), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_73), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_152), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_105), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_127), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_10), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_66), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_218), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_192), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_74), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_96), .Y(n_395) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_77), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_162), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_69), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_221), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_214), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_171), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_78), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_147), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_269), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_275), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_212), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_53), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_26), .B(n_207), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_27), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_148), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_206), .Y(n_411) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_259), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_7), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_247), .Y(n_414) );
INVxp33_ASAP7_75t_L g415 ( .A(n_243), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_28), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_42), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_5), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_63), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_6), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_39), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_85), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_14), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_27), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_159), .B(n_16), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_82), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_124), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_87), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_87), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_57), .Y(n_430) );
INVxp33_ASAP7_75t_SL g431 ( .A(n_145), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_71), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_12), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_244), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_86), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_282), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_35), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_77), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_83), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_55), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_241), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_258), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_288), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_119), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_100), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_15), .Y(n_446) );
INVxp33_ASAP7_75t_L g447 ( .A(n_106), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_238), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_362), .B(n_0), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_362), .B(n_0), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_392), .B(n_1), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_331), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_392), .B(n_313), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_300), .B(n_1), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_302), .A2(n_2), .B(n_3), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_308), .B(n_2), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_331), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_302), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_377), .B(n_3), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_335), .A2(n_4), .B1(n_7), .B2(n_8), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_314), .Y(n_461) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_314), .A2(n_4), .B(n_8), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_318), .Y(n_463) );
INVx3_ASAP7_75t_L g464 ( .A(n_313), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_331), .Y(n_465) );
INVx6_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_300), .B(n_9), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_415), .B(n_10), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_331), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_318), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_319), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_319), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_320), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_390), .B(n_11), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_390), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_317), .B(n_11), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_320), .Y(n_477) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_321), .B(n_101), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_331), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_341), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_321), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_423), .B(n_12), .Y(n_482) );
AND2x2_ASAP7_75t_SL g483 ( .A(n_448), .B(n_102), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_480), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
AO22x2_ASAP7_75t_L g486 ( .A1(n_450), .A2(n_448), .B1(n_322), .B2(n_326), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_475), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_453), .B(n_371), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_480), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_453), .B(n_316), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_480), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_453), .B(n_371), .Y(n_492) );
AND2x6_ASAP7_75t_L g493 ( .A(n_450), .B(n_322), .Y(n_493) );
AND2x6_ASAP7_75t_L g494 ( .A(n_450), .B(n_323), .Y(n_494) );
NAND3xp33_ASAP7_75t_L g495 ( .A(n_449), .B(n_433), .C(n_333), .Y(n_495) );
INVx4_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_480), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_480), .Y(n_498) );
BUFx3_ASAP7_75t_L g499 ( .A(n_466), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_466), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_479), .Y(n_501) );
AND2x4_ASAP7_75t_SL g502 ( .A(n_474), .B(n_305), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_453), .B(n_447), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_453), .B(n_402), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_480), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_453), .B(n_315), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_475), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_480), .Y(n_508) );
AND2x6_ASAP7_75t_L g509 ( .A(n_450), .B(n_323), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_454), .A2(n_394), .B1(n_417), .B2(n_396), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_450), .B(n_350), .Y(n_511) );
INVx4_ASAP7_75t_SL g512 ( .A(n_466), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_479), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_453), .B(n_402), .Y(n_514) );
BUFx4f_ASAP7_75t_L g515 ( .A(n_474), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_464), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_479), .Y(n_517) );
AND2x6_ASAP7_75t_L g518 ( .A(n_450), .B(n_326), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_458), .B(n_352), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
INVx4_ASAP7_75t_L g521 ( .A(n_451), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_479), .Y(n_522) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_465), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_458), .B(n_373), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_449), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_464), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_458), .B(n_353), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_461), .B(n_431), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_461), .B(n_365), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_451), .B(n_332), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_519), .B(n_490), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_525), .B(n_451), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_486), .A2(n_483), .B1(n_478), .B2(n_474), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_496), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_530), .B(n_451), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_529), .B(n_451), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_496), .B(n_454), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_493), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_487), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_503), .B(n_451), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_515), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_493), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_527), .B(n_451), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_493), .Y(n_545) );
INVx4_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_521), .Y(n_547) );
BUFx3_ASAP7_75t_L g548 ( .A(n_515), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_528), .B(n_454), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_487), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_530), .B(n_454), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_486), .A2(n_483), .B1(n_478), .B2(n_474), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_521), .B(n_478), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
BUFx8_ASAP7_75t_L g556 ( .A(n_493), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_506), .B(n_467), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_502), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_489), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_521), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_502), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_507), .B(n_449), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_493), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_530), .B(n_478), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_488), .B(n_467), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_486), .A2(n_483), .B1(n_478), .B2(n_474), .Y(n_570) );
INVx4_ASAP7_75t_L g571 ( .A(n_494), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_486), .A2(n_483), .B1(n_474), .B2(n_467), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_488), .B(n_467), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_497), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_516), .B(n_461), .Y(n_575) );
BUFx5_ASAP7_75t_L g576 ( .A(n_494), .Y(n_576) );
AND2x6_ASAP7_75t_L g577 ( .A(n_488), .B(n_476), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_494), .A2(n_483), .B1(n_474), .B2(n_482), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_492), .B(n_476), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_492), .B(n_474), .Y(n_580) );
BUFx4f_ASAP7_75t_L g581 ( .A(n_494), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_510), .Y(n_582) );
BUFx2_ASAP7_75t_L g583 ( .A(n_494), .Y(n_583) );
BUFx4f_ASAP7_75t_L g584 ( .A(n_494), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_509), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_492), .B(n_476), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_509), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_497), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_509), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_509), .A2(n_518), .B1(n_474), .B2(n_511), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_498), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_504), .B(n_476), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_504), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_510), .B(n_456), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_509), .Y(n_595) );
OR2x6_ASAP7_75t_L g596 ( .A(n_504), .B(n_514), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_509), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_495), .B(n_482), .Y(n_598) );
BUFx2_ASAP7_75t_L g599 ( .A(n_518), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_498), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_524), .A2(n_482), .B(n_459), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_514), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_518), .A2(n_482), .B1(n_455), .B2(n_462), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_514), .B(n_463), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_518), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_518), .A2(n_455), .B1(n_462), .B2(n_463), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_518), .Y(n_607) );
AO22x1_ASAP7_75t_L g608 ( .A1(n_516), .A2(n_459), .B1(n_456), .B2(n_325), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_505), .B(n_463), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_505), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_508), .A2(n_455), .B1(n_462), .B2(n_470), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_508), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_526), .B(n_456), .Y(n_613) );
OR2x4_ASAP7_75t_L g614 ( .A(n_526), .B(n_468), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_485), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_485), .A2(n_455), .B1(n_462), .B2(n_470), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_512), .B(n_459), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_512), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_499), .B(n_468), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_512), .Y(n_620) );
INVx4_ASAP7_75t_L g621 ( .A(n_512), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_577), .A2(n_357), .B1(n_413), .B2(n_355), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_531), .B(n_460), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_571), .B(n_332), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_573), .Y(n_625) );
INVx8_ASAP7_75t_L g626 ( .A(n_577), .Y(n_626) );
AO21x2_ASAP7_75t_L g627 ( .A1(n_570), .A2(n_471), .B(n_470), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_593), .Y(n_628) );
BUFx2_ASAP7_75t_R g629 ( .A(n_540), .Y(n_629) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_595), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_540), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_541), .A2(n_500), .B(n_499), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_551), .Y(n_633) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_596), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_573), .Y(n_635) );
NOR4xp25_ASAP7_75t_L g636 ( .A(n_566), .B(n_430), .C(n_312), .D(n_364), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_559), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_602), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_577), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_564), .B(n_460), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_577), .Y(n_642) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_577), .A2(n_446), .B1(n_462), .B2(n_455), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g644 ( .A(n_571), .B(n_460), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_552), .B(n_471), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_594), .B(n_330), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_563), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_596), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_533), .A2(n_472), .B1(n_473), .B2(n_471), .Y(n_649) );
OAI21x1_ASAP7_75t_L g650 ( .A1(n_616), .A2(n_473), .B(n_472), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_578), .A2(n_444), .B1(n_346), .B2(n_333), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_553), .A2(n_473), .B1(n_477), .B2(n_472), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_577), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_594), .B(n_330), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_552), .B(n_477), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_595), .Y(n_656) );
NOR2x1_ASAP7_75t_SL g657 ( .A(n_571), .B(n_477), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_577), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_552), .B(n_368), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_556), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_549), .B(n_368), .Y(n_661) );
INVx3_ASAP7_75t_SL g662 ( .A(n_561), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_556), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_563), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_567), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_567), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_573), .B(n_306), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_596), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_574), .Y(n_669) );
BUFx2_ASAP7_75t_L g670 ( .A(n_556), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_596), .Y(n_671) );
INVx4_ASAP7_75t_L g672 ( .A(n_560), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_578), .A2(n_481), .B1(n_381), .B2(n_424), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_574), .Y(n_674) );
BUFx8_ASAP7_75t_L g675 ( .A(n_535), .Y(n_675) );
INVx2_ASAP7_75t_SL g676 ( .A(n_614), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_536), .A2(n_481), .B1(n_337), .B2(n_344), .Y(n_677) );
AO32x2_ASAP7_75t_L g678 ( .A1(n_546), .A2(n_462), .A3(n_455), .B1(n_464), .B2(n_466), .Y(n_678) );
INVx4_ASAP7_75t_L g679 ( .A(n_560), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_537), .B(n_481), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_535), .B(n_384), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_581), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_588), .Y(n_683) );
AND2x4_ASAP7_75t_L g684 ( .A(n_535), .B(n_546), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_544), .A2(n_337), .B1(n_344), .B2(n_336), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_614), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_546), .B(n_432), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_538), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_581), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_581), .Y(n_690) );
CKINVDCx14_ASAP7_75t_R g691 ( .A(n_561), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_588), .Y(n_692) );
CKINVDCx6p67_ASAP7_75t_R g693 ( .A(n_582), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_614), .Y(n_694) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_538), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_543), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_554), .A2(n_374), .B(n_386), .C(n_307), .Y(n_697) );
INVx3_ASAP7_75t_SL g698 ( .A(n_597), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_572), .A2(n_462), .B1(n_455), .B2(n_464), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_532), .A2(n_464), .B1(n_351), .B2(n_359), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_560), .Y(n_701) );
CKINVDCx8_ASAP7_75t_R g702 ( .A(n_597), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_604), .Y(n_703) );
BUFx2_ASAP7_75t_L g704 ( .A(n_558), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_537), .Y(n_705) );
OAI222xp33_ASAP7_75t_L g706 ( .A1(n_590), .A2(n_420), .B1(n_351), .B2(n_440), .C1(n_439), .C2(n_438), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_598), .A2(n_381), .B1(n_424), .B2(n_372), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_609), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_608), .B(n_372), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_580), .A2(n_328), .B1(n_347), .B2(n_324), .Y(n_711) );
OR2x6_ASAP7_75t_L g712 ( .A(n_543), .B(n_336), .Y(n_712) );
INVx3_ASAP7_75t_L g713 ( .A(n_560), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_550), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_550), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_617), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_613), .B(n_359), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_601), .B(n_391), .Y(n_718) );
INVx3_ASAP7_75t_L g719 ( .A(n_560), .Y(n_719) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_584), .Y(n_720) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_590), .B(n_324), .Y(n_721) );
BUFx2_ASAP7_75t_L g722 ( .A(n_617), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_608), .Y(n_723) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_603), .B(n_606), .C(n_611), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_580), .A2(n_464), .B1(n_419), .B2(n_420), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_584), .Y(n_726) );
NOR2x1_ASAP7_75t_SL g727 ( .A(n_565), .B(n_327), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_568), .A2(n_419), .B1(n_421), .B2(n_418), .Y(n_728) );
INVx3_ASAP7_75t_L g729 ( .A(n_534), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_557), .A2(n_421), .B1(n_422), .B2(n_418), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_591), .Y(n_731) );
INVx5_ASAP7_75t_L g732 ( .A(n_621), .Y(n_732) );
O2A1O1Ixp5_ASAP7_75t_L g733 ( .A1(n_619), .A2(n_356), .B(n_410), .C(n_341), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_555), .A2(n_500), .B(n_501), .Y(n_734) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_584), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_555), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_605), .A2(n_328), .B1(n_354), .B2(n_347), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_534), .Y(n_738) );
BUFx3_ASAP7_75t_L g739 ( .A(n_576), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_579), .B(n_354), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_569), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_569), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_586), .B(n_363), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_545), .Y(n_744) );
INVx5_ASAP7_75t_L g745 ( .A(n_621), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_592), .A2(n_428), .B1(n_435), .B2(n_422), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_605), .A2(n_376), .B1(n_385), .B2(n_363), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_600), .Y(n_748) );
BUFx4f_ASAP7_75t_L g749 ( .A(n_545), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_600), .Y(n_750) );
INVxp67_ASAP7_75t_L g751 ( .A(n_562), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_562), .Y(n_752) );
AND3x1_ASAP7_75t_SL g753 ( .A(n_612), .B(n_435), .C(n_428), .Y(n_753) );
INVx3_ASAP7_75t_L g754 ( .A(n_534), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_612), .Y(n_755) );
OR2x6_ASAP7_75t_L g756 ( .A(n_626), .B(n_583), .Y(n_756) );
CKINVDCx6p67_ASAP7_75t_R g757 ( .A(n_662), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_676), .B(n_542), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g759 ( .A1(n_623), .A2(n_610), .B1(n_575), .B2(n_548), .C(n_542), .Y(n_759) );
NAND2x1p5_ASAP7_75t_L g760 ( .A(n_749), .B(n_583), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_637), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_626), .A2(n_548), .B1(n_610), .B2(n_599), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_646), .B(n_575), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_623), .A2(n_547), .B1(n_539), .B2(n_599), .C(n_407), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_686), .B(n_565), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_641), .A2(n_539), .B1(n_547), .B2(n_587), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_637), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_622), .A2(n_547), .B1(n_539), .B2(n_576), .Y(n_768) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_749), .B(n_587), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_633), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_628), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_638), .Y(n_772) );
INVx6_ASAP7_75t_L g773 ( .A(n_675), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_654), .B(n_576), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_691), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_631), .B(n_587), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_706), .A2(n_398), .B(n_409), .C(n_395), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_622), .A2(n_607), .B1(n_576), .B2(n_589), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_733), .B(n_724), .C(n_643), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_644), .A2(n_607), .B1(n_576), .B2(n_589), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_640), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_649), .A2(n_585), .B1(n_438), .B2(n_439), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_681), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_681), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_662), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_708), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_659), .B(n_437), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_624), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_644), .A2(n_607), .B1(n_576), .B2(n_585), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_703), .B(n_576), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_626), .A2(n_576), .B1(n_385), .B2(n_403), .Y(n_791) );
OR2x6_ASAP7_75t_L g792 ( .A(n_624), .B(n_621), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_694), .B(n_615), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_693), .B(n_615), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_684), .B(n_620), .Y(n_795) );
INVx1_ASAP7_75t_SL g796 ( .A(n_722), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g797 ( .A1(n_706), .A2(n_416), .B(n_440), .C(n_437), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_640), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_667), .Y(n_799) );
NOR2x1_ASAP7_75t_SL g800 ( .A(n_624), .B(n_620), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_651), .B(n_303), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_625), .A2(n_466), .B1(n_329), .B2(n_334), .Y(n_802) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_650), .A2(n_618), .B(n_513), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_667), .A2(n_466), .B1(n_329), .B2(n_334), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_712), .Y(n_805) );
OAI222xp33_ASAP7_75t_L g806 ( .A1(n_673), .A2(n_426), .B1(n_303), .B2(n_429), .C1(n_367), .C2(n_360), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_712), .A2(n_403), .B1(n_436), .B2(n_376), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_714), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_705), .A2(n_635), .B1(n_684), .B2(n_723), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_629), .Y(n_810) );
OR2x6_ASAP7_75t_L g811 ( .A(n_712), .B(n_660), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_634), .A2(n_466), .B1(n_338), .B2(n_339), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_716), .A2(n_441), .B1(n_436), .B2(n_412), .Y(n_813) );
INVx1_ASAP7_75t_SL g814 ( .A(n_634), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_715), .B(n_360), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_649), .A2(n_426), .B1(n_429), .B2(n_367), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_675), .Y(n_817) );
A2O1A1Ixp33_ASAP7_75t_L g818 ( .A1(n_697), .A2(n_338), .B(n_339), .C(n_327), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_736), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_647), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_741), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_725), .B(n_441), .Y(n_822) );
CKINVDCx11_ASAP7_75t_R g823 ( .A(n_702), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_704), .B(n_618), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_742), .A2(n_393), .B(n_342), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_648), .B(n_340), .Y(n_826) );
OR2x2_ASAP7_75t_L g827 ( .A(n_661), .B(n_13), .Y(n_827) );
INVx3_ASAP7_75t_L g828 ( .A(n_672), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_691), .Y(n_829) );
AND2x6_ASAP7_75t_L g830 ( .A(n_682), .B(n_340), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_647), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_716), .A2(n_304), .B1(n_310), .B2(n_309), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_652), .A2(n_343), .B1(n_345), .B2(n_342), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_687), .A2(n_345), .B1(n_349), .B2(n_343), .Y(n_834) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_663), .A2(n_445), .B1(n_414), .B2(n_358), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_668), .B(n_349), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_748), .Y(n_837) );
BUFx2_ASAP7_75t_L g838 ( .A(n_670), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_733), .B(n_425), .C(n_408), .Y(n_839) );
AND2x4_ASAP7_75t_L g840 ( .A(n_671), .B(n_358), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_687), .A2(n_427), .B1(n_434), .B2(n_361), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_639), .B(n_361), .Y(n_842) );
BUFx2_ASAP7_75t_L g843 ( .A(n_672), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_652), .A2(n_434), .B1(n_442), .B2(n_427), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_750), .Y(n_845) );
AOI221x1_ASAP7_75t_L g846 ( .A1(n_718), .A2(n_442), .B1(n_443), .B2(n_311), .C(n_401), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_643), .A2(n_443), .B1(n_369), .B2(n_375), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_642), .A2(n_370), .B1(n_379), .B2(n_378), .Y(n_848) );
OR2x6_ASAP7_75t_L g849 ( .A(n_653), .B(n_356), .Y(n_849) );
INVx4_ASAP7_75t_SL g850 ( .A(n_698), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_710), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_717), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_680), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_707), .B(n_13), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_753), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_658), .A2(n_382), .B1(n_383), .B2(n_380), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_645), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_746), .B(n_14), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g859 ( .A1(n_711), .A2(n_445), .B1(n_348), .B2(n_366), .Y(n_859) );
AND2x2_ASAP7_75t_L g860 ( .A(n_746), .B(n_15), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_657), .A2(n_301), .B1(n_388), .B2(n_387), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_725), .B(n_389), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_728), .B(n_17), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g864 ( .A1(n_721), .A2(n_655), .B1(n_743), .B2(n_740), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_685), .A2(n_399), .B(n_400), .C(n_397), .Y(n_865) );
OR2x6_ASAP7_75t_L g866 ( .A(n_688), .B(n_695), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_688), .A2(n_405), .B1(n_406), .B2(n_404), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_627), .A2(n_411), .B1(n_410), .B2(n_479), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_751), .B(n_17), .Y(n_869) );
OAI21x1_ASAP7_75t_L g870 ( .A1(n_734), .A2(n_457), .B(n_452), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_755), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_664), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_755), .Y(n_873) );
INVx4_ASAP7_75t_L g874 ( .A(n_732), .Y(n_874) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_737), .A2(n_479), .B1(n_19), .B2(n_21), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_728), .B(n_18), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_627), .A2(n_452), .B1(n_457), .B2(n_465), .Y(n_877) );
A2O1A1Ixp33_ASAP7_75t_L g878 ( .A1(n_718), .A2(n_452), .B(n_457), .C(n_520), .Y(n_878) );
INVx3_ASAP7_75t_SL g879 ( .A(n_698), .Y(n_879) );
BUFx12f_ASAP7_75t_L g880 ( .A(n_679), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_664), .Y(n_881) );
INVx4_ASAP7_75t_L g882 ( .A(n_732), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_695), .A2(n_18), .B1(n_19), .B2(n_21), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_700), .B(n_22), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_700), .B(n_23), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_696), .A2(n_452), .B1(n_457), .B2(n_465), .Y(n_886) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_730), .A2(n_452), .B1(n_457), .B2(n_501), .C(n_513), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_665), .Y(n_888) );
OAI21x1_ASAP7_75t_SL g889 ( .A1(n_727), .A2(n_23), .B(n_24), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_696), .A2(n_469), .B1(n_465), .B2(n_520), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_677), .A2(n_465), .B1(n_469), .B2(n_517), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_665), .A2(n_522), .B(n_517), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_751), .B(n_24), .Y(n_893) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_685), .A2(n_522), .B1(n_469), .B2(n_465), .C(n_523), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_752), .A2(n_469), .B1(n_465), .B2(n_523), .Y(n_895) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_677), .A2(n_26), .B1(n_28), .B2(n_29), .Y(n_896) );
INVx6_ASAP7_75t_L g897 ( .A(n_679), .Y(n_897) );
INVx6_ASAP7_75t_L g898 ( .A(n_732), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_666), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_699), .A2(n_465), .B1(n_469), .B2(n_31), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_858), .A2(n_730), .B1(n_666), .B2(n_674), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_771), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g903 ( .A1(n_852), .A2(n_636), .B1(n_699), .B2(n_747), .C(n_692), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_785), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_855), .A2(n_753), .B1(n_752), .B2(n_674), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_851), .A2(n_683), .B(n_692), .C(n_669), .Y(n_906) );
BUFx4f_ASAP7_75t_SL g907 ( .A(n_757), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_772), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_786), .Y(n_909) );
OAI33xp33_ASAP7_75t_L g910 ( .A1(n_896), .A2(n_669), .A3(n_683), .B1(n_709), .B2(n_731), .B3(n_678), .Y(n_910) );
AOI21xp5_ASAP7_75t_L g911 ( .A1(n_864), .A2(n_731), .B(n_709), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_796), .B(n_678), .Y(n_912) );
OA21x2_ASAP7_75t_L g913 ( .A1(n_779), .A2(n_803), .B(n_870), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_761), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_860), .A2(n_754), .B1(n_729), .B2(n_744), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_863), .A2(n_754), .B1(n_729), .B2(n_744), .Y(n_916) );
OR2x6_ASAP7_75t_L g917 ( .A(n_811), .B(n_744), .Y(n_917) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_787), .A2(n_738), .B1(n_632), .B2(n_701), .C(n_713), .Y(n_918) );
INVx6_ASAP7_75t_L g919 ( .A(n_880), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_853), .B(n_732), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_857), .B(n_701), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_811), .B(n_745), .Y(n_922) );
HB1xp67_ASAP7_75t_L g923 ( .A(n_866), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_799), .Y(n_924) );
AOI321xp33_ASAP7_75t_L g925 ( .A1(n_847), .A2(n_713), .A3(n_719), .B1(n_32), .B2(n_33), .C(n_34), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_796), .B(n_678), .Y(n_926) );
AOI211xp5_ASAP7_75t_L g927 ( .A1(n_859), .A2(n_719), .B(n_744), .C(n_465), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_801), .B(n_630), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_808), .B(n_630), .Y(n_929) );
OAI31xp33_ASAP7_75t_L g930 ( .A1(n_807), .A2(n_739), .A3(n_678), .B(n_32), .Y(n_930) );
INVx3_ASAP7_75t_L g931 ( .A(n_874), .Y(n_931) );
AOI211xp5_ASAP7_75t_L g932 ( .A1(n_806), .A2(n_847), .B(n_876), .C(n_875), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_869), .A2(n_739), .B1(n_689), .B2(n_735), .Y(n_933) );
OAI21xp5_ASAP7_75t_L g934 ( .A1(n_779), .A2(n_745), .B(n_656), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_819), .B(n_821), .Y(n_935) );
NAND2xp5_ASAP7_75t_SL g936 ( .A(n_805), .B(n_745), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_767), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_805), .A2(n_630), .B1(n_656), .B2(n_745), .Y(n_938) );
OAI211xp5_ASAP7_75t_L g939 ( .A1(n_861), .A2(n_465), .B(n_469), .C(n_630), .Y(n_939) );
INVx3_ASAP7_75t_L g940 ( .A(n_874), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_794), .B(n_656), .Y(n_941) );
A2O1A1Ixp33_ASAP7_75t_L g942 ( .A1(n_763), .A2(n_735), .B(n_726), .C(n_720), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_854), .A2(n_656), .B1(n_726), .B2(n_720), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_792), .A2(n_735), .B1(n_726), .B2(n_720), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_792), .A2(n_735), .B1(n_726), .B2(n_720), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_884), .A2(n_690), .B1(n_689), .B2(n_682), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_884), .A2(n_690), .B1(n_689), .B2(n_682), .Y(n_947) );
AO21x1_ASAP7_75t_L g948 ( .A1(n_900), .A2(n_29), .B(n_30), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_770), .B(n_33), .Y(n_949) );
OA21x2_ASAP7_75t_L g950 ( .A1(n_803), .A2(n_469), .B(n_523), .Y(n_950) );
INVx4_ASAP7_75t_SL g951 ( .A(n_792), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_777), .A2(n_690), .B1(n_689), .B2(n_682), .C(n_469), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g953 ( .A1(n_869), .A2(n_690), .B1(n_469), .B2(n_37), .Y(n_953) );
AND2x4_ASAP7_75t_SL g954 ( .A(n_811), .B(n_469), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_837), .B(n_34), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_788), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_956) );
OR2x2_ASAP7_75t_L g957 ( .A(n_827), .B(n_36), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_790), .A2(n_523), .B(n_104), .Y(n_958) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_867), .A2(n_759), .B1(n_841), .B2(n_834), .C(n_764), .Y(n_959) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_782), .A2(n_523), .B1(n_39), .B2(n_40), .Y(n_960) );
HB1xp67_ASAP7_75t_L g961 ( .A(n_866), .Y(n_961) );
OAI211xp5_ASAP7_75t_L g962 ( .A1(n_835), .A2(n_883), .B(n_832), .C(n_804), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_845), .Y(n_963) );
OAI22xp5_ASAP7_75t_SL g964 ( .A1(n_810), .A2(n_38), .B1(n_40), .B2(n_42), .Y(n_964) );
OAI211xp5_ASAP7_75t_L g965 ( .A1(n_865), .A2(n_43), .B(n_44), .C(n_45), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_885), .A2(n_44), .B1(n_46), .B2(n_47), .Y(n_966) );
OAI222xp33_ASAP7_75t_L g967 ( .A1(n_900), .A2(n_46), .B1(n_47), .B2(n_48), .C1(n_49), .C2(n_50), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_783), .Y(n_968) );
INVxp67_ASAP7_75t_L g969 ( .A(n_866), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_784), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_885), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_781), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_844), .B(n_52), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_849), .A2(n_52), .B1(n_54), .B2(n_55), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_817), .B(n_54), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_849), .A2(n_782), .B1(n_768), .B2(n_762), .Y(n_976) );
AO221x1_ASAP7_75t_L g977 ( .A1(n_889), .A2(n_56), .B1(n_57), .B2(n_58), .C(n_59), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_798), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_813), .B(n_56), .Y(n_979) );
AOI21xp33_ASAP7_75t_L g980 ( .A1(n_774), .A2(n_58), .B(n_59), .Y(n_980) );
HB1xp67_ASAP7_75t_L g981 ( .A(n_871), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_833), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_838), .B(n_61), .Y(n_983) );
INVx4_ASAP7_75t_L g984 ( .A(n_773), .Y(n_984) );
INVx2_ASAP7_75t_L g985 ( .A(n_820), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_893), .A2(n_62), .B1(n_63), .B2(n_64), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_833), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_987) );
O2A1O1Ixp5_ASAP7_75t_L g988 ( .A1(n_839), .A2(n_181), .B(n_295), .C(n_294), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_773), .B(n_65), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_873), .B(n_67), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_879), .B(n_67), .Y(n_991) );
AND2x4_ASAP7_75t_L g992 ( .A(n_850), .B(n_68), .Y(n_992) );
AO31x2_ASAP7_75t_L g993 ( .A1(n_846), .A2(n_891), .A3(n_816), .B(n_878), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_793), .B(n_68), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_793), .B(n_69), .Y(n_995) );
AOI222xp33_ASAP7_75t_L g996 ( .A1(n_816), .A2(n_70), .B1(n_71), .B2(n_72), .C1(n_73), .C2(n_74), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_831), .Y(n_997) );
BUFx3_ASAP7_75t_L g998 ( .A(n_775), .Y(n_998) );
NAND2xp33_ASAP7_75t_R g999 ( .A(n_843), .B(n_70), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_862), .A2(n_72), .B1(n_75), .B2(n_76), .Y(n_1000) );
OAI21x1_ASAP7_75t_L g1001 ( .A1(n_877), .A2(n_187), .B(n_293), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_797), .A2(n_75), .B1(n_79), .B2(n_80), .C(n_81), .Y(n_1002) );
OAI211xp5_ASAP7_75t_L g1003 ( .A1(n_778), .A2(n_80), .B(n_82), .C(n_83), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_814), .B(n_84), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_830), .A2(n_84), .B1(n_88), .B2(n_89), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_829), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_809), .A2(n_88), .B1(n_89), .B2(n_90), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_842), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_814), .B(n_91), .Y(n_1009) );
AOI21xp33_ASAP7_75t_L g1010 ( .A1(n_776), .A2(n_92), .B(n_93), .Y(n_1010) );
OAI21x1_ASAP7_75t_L g1011 ( .A1(n_895), .A2(n_198), .B(n_292), .Y(n_1011) );
NAND2x1_ASAP7_75t_L g1012 ( .A(n_882), .B(n_103), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_825), .A2(n_93), .B1(n_94), .B2(n_95), .C(n_96), .Y(n_1013) );
AOI21xp5_ASAP7_75t_L g1014 ( .A1(n_790), .A2(n_200), .B(n_289), .Y(n_1014) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_830), .A2(n_94), .B1(n_95), .B2(n_97), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g1016 ( .A1(n_849), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_842), .A2(n_98), .B1(n_99), .B2(n_107), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_815), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_872), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_891), .A2(n_108), .B1(n_110), .B2(n_111), .Y(n_1020) );
AOI21xp33_ASAP7_75t_L g1021 ( .A1(n_822), .A2(n_839), .B(n_868), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_815), .Y(n_1022) );
BUFx4f_ASAP7_75t_SL g1023 ( .A(n_882), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_826), .B(n_112), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1025 ( .A1(n_818), .A2(n_113), .B1(n_114), .B2(n_115), .C(n_116), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_899), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_766), .A2(n_118), .B1(n_122), .B2(n_128), .C(n_129), .Y(n_1027) );
BUFx6f_ASAP7_75t_L g1028 ( .A(n_898), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_881), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_826), .A2(n_133), .B1(n_135), .B2(n_136), .C(n_137), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_836), .Y(n_1031) );
OAI33xp33_ASAP7_75t_L g1032 ( .A1(n_1016), .A2(n_888), .A3(n_836), .B1(n_840), .B2(n_830), .B3(n_848), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_994), .B(n_840), .Y(n_1033) );
AOI222xp33_ASAP7_75t_L g1034 ( .A1(n_964), .A2(n_823), .B1(n_850), .B2(n_758), .C1(n_830), .C2(n_856), .Y(n_1034) );
OAI222xp33_ASAP7_75t_L g1035 ( .A1(n_953), .A2(n_760), .B1(n_791), .B2(n_756), .C1(n_828), .C2(n_812), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_909), .Y(n_1036) );
OAI33xp33_ASAP7_75t_L g1037 ( .A1(n_1016), .A2(n_800), .A3(n_802), .B1(n_850), .B2(n_894), .B3(n_897), .Y(n_1037) );
OAI211xp5_ASAP7_75t_SL g1038 ( .A1(n_975), .A2(n_887), .B(n_828), .C(n_886), .Y(n_1038) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_919), .Y(n_1039) );
BUFx3_ASAP7_75t_L g1040 ( .A(n_1023), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_902), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_957), .B(n_760), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_995), .B(n_758), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_951), .B(n_795), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_908), .Y(n_1045) );
INVx4_ASAP7_75t_L g1046 ( .A(n_907), .Y(n_1046) );
AOI222xp33_ASAP7_75t_L g1047 ( .A1(n_907), .A2(n_765), .B1(n_824), .B2(n_795), .C1(n_898), .C2(n_897), .Y(n_1047) );
OAI221xp5_ASAP7_75t_SL g1048 ( .A1(n_925), .A2(n_789), .B1(n_780), .B2(n_756), .C(n_890), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_963), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_950), .Y(n_1050) );
OAI31xp33_ASAP7_75t_SL g1051 ( .A1(n_976), .A2(n_765), .A3(n_769), .B(n_756), .Y(n_1051) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_959), .A2(n_769), .B1(n_892), .B2(n_142), .C(n_146), .Y(n_1052) );
AND2x6_ASAP7_75t_L g1053 ( .A(n_922), .B(n_139), .Y(n_1053) );
INVx5_ASAP7_75t_L g1054 ( .A(n_917), .Y(n_1054) );
OAI33xp33_ASAP7_75t_L g1055 ( .A1(n_956), .A2(n_141), .A3(n_149), .B1(n_150), .B2(n_151), .B3(n_153), .Y(n_1055) );
AOI322xp5_ASAP7_75t_L g1056 ( .A1(n_982), .A2(n_154), .A3(n_155), .B1(n_160), .B2(n_164), .C1(n_165), .C2(n_167), .Y(n_1056) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_967), .A2(n_170), .B1(n_172), .B2(n_173), .C(n_174), .Y(n_1057) );
AO21x2_ASAP7_75t_L g1058 ( .A1(n_934), .A2(n_175), .B(n_177), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_977), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_1059) );
AND2x6_ASAP7_75t_L g1060 ( .A(n_922), .B(n_185), .Y(n_1060) );
AOI222xp33_ASAP7_75t_L g1061 ( .A1(n_967), .A2(n_188), .B1(n_190), .B2(n_191), .C1(n_194), .C2(n_197), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_935), .Y(n_1062) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_951), .B(n_201), .Y(n_1063) );
AOI31xp33_ASAP7_75t_SL g1064 ( .A1(n_996), .A2(n_203), .A3(n_205), .B(n_208), .Y(n_1064) );
OAI221xp5_ASAP7_75t_L g1065 ( .A1(n_932), .A2(n_209), .B1(n_210), .B2(n_215), .C(n_217), .Y(n_1065) );
INVx3_ASAP7_75t_L g1066 ( .A(n_1023), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_953), .A2(n_219), .B1(n_223), .B2(n_224), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_1004), .B(n_296), .Y(n_1068) );
OA21x2_ASAP7_75t_L g1069 ( .A1(n_988), .A2(n_225), .B(n_226), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_981), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_950), .Y(n_1071) );
NOR2xp33_ASAP7_75t_R g1072 ( .A(n_999), .B(n_228), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_911), .A2(n_229), .B(n_230), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_949), .B(n_231), .Y(n_1074) );
OA21x2_ASAP7_75t_L g1075 ( .A1(n_988), .A2(n_233), .B(n_234), .Y(n_1075) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1029), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_979), .B(n_235), .Y(n_1077) );
AOI21xp33_ASAP7_75t_SL g1078 ( .A1(n_904), .A2(n_236), .B(n_237), .Y(n_1078) );
AOI32xp33_ASAP7_75t_L g1079 ( .A1(n_1005), .A2(n_239), .A3(n_242), .B1(n_245), .B2(n_246), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_983), .B(n_248), .Y(n_1080) );
NOR2xp33_ASAP7_75t_L g1081 ( .A(n_962), .B(n_249), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_948), .A2(n_252), .B1(n_254), .B2(n_260), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_1018), .A2(n_262), .B1(n_263), .B2(n_265), .Y(n_1083) );
OAI211xp5_ASAP7_75t_L g1084 ( .A1(n_1005), .A2(n_266), .B(n_270), .C(n_272), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_981), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1022), .B(n_273), .Y(n_1086) );
AND4x1_ASAP7_75t_L g1087 ( .A(n_982), .B(n_274), .C(n_276), .D(n_277), .Y(n_1087) );
OR2x2_ASAP7_75t_L g1088 ( .A(n_997), .B(n_278), .Y(n_1088) );
OAI221xp5_ASAP7_75t_L g1089 ( .A1(n_905), .A2(n_279), .B1(n_280), .B2(n_281), .C(n_283), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_989), .B(n_284), .Y(n_1090) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_919), .Y(n_1091) );
NAND3xp33_ASAP7_75t_L g1092 ( .A(n_1013), .B(n_285), .C(n_287), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_997), .B(n_955), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_923), .B(n_961), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_923), .Y(n_1095) );
INVx2_ASAP7_75t_L g1096 ( .A(n_914), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_1002), .A2(n_974), .B1(n_987), .B2(n_1010), .C(n_903), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_991), .B(n_920), .Y(n_1098) );
AOI221x1_ASAP7_75t_SL g1099 ( .A1(n_992), .A2(n_968), .B1(n_970), .B2(n_924), .C(n_980), .Y(n_1099) );
AO21x2_ASAP7_75t_L g1100 ( .A1(n_1021), .A2(n_912), .B(n_926), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_990), .Y(n_1101) );
OAI211xp5_ASAP7_75t_L g1102 ( .A1(n_1015), .A2(n_986), .B(n_987), .C(n_1000), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_960), .A2(n_1007), .B1(n_917), .B2(n_969), .Y(n_1103) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_930), .A2(n_927), .B1(n_965), .B2(n_971), .C(n_966), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1009), .Y(n_1105) );
OAI31xp33_ASAP7_75t_SL g1106 ( .A1(n_992), .A2(n_1020), .A3(n_1015), .B(n_939), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_937), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_1031), .A2(n_966), .B1(n_971), .B2(n_1000), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_941), .B(n_901), .Y(n_1109) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_917), .A2(n_969), .B1(n_961), .B2(n_1020), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_920), .B(n_954), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_972), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1113 ( .A1(n_910), .A2(n_973), .B1(n_901), .B2(n_1008), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_910), .A2(n_952), .B1(n_1017), .B2(n_951), .Y(n_1114) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_919), .Y(n_1115) );
OAI31xp33_ASAP7_75t_L g1116 ( .A1(n_1003), .A2(n_1024), .A3(n_1006), .B(n_944), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1117 ( .A1(n_906), .A2(n_942), .B(n_946), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_984), .B(n_928), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1119 ( .A1(n_921), .A2(n_918), .B1(n_915), .B2(n_916), .Y(n_1119) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_978), .B(n_985), .Y(n_1120) );
INVx3_ASAP7_75t_L g1121 ( .A(n_931), .Y(n_1121) );
AOI211xp5_ASAP7_75t_L g1122 ( .A1(n_998), .A2(n_936), .B(n_1030), .C(n_1027), .Y(n_1122) );
AOI33xp33_ASAP7_75t_L g1123 ( .A1(n_915), .A2(n_916), .A3(n_943), .B1(n_933), .B2(n_946), .B3(n_947), .Y(n_1123) );
OA222x2_ASAP7_75t_L g1124 ( .A1(n_931), .A2(n_940), .B1(n_929), .B2(n_993), .C1(n_1026), .C2(n_1019), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_940), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_984), .B(n_1028), .Y(n_1126) );
OAI21x1_ASAP7_75t_L g1127 ( .A1(n_1001), .A2(n_958), .B(n_1011), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1028), .Y(n_1128) );
OAI321xp33_ASAP7_75t_L g1129 ( .A1(n_943), .A2(n_947), .A3(n_1025), .B1(n_945), .B2(n_938), .C(n_1014), .Y(n_1129) );
OAI33xp33_ASAP7_75t_L g1130 ( .A1(n_993), .A2(n_1016), .A3(n_956), .B1(n_974), .B2(n_896), .B3(n_964), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_993), .Y(n_1131) );
INVx2_ASAP7_75t_L g1132 ( .A(n_993), .Y(n_1132) );
AOI222xp33_ASAP7_75t_L g1133 ( .A1(n_1028), .A2(n_623), .B1(n_641), .B2(n_654), .C1(n_646), .C2(n_964), .Y(n_1133) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1028), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1012), .Y(n_1135) );
NAND3xp33_ASAP7_75t_L g1136 ( .A(n_913), .B(n_835), .C(n_996), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1085), .B(n_913), .Y(n_1137) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1050), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1036), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1085), .B(n_1070), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1041), .Y(n_1141) );
BUFx2_ASAP7_75t_L g1142 ( .A(n_1095), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1076), .B(n_1131), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1063), .B(n_1054), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1045), .Y(n_1145) );
INVx4_ASAP7_75t_L g1146 ( .A(n_1054), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1131), .Y(n_1147) );
AOI31xp33_ASAP7_75t_L g1148 ( .A1(n_1034), .A2(n_1133), .A3(n_1047), .B(n_1032), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_1130), .A2(n_1032), .B1(n_1103), .B2(n_1037), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1062), .B(n_1049), .Y(n_1150) );
BUFx3_ASAP7_75t_L g1151 ( .A(n_1040), .Y(n_1151) );
INVx3_ASAP7_75t_L g1152 ( .A(n_1050), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1076), .B(n_1096), .Y(n_1153) );
AOI222xp33_ASAP7_75t_L g1154 ( .A1(n_1130), .A2(n_1102), .B1(n_1101), .B2(n_1097), .C1(n_1035), .C2(n_1103), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1094), .B(n_1095), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1120), .Y(n_1156) );
INVx3_ASAP7_75t_L g1157 ( .A(n_1071), .Y(n_1157) );
AOI33xp33_ASAP7_75t_L g1158 ( .A1(n_1105), .A2(n_1108), .A3(n_1110), .B1(n_1039), .B2(n_1091), .B3(n_1059), .Y(n_1158) );
NAND2xp5_ASAP7_75t_SL g1159 ( .A(n_1106), .B(n_1072), .Y(n_1159) );
AO21x2_ASAP7_75t_L g1160 ( .A1(n_1117), .A2(n_1110), .B(n_1071), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1112), .B(n_1033), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1096), .B(n_1107), .Y(n_1162) );
NAND4xp25_ASAP7_75t_L g1163 ( .A(n_1099), .B(n_1116), .C(n_1051), .D(n_1108), .Y(n_1163) );
NAND4xp25_ASAP7_75t_SL g1164 ( .A(n_1079), .B(n_1061), .C(n_1072), .D(n_1042), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1107), .B(n_1132), .Y(n_1165) );
AOI31xp33_ASAP7_75t_SL g1166 ( .A1(n_1122), .A2(n_1081), .A3(n_1046), .B(n_1068), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1100), .B(n_1124), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1100), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1109), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1135), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1118), .B(n_1098), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1093), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1134), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1128), .B(n_1111), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1125), .B(n_1121), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1088), .B(n_1121), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1118), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1126), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1058), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_1037), .A2(n_1104), .B1(n_1136), .B2(n_1081), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_1038), .A2(n_1052), .B1(n_1057), .B2(n_1043), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1113), .B(n_1119), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_1040), .A2(n_1066), .B1(n_1077), .B2(n_1060), .Y(n_1183) );
INVx2_ASAP7_75t_L g1184 ( .A(n_1058), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1113), .B(n_1119), .Y(n_1185) );
AND2x4_ASAP7_75t_L g1186 ( .A(n_1063), .B(n_1054), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1090), .B(n_1123), .Y(n_1187) );
CKINVDCx16_ASAP7_75t_R g1188 ( .A(n_1046), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1123), .B(n_1044), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1044), .B(n_1080), .Y(n_1190) );
NOR2xp67_ASAP7_75t_L g1191 ( .A(n_1066), .B(n_1054), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1115), .B(n_1048), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1074), .B(n_1086), .Y(n_1193) );
AOI211xp5_ASAP7_75t_L g1194 ( .A1(n_1064), .A2(n_1065), .B(n_1067), .C(n_1089), .Y(n_1194) );
AOI31xp33_ASAP7_75t_SL g1195 ( .A1(n_1082), .A2(n_1114), .A3(n_1083), .B(n_1060), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1053), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1114), .B(n_1053), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1198 ( .A(n_1082), .B(n_1092), .Y(n_1198) );
INVxp67_ASAP7_75t_SL g1199 ( .A(n_1087), .Y(n_1199) );
OAI211xp5_ASAP7_75t_SL g1200 ( .A1(n_1059), .A2(n_1056), .B(n_1083), .C(n_1084), .Y(n_1200) );
NAND3xp33_ASAP7_75t_L g1201 ( .A(n_1078), .B(n_1073), .C(n_1075), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1053), .Y(n_1202) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1069), .B(n_1075), .Y(n_1203) );
BUFx3_ASAP7_75t_L g1204 ( .A(n_1053), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1205 ( .A(n_1055), .B(n_1053), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1060), .Y(n_1206) );
NAND2xp5_ASAP7_75t_SL g1207 ( .A(n_1129), .B(n_1060), .Y(n_1207) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_1060), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1069), .B(n_1075), .Y(n_1209) );
AOI22xp33_ASAP7_75t_SL g1210 ( .A1(n_1069), .A2(n_1072), .B1(n_855), .B2(n_1060), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1127), .Y(n_1211) );
AND2x4_ASAP7_75t_L g1212 ( .A(n_1055), .B(n_1085), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1036), .Y(n_1213) );
NOR2xp67_ASAP7_75t_L g1214 ( .A(n_1046), .B(n_1066), .Y(n_1214) );
AND2x4_ASAP7_75t_SL g1215 ( .A(n_1066), .B(n_1046), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1036), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1036), .Y(n_1217) );
INVx4_ASAP7_75t_L g1218 ( .A(n_1054), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1085), .Y(n_1219) );
NAND4xp25_ASAP7_75t_L g1220 ( .A(n_1133), .B(n_460), .C(n_1099), .D(n_1034), .Y(n_1220) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_1208), .Y(n_1221) );
INVx1_ASAP7_75t_SL g1222 ( .A(n_1188), .Y(n_1222) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_1164), .A2(n_1159), .B1(n_1220), .B2(n_1163), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1219), .Y(n_1224) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1219), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1172), .B(n_1156), .Y(n_1226) );
AOI211xp5_ASAP7_75t_L g1227 ( .A1(n_1166), .A2(n_1195), .B(n_1207), .C(n_1192), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1143), .B(n_1165), .Y(n_1228) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1138), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1143), .B(n_1165), .Y(n_1230) );
INVx2_ASAP7_75t_L g1231 ( .A(n_1152), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1140), .B(n_1155), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1137), .B(n_1169), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1140), .B(n_1155), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1152), .Y(n_1235) );
NOR3xp33_ASAP7_75t_SL g1236 ( .A(n_1199), .B(n_1200), .C(n_1205), .Y(n_1236) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1137), .B(n_1169), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1177), .B(n_1150), .Y(n_1238) );
NAND5xp2_ASAP7_75t_L g1239 ( .A(n_1154), .B(n_1180), .C(n_1210), .D(n_1194), .E(n_1149), .Y(n_1239) );
OAI33xp33_ASAP7_75t_L g1240 ( .A1(n_1139), .A2(n_1141), .A3(n_1217), .B1(n_1216), .B2(n_1145), .B3(n_1213), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1157), .B(n_1153), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1157), .B(n_1153), .Y(n_1242) );
AOI21xp33_ASAP7_75t_L g1243 ( .A1(n_1148), .A2(n_1192), .B(n_1185), .Y(n_1243) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1162), .Y(n_1244) );
INVx1_ASAP7_75t_SL g1245 ( .A(n_1151), .Y(n_1245) );
OAI33xp33_ASAP7_75t_L g1246 ( .A1(n_1161), .A2(n_1171), .A3(n_1178), .B1(n_1147), .B2(n_1193), .B3(n_1176), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1142), .B(n_1147), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1142), .B(n_1160), .Y(n_1248) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_1181), .A2(n_1193), .B1(n_1183), .B2(n_1214), .C(n_1185), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1162), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1170), .Y(n_1251) );
NAND4xp25_ASAP7_75t_L g1252 ( .A(n_1167), .B(n_1158), .C(n_1189), .D(n_1187), .Y(n_1252) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_1151), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1182), .B(n_1187), .Y(n_1254) );
AND2x4_ASAP7_75t_L g1255 ( .A(n_1208), .B(n_1204), .Y(n_1255) );
NAND4xp25_ASAP7_75t_L g1256 ( .A(n_1158), .B(n_1167), .C(n_1182), .D(n_1189), .Y(n_1256) );
BUFx2_ASAP7_75t_L g1257 ( .A(n_1204), .Y(n_1257) );
AND2x4_ASAP7_75t_L g1258 ( .A(n_1196), .B(n_1206), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1160), .B(n_1168), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1160), .B(n_1173), .Y(n_1260) );
NAND3xp33_ASAP7_75t_SL g1261 ( .A(n_1198), .B(n_1190), .C(n_1202), .Y(n_1261) );
INVx3_ASAP7_75t_L g1262 ( .A(n_1144), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1173), .B(n_1170), .Y(n_1263) );
INVx3_ASAP7_75t_L g1264 ( .A(n_1144), .Y(n_1264) );
AOI221x1_ASAP7_75t_L g1265 ( .A1(n_1201), .A2(n_1179), .B1(n_1212), .B2(n_1211), .C(n_1168), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1190), .B(n_1215), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1174), .B(n_1175), .Y(n_1267) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_1212), .Y(n_1268) );
AOI32xp33_ASAP7_75t_L g1269 ( .A1(n_1215), .A2(n_1197), .A3(n_1212), .B1(n_1144), .B2(n_1186), .Y(n_1269) );
OAI31xp33_ASAP7_75t_L g1270 ( .A1(n_1197), .A2(n_1186), .A3(n_1176), .B(n_1198), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1174), .B(n_1175), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1272 ( .A(n_1146), .B(n_1218), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1186), .B(n_1179), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_1191), .Y(n_1274) );
NOR2xp33_ASAP7_75t_L g1275 ( .A(n_1146), .B(n_1218), .Y(n_1275) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1146), .B(n_1218), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1184), .B(n_1209), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1184), .B(n_1209), .Y(n_1278) );
OAI31xp33_ASAP7_75t_L g1279 ( .A1(n_1203), .A2(n_1164), .A3(n_1159), .B(n_1220), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1203), .B(n_1143), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1140), .B(n_1155), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1143), .B(n_1165), .Y(n_1282) );
AND2x2_ASAP7_75t_SL g1283 ( .A(n_1221), .B(n_1255), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1228), .B(n_1230), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1228), .B(n_1230), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1224), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1224), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1282), .B(n_1280), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1282), .B(n_1280), .Y(n_1289) );
AOI211xp5_ASAP7_75t_L g1290 ( .A1(n_1279), .A2(n_1239), .B(n_1243), .C(n_1227), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1232), .B(n_1281), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1241), .B(n_1242), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1232), .B(n_1281), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1225), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1254), .B(n_1233), .Y(n_1295) );
OAI21xp33_ASAP7_75t_L g1296 ( .A1(n_1223), .A2(n_1256), .B(n_1252), .Y(n_1296) );
NOR3xp33_ASAP7_75t_L g1297 ( .A(n_1227), .B(n_1249), .C(n_1256), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1225), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1234), .B(n_1244), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1251), .Y(n_1300) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1277), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1241), .B(n_1242), .Y(n_1302) );
INVx1_ASAP7_75t_SL g1303 ( .A(n_1245), .Y(n_1303) );
AND2x4_ASAP7_75t_SL g1304 ( .A(n_1255), .B(n_1262), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1234), .B(n_1244), .Y(n_1305) );
OR2x6_ASAP7_75t_L g1306 ( .A(n_1255), .B(n_1221), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1233), .B(n_1237), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1237), .B(n_1250), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1247), .B(n_1267), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1247), .B(n_1248), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1271), .B(n_1260), .Y(n_1311) );
AND2x4_ASAP7_75t_L g1312 ( .A(n_1258), .B(n_1273), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1251), .B(n_1260), .Y(n_1313) );
AND2x4_ASAP7_75t_L g1314 ( .A(n_1258), .B(n_1273), .Y(n_1314) );
NAND2xp5_ASAP7_75t_SL g1315 ( .A(n_1279), .B(n_1269), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_1277), .B(n_1278), .Y(n_1316) );
XOR2xp5_ASAP7_75t_L g1317 ( .A(n_1222), .B(n_1274), .Y(n_1317) );
XNOR2xp5_ASAP7_75t_L g1318 ( .A(n_1236), .B(n_1255), .Y(n_1318) );
INVx3_ASAP7_75t_L g1319 ( .A(n_1273), .Y(n_1319) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_1276), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1263), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1322 ( .A(n_1320), .B(n_1238), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1310), .B(n_1248), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1311), .B(n_1273), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1320), .B(n_1226), .Y(n_1325) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_1296), .A2(n_1246), .B1(n_1240), .B2(n_1261), .C(n_1270), .Y(n_1326) );
O2A1O1Ixp33_ASAP7_75t_L g1327 ( .A1(n_1290), .A2(n_1253), .B(n_1270), .C(n_1268), .Y(n_1327) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_1290), .A2(n_1269), .B1(n_1266), .B2(n_1257), .C(n_1276), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1316), .B(n_1263), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1313), .Y(n_1330) );
INVx1_ASAP7_75t_SL g1331 ( .A(n_1303), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1291), .Y(n_1332) );
NAND2xp5_ASAP7_75t_SL g1333 ( .A(n_1297), .B(n_1275), .Y(n_1333) );
OR2x2_ASAP7_75t_L g1334 ( .A(n_1310), .B(n_1259), .Y(n_1334) );
NAND2xp33_ASAP7_75t_SL g1335 ( .A(n_1315), .B(n_1318), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1295), .B(n_1229), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1295), .B(n_1265), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1284), .B(n_1265), .Y(n_1338) );
AOI22x1_ASAP7_75t_L g1339 ( .A1(n_1317), .A2(n_1257), .B1(n_1262), .B2(n_1264), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1291), .Y(n_1340) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1313), .Y(n_1341) );
NAND4xp25_ASAP7_75t_L g1342 ( .A(n_1296), .B(n_1272), .C(n_1259), .D(n_1262), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1300), .Y(n_1343) );
INVx1_ASAP7_75t_SL g1344 ( .A(n_1303), .Y(n_1344) );
XNOR2xp5_ASAP7_75t_L g1345 ( .A(n_1317), .B(n_1264), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1284), .B(n_1264), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1293), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_1297), .A2(n_1231), .B1(n_1235), .B2(n_1318), .Y(n_1348) );
AOI322xp5_ASAP7_75t_L g1349 ( .A1(n_1285), .A2(n_1288), .A3(n_1289), .B1(n_1307), .B2(n_1283), .C1(n_1308), .C2(n_1302), .Y(n_1349) );
XNOR2x1_ASAP7_75t_L g1350 ( .A(n_1293), .B(n_1235), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1285), .B(n_1288), .Y(n_1351) );
OAI21xp5_ASAP7_75t_SL g1352 ( .A1(n_1304), .A2(n_1319), .B(n_1312), .Y(n_1352) );
AO22x1_ASAP7_75t_L g1353 ( .A1(n_1319), .A2(n_1314), .B1(n_1312), .B2(n_1289), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_1283), .A2(n_1306), .B1(n_1304), .B2(n_1307), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1300), .Y(n_1355) );
XNOR2x2_ASAP7_75t_SL g1356 ( .A(n_1309), .B(n_1283), .Y(n_1356) );
XOR2xp5_ASAP7_75t_L g1357 ( .A(n_1309), .B(n_1299), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1308), .Y(n_1358) );
AOI221xp5_ASAP7_75t_L g1359 ( .A1(n_1321), .A2(n_1286), .B1(n_1287), .B2(n_1294), .C(n_1298), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1321), .B(n_1301), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1299), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1362 ( .A(n_1301), .B(n_1292), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1301), .B(n_1305), .Y(n_1363) );
OAI221xp5_ASAP7_75t_L g1364 ( .A1(n_1335), .A2(n_1328), .B1(n_1342), .B2(n_1326), .C(n_1333), .Y(n_1364) );
NOR2xp33_ASAP7_75t_SL g1365 ( .A(n_1339), .B(n_1354), .Y(n_1365) );
INVxp67_ASAP7_75t_L g1366 ( .A(n_1335), .Y(n_1366) );
OA22x2_ASAP7_75t_L g1367 ( .A1(n_1345), .A2(n_1352), .B1(n_1356), .B2(n_1357), .Y(n_1367) );
O2A1O1Ixp33_ASAP7_75t_L g1368 ( .A1(n_1327), .A2(n_1344), .B(n_1331), .C(n_1338), .Y(n_1368) );
XNOR2xp5_ASAP7_75t_L g1369 ( .A(n_1345), .B(n_1350), .Y(n_1369) );
NOR2xp67_ASAP7_75t_L g1370 ( .A(n_1353), .B(n_1337), .Y(n_1370) );
OAI211xp5_ASAP7_75t_L g1371 ( .A1(n_1348), .A2(n_1339), .B(n_1349), .C(n_1357), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1341), .Y(n_1372) );
INVx2_ASAP7_75t_L g1373 ( .A(n_1334), .Y(n_1373) );
AOI21xp5_ASAP7_75t_L g1374 ( .A1(n_1353), .A2(n_1350), .B(n_1322), .Y(n_1374) );
XNOR2xp5_ASAP7_75t_L g1375 ( .A(n_1347), .B(n_1332), .Y(n_1375) );
AOI21xp5_ASAP7_75t_L g1376 ( .A1(n_1325), .A2(n_1306), .B(n_1359), .Y(n_1376) );
NOR2x1_ASAP7_75t_L g1377 ( .A(n_1306), .B(n_1351), .Y(n_1377) );
AOI211x1_ASAP7_75t_L g1378 ( .A1(n_1364), .A2(n_1340), .B(n_1346), .C(n_1362), .Y(n_1378) );
O2A1O1Ixp33_ASAP7_75t_L g1379 ( .A1(n_1366), .A2(n_1323), .B(n_1358), .C(n_1330), .Y(n_1379) );
O2A1O1Ixp33_ASAP7_75t_L g1380 ( .A1(n_1368), .A2(n_1371), .B(n_1374), .C(n_1365), .Y(n_1380) );
OAI221xp5_ASAP7_75t_L g1381 ( .A1(n_1367), .A2(n_1323), .B1(n_1334), .B2(n_1341), .C(n_1330), .Y(n_1381) );
INVx1_ASAP7_75t_SL g1382 ( .A(n_1377), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1370), .B(n_1324), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_1367), .A2(n_1306), .B1(n_1304), .B2(n_1324), .Y(n_1384) );
OAI211xp5_ASAP7_75t_L g1385 ( .A1(n_1376), .A2(n_1319), .B(n_1336), .C(n_1360), .Y(n_1385) );
NAND4xp25_ASAP7_75t_SL g1386 ( .A(n_1365), .B(n_1361), .C(n_1363), .D(n_1329), .Y(n_1386) );
AOI22xp5_ASAP7_75t_L g1387 ( .A1(n_1381), .A2(n_1369), .B1(n_1375), .B2(n_1373), .Y(n_1387) );
AND2x4_ASAP7_75t_L g1388 ( .A(n_1383), .B(n_1372), .Y(n_1388) );
BUFx6f_ASAP7_75t_L g1389 ( .A(n_1383), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1379), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1391 ( .A(n_1380), .B(n_1355), .C(n_1343), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1378), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1389), .Y(n_1393) );
NOR3xp33_ASAP7_75t_L g1394 ( .A(n_1391), .B(n_1386), .C(n_1384), .Y(n_1394) );
NAND3xp33_ASAP7_75t_SL g1395 ( .A(n_1387), .B(n_1382), .C(n_1385), .Y(n_1395) );
NOR4xp25_ASAP7_75t_L g1396 ( .A(n_1392), .B(n_1363), .C(n_1355), .D(n_1343), .Y(n_1396) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1393), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1395), .Y(n_1398) );
BUFx2_ASAP7_75t_L g1399 ( .A(n_1394), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1397), .Y(n_1400) );
AND3x4_ASAP7_75t_L g1401 ( .A(n_1397), .B(n_1396), .C(n_1388), .Y(n_1401) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1398), .A2(n_1390), .B1(n_1388), .B2(n_1306), .Y(n_1402) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1400), .Y(n_1403) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_1402), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1401), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g1406 ( .A(n_1403), .Y(n_1406) );
AOI22xp33_ASAP7_75t_SL g1407 ( .A1(n_1406), .A2(n_1399), .B1(n_1404), .B2(n_1405), .Y(n_1407) );
endmodule