module fake_jpeg_28799_n_239 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_2),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_2),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_35),
.Y(n_73)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_22),
.Y(n_48)
);

CKINVDCx9p33_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_3),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_30),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_52),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_28),
.B1(n_26),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_53),
.A2(n_59),
.B1(n_62),
.B2(n_65),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_17),
.B(n_33),
.C(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_35),
.B1(n_27),
.B2(n_29),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_33),
.B1(n_22),
.B2(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_70),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_3),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_34),
.B(n_5),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_4),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_16),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_24),
.B1(n_32),
.B2(n_19),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_102),
.B(n_109),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_92),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_74),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_24),
.A3(n_34),
.B1(n_7),
.B2(n_9),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_95),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_55),
.B(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_107),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_15),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_58),
.A2(n_42),
.B(n_36),
.C(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_15),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_74),
.C(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_5),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_51),
.B1(n_81),
.B2(n_54),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_125),
.B1(n_130),
.B2(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_121),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_98),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_80),
.B(n_70),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_124),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_80),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_42),
.B1(n_36),
.B2(n_72),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_43),
.B1(n_42),
.B2(n_57),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_84),
.B1(n_100),
.B2(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_43),
.B1(n_69),
.B2(n_34),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_69),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_135),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_69),
.B1(n_66),
.B2(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_69),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_66),
.B1(n_7),
.B2(n_9),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_84),
.B1(n_104),
.B2(n_91),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_121),
.B(n_109),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_120),
.B(n_105),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_109),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_130),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_138),
.B(n_89),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_146),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_116),
.B1(n_127),
.B2(n_131),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_161),
.C(n_96),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_87),
.B1(n_82),
.B2(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_154),
.B1(n_162),
.B2(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_158),
.Y(n_170)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_106),
.B1(n_105),
.B2(n_96),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_129),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_111),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_111),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_168),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_147),
.B(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_164),
.B1(n_178),
.B2(n_160),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_133),
.B1(n_131),
.B2(n_114),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_114),
.B1(n_125),
.B2(n_106),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_139),
.B(n_154),
.Y(n_182)
);

XOR2x2_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_119),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_156),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_111),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_189),
.B(n_173),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_157),
.C(n_148),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_197),
.C(n_167),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_149),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_196),
.B1(n_156),
.B2(n_179),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_165),
.B(n_140),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_205),
.B(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_209),
.C(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_203),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_183),
.A2(n_165),
.B1(n_181),
.B2(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_160),
.B1(n_176),
.B2(n_175),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_186),
.Y(n_207)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_175),
.C(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_211),
.Y(n_224)
);

AOI31xp67_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_185),
.A3(n_195),
.B(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_209),
.C(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_212),
.B(n_215),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_186),
.C(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_204),
.B1(n_205),
.B2(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_194),
.C(n_159),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_221),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_222),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_214),
.C(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_66),
.C(n_11),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_208),
.A3(n_153),
.B1(n_152),
.B2(n_144),
.C1(n_13),
.C2(n_7),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_10),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_232),
.C(n_226),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_227),
.A2(n_220),
.B1(n_11),
.B2(n_12),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_233),
.B1(n_228),
.B2(n_13),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_225),
.C(n_10),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_236),
.Y(n_239)
);


endmodule