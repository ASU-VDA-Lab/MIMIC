module real_jpeg_31455_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_542, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_542;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_0),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_0),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_1),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_1),
.A2(n_137),
.B1(n_178),
.B2(n_183),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_1),
.A2(n_69),
.B1(n_137),
.B2(n_534),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_2),
.A2(n_115),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_2),
.A2(n_115),
.B1(n_395),
.B2(n_399),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_2),
.A2(n_115),
.B1(n_439),
.B2(n_443),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_3),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_3),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_244),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_3),
.A2(n_244),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_6),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_6),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_7),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_7),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_7),
.A2(n_74),
.B1(n_107),
.B2(n_110),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_7),
.A2(n_74),
.B1(n_285),
.B2(n_287),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_7),
.A2(n_74),
.B1(n_375),
.B2(n_379),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_8),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_8),
.A2(n_63),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_8),
.A2(n_63),
.B1(n_343),
.B2(n_348),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_8),
.A2(n_63),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_9),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_11),
.Y(n_192)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

AO22x1_ASAP7_75t_L g522 ( 
.A1(n_12),
.A2(n_224),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_14),
.A2(n_149),
.B1(n_209),
.B2(n_213),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g231 ( 
.A1(n_15),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_154),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_16),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_16),
.B(n_122),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_16),
.A2(n_302),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

OAI21xp33_ASAP7_75t_L g480 ( 
.A1(n_16),
.A2(n_227),
.B(n_427),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_505),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_332),
.B(n_501),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_273),
.B(n_306),
.Y(n_20)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_21),
.Y(n_503)
);

XNOR2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_173),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_22),
.B(n_174),
.C(n_509),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.C(n_123),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_23),
.A2(n_24),
.B1(n_79),
.B2(n_80),
.Y(n_276)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_58),
.B(n_66),
.Y(n_24)
);

OAI22x1_ASAP7_75t_L g255 ( 
.A1(n_25),
.A2(n_256),
.B1(n_257),
.B2(n_265),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_25),
.A2(n_66),
.B(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22x1_ASAP7_75t_L g291 ( 
.A1(n_26),
.A2(n_292),
.B1(n_296),
.B2(n_297),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_26),
.B(n_68),
.Y(n_330)
);

AOI22x1_ASAP7_75t_L g532 ( 
.A1(n_26),
.A2(n_67),
.B1(n_258),
.B2(n_533),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

AOI22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_31),
.Y(n_369)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_34),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_40),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_41),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_51),
.B2(n_55),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_46),
.Y(n_405)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_56),
.Y(n_537)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_57),
.Y(n_264)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_58),
.Y(n_296)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_60),
.Y(n_293)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_62),
.Y(n_295)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_68),
.Y(n_256)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_72),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_73),
.Y(n_409)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_78),
.Y(n_365)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_113),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_106),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_82),
.A2(n_114),
.B1(n_122),
.B2(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_82),
.A2(n_299),
.B(n_304),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_82),
.B(n_267),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_96),
.Y(n_301)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_106),
.B(n_122),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g272 ( 
.A(n_121),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_123),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_152),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_125),
.B(n_152),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_132),
.B1(n_141),
.B2(n_144),
.Y(n_125)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_126),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_126),
.B(n_144),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_126),
.B(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_126),
.A2(n_437),
.B1(n_446),
.B2(n_448),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_126),
.A2(n_231),
.B(n_517),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_127),
.Y(n_447)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g429 ( 
.A(n_128),
.Y(n_429)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_131),
.Y(n_426)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_131),
.Y(n_488)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_133),
.A2(n_227),
.B1(n_318),
.B2(n_324),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_140),
.Y(n_320)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_140),
.Y(n_442)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_143),
.Y(n_517)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AO32x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_157),
.A3(n_160),
.B1(n_164),
.B2(n_165),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_156),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_164),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2x1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_237),
.Y(n_173)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_218),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_176),
.B(n_218),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_187),
.B1(n_208),
.B2(n_216),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_187),
.B1(n_216),
.B2(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_184),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_186),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_187),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_187),
.B(n_208),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_200),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_197),
.Y(n_459)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_205),
.B2(n_207),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_202),
.Y(n_290)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_202),
.Y(n_350)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_207),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_214),
.B(n_302),
.Y(n_461)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_216),
.A2(n_341),
.B1(n_342),
.B2(n_394),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_216),
.A2(n_394),
.B(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_216),
.B(n_302),
.Y(n_477)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_217),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_217),
.B(n_284),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_217),
.B(n_522),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_228),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_249),
.B(n_253),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_224),
.B(n_225),
.Y(n_219)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_220),
.Y(n_421)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_227),
.A2(n_420),
.B(n_427),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

BUFx4f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_235),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_237),
.Y(n_509)
);

XOR2x1_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_254),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g511 ( 
.A(n_238),
.B(n_266),
.C(n_512),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_248),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_247),
.Y(n_357)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_247),
.Y(n_361)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_252),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_266),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_255),
.Y(n_512)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_265),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_265),
.A2(n_329),
.B(n_330),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_265),
.B(n_302),
.Y(n_430)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_274),
.B(n_503),
.C(n_504),
.Y(n_502)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_280),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_291),
.C(n_298),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_281),
.B(n_291),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_283),
.B(n_284),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_283),
.B(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_302),
.B(n_303),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_355),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_359),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_SL g474 ( 
.A1(n_302),
.A2(n_344),
.B(n_461),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_302),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_305),
.B(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_307),
.B(n_309),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_310),
.B(n_383),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_328),
.B(n_331),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_327),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_327),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_318),
.A2(n_371),
.B(n_373),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_325),
.Y(n_485)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_328),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_385),
.B(n_499),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_382),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_336),
.B(n_500),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_339),
.C(n_352),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_337),
.B(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_339),
.A2(n_340),
.B1(n_352),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B(n_351),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_347),
.Y(n_471)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_351),
.B(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_370),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_370),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_357),
.B1(n_358),
.B2(n_362),
.Y(n_353)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_SL g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_373),
.A2(n_438),
.B(n_447),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_410),
.B(n_498),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_387),
.B(n_390),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.C(n_401),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_391),
.A2(n_413),
.B1(n_414),
.B2(n_416),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_401),
.Y(n_414)
);

BUFx4f_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

OAI321xp33_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_434),
.A3(n_491),
.B1(n_495),
.B2(n_496),
.C(n_542),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_415),
.B(n_417),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_417),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_430),
.C(n_431),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_494),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_430),
.B(n_432),
.Y(n_494)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_475),
.B(n_490),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_449),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_436),
.B(n_449),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_472),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_472),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_460),
.B1(n_462),
.B2(n_467),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_456),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_468),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_479),
.B(n_489),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_477),
.B(n_478),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_486),
.Y(n_481)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_493),
.Y(n_495)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_538),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_510),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_510),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_527),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_518),
.B1(n_519),
.B2(n_526),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_516),
.Y(n_526)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_525),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_532),
.Y(n_529)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);


endmodule