module real_jpeg_5295_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_0),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_0),
.A2(n_66),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_0),
.A2(n_66),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_0),
.A2(n_66),
.B1(n_290),
.B2(n_389),
.Y(n_388)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g448 ( 
.A(n_1),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_3),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_102),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_102),
.B1(n_192),
.B2(n_195),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_4),
.A2(n_50),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g359 ( 
.A1(n_4),
.A2(n_50),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_4),
.A2(n_50),
.B1(n_164),
.B2(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_5),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_5),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_128),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_128),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_5),
.A2(n_128),
.B1(n_304),
.B2(n_312),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_134),
.B1(n_136),
.B2(n_140),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_6),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_6),
.A2(n_140),
.B1(n_164),
.B2(n_167),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_140),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_7),
.Y(n_406)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_8),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_9),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_9),
.A2(n_207),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_9),
.A2(n_207),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_9),
.A2(n_207),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_14),
.A2(n_248),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_14),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_14),
.A2(n_250),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_14),
.A2(n_250),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_14),
.A2(n_250),
.B1(n_352),
.B2(n_426),
.Y(n_425)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_16),
.A2(n_237),
.B1(n_238),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_16),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_16),
.B(n_275),
.C(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_16),
.B(n_115),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_16),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_16),
.B(n_168),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_16),
.B(n_347),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_17),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_18),
.A2(n_120),
.B1(n_238),
.B2(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_18),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_18),
.A2(n_296),
.B1(n_311),
.B2(n_316),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_18),
.A2(n_46),
.B1(n_296),
.B2(n_354),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_18),
.A2(n_32),
.B1(n_33),
.B2(n_296),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_496),
.B(n_498),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_211),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_210),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_157),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_24),
.B(n_157),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_141),
.B2(n_142),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_67),
.C(n_103),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_27),
.A2(n_143),
.B1(n_144),
.B2(n_156),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_27),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_27),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_48),
.B1(n_57),
.B2(n_59),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_28),
.A2(n_57),
.B1(n_59),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_28),
.A2(n_247),
.B(n_252),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_28),
.A2(n_39),
.B1(n_247),
.B2(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_29),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_29),
.A2(n_420),
.B(n_422),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_30)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_33),
.Y(n_154)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_34),
.Y(n_403)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_39),
.B(n_264),
.Y(n_386)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_41),
.Y(n_344)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_43),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_44),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_44),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_44),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_44),
.Y(n_243)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_49),
.B(n_58),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_51),
.B(n_264),
.Y(n_408)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_57),
.A2(n_205),
.B(n_451),
.Y(n_466)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_58),
.B(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g421 ( 
.A(n_62),
.Y(n_421)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_67),
.A2(n_68),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_67),
.A2(n_68),
.B1(n_103),
.B2(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_87),
.B(n_96),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_69),
.A2(n_263),
.B(n_265),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_69),
.A2(n_87),
.B1(n_295),
.B2(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_69),
.A2(n_265),
.B(n_338),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_69),
.A2(n_87),
.B1(n_428),
.B2(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_70),
.A2(n_163),
.B1(n_168),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_70),
.A2(n_168),
.B1(n_198),
.B2(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_70),
.B(n_266),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_87),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_74),
.Y(n_269)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_75),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_75),
.Y(n_431)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_76),
.Y(n_238)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_76),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx5_ASAP7_75t_SL g368 ( 
.A(n_84),
.Y(n_368)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_85),
.Y(n_267)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_87),
.A2(n_295),
.B(n_297),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_87),
.A2(n_297),
.B(n_428),
.Y(n_427)
);

AOI22x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_90),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_91),
.Y(n_318)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_92),
.Y(n_277)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_125),
.B1(n_132),
.B2(n_133),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_132),
.B1(n_133),
.B2(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_105),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_105),
.A2(n_132),
.B1(n_173),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_105),
.A2(n_132),
.B1(n_382),
.B2(n_425),
.Y(n_424)
);

OR2x2_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_115),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_106)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_107),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_114),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_114),
.Y(n_426)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_115),
.A2(n_126),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_115),
.A2(n_171),
.B1(n_384),
.B2(n_453),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_118),
.Y(n_369)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g370 ( 
.A(n_120),
.B(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_132),
.B(n_351),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_132),
.A2(n_382),
.B(n_383),
.Y(n_381)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_135),
.Y(n_353)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_139),
.Y(n_349)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_179),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_158),
.B(n_161),
.CI(n_179),
.CON(n_213),
.SN(n_213)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_170),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_168),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_171),
.A2(n_343),
.B(n_350),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_171),
.B(n_384),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_171),
.A2(n_350),
.B(n_469),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_174),
.B(n_405),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B(n_203),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_197),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_203),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_181),
.A2(n_197),
.B1(n_219),
.B2(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_189),
.B(n_191),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_191),
.B1(n_226),
.B2(n_232),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_182),
.A2(n_280),
.B(n_286),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_182),
.A2(n_264),
.B(n_286),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_182),
.A2(n_189),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_183),
.B(n_288),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_183),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_183),
.A2(n_359),
.B1(n_388),
.B2(n_391),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_183),
.A2(n_413),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_185),
.Y(n_327)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_185),
.Y(n_392)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_186),
.Y(n_304)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_189),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_189),
.A2(n_310),
.B(n_319),
.Y(n_309)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_192),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_197),
.Y(n_440)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_202),
.Y(n_340)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_253),
.B(n_495),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_213),
.B(n_214),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_213),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.C(n_223),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_220),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_223),
.B(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_239),
.C(n_246),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_224),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_225),
.B(n_235),
.Y(n_463)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_226),
.Y(n_446)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_227),
.Y(n_360)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_236),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_239),
.B(n_246),
.Y(n_438)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_240),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_245),
.Y(n_355)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_245),
.Y(n_367)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_252),
.Y(n_422)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI311xp33_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_434),
.A3(n_471),
.B1(n_489),
.C1(n_490),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_395),
.B(n_433),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_373),
.B(n_394),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_332),
.B(n_372),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_300),
.B(n_331),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_278),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_262),
.A2(n_270),
.B1(n_271),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_264),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_SL g420 ( 
.A1(n_264),
.A2(n_408),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_292),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_293),
.C(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_282),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_298),
.B2(n_299),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_322),
.B(n_330),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_308),
.B(n_321),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_310),
.Y(n_324)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_319),
.A2(n_358),
.B(n_363),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_328),
.Y(n_330)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_334),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_356),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_341),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_341),
.C(n_356),
.Y(n_374)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_346),
.A2(n_366),
.A3(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_365)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_347),
.Y(n_402)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_365),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_365),
.Y(n_379)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_374),
.B(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_380),
.B2(n_393),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_379),
.C(n_393),
.Y(n_396)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_385),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_386),
.C(n_387),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_388),
.Y(n_411)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_396),
.B(n_397),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_417),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_398)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_399),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_409),
.B2(n_410),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_401),
.B(n_409),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_403),
.A3(n_404),
.B1(n_407),
.B2(n_408),
.Y(n_401)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_414),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_414),
.B(n_416),
.C(n_417),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_423),
.B2(n_432),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_418),
.B(n_424),
.C(n_427),
.Y(n_480)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_427),
.Y(n_423)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_457),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_SL g490 ( 
.A1(n_435),
.A2(n_457),
.B(n_491),
.C(n_494),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_454),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_436),
.B(n_454),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.C(n_441),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_437),
.B(n_439),
.CI(n_441),
.CON(n_470),
.SN(n_470)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_449),
.C(n_452),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_445),
.Y(n_479)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_452),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_470),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_470),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_464),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_460),
.B1(n_463),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.C(n_468),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_467),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_470),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_473),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_481),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.C(n_480),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_486),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_496),
.Y(n_499)
);

INVx13_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);


endmodule