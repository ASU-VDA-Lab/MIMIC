module fake_jpeg_28732_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_0),
.CON(n_43),
.SN(n_43)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_46),
.Y(n_89)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_21),
.B(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_70),
.B1(n_76),
.B2(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_30),
.B1(n_15),
.B2(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_32),
.B1(n_22),
.B2(n_15),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_27),
.B1(n_32),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_54),
.B1(n_50),
.B2(n_53),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_60),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_92),
.B(n_103),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_55),
.B1(n_40),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_93),
.A2(n_126),
.B1(n_73),
.B2(n_87),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_63),
.A2(n_49),
.B1(n_59),
.B2(n_38),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_58),
.B(n_14),
.C(n_26),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_110),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_106),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_41),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_113),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_25),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_114),
.C(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_28),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_67),
.C(n_62),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_19),
.B1(n_25),
.B2(n_37),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_68),
.B(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_25),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_8),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_25),
.C(n_48),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_37),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_37),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_69),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_131),
.B1(n_73),
.B2(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_37),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_65),
.B(n_2),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_136),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_159),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_87),
.B1(n_68),
.B2(n_91),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_153),
.B1(n_128),
.B2(n_116),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_154),
.B1(n_158),
.B2(n_163),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_107),
.B1(n_106),
.B2(n_103),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_95),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_8),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_92),
.A2(n_120),
.B1(n_113),
.B2(n_114),
.Y(n_163)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_92),
.B(n_117),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_169),
.A2(n_170),
.B(n_195),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_119),
.B(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_111),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_102),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_177),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_144),
.B1(n_152),
.B2(n_142),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_105),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_102),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g211 ( 
.A(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_112),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_121),
.C(n_118),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_188),
.C(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_140),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_97),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_122),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_135),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_104),
.B(n_98),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_195),
.B(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_166),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_100),
.B(n_96),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_SL g196 ( 
.A(n_146),
.B(n_154),
.C(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_139),
.B(n_152),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_143),
.B1(n_144),
.B2(n_136),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_206),
.B1(n_209),
.B2(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_193),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_208),
.B1(n_192),
.B2(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_144),
.B1(n_108),
.B2(n_134),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_138),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_210),
.C(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_134),
.B1(n_162),
.B2(n_138),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_167),
.A2(n_162),
.B1(n_172),
.B2(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_213),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_187),
.B(n_168),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_171),
.C(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_167),
.A2(n_175),
.B1(n_174),
.B2(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_168),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_184),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_173),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_218),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_238),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_227),
.A2(n_235),
.B(n_202),
.Y(n_266)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_189),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_198),
.A2(n_175),
.B1(n_182),
.B2(n_185),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_237),
.B1(n_246),
.B2(n_213),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_206),
.B1(n_223),
.B2(n_203),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_236),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_178),
.B1(n_191),
.B2(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_178),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_205),
.A3(n_222),
.B1(n_217),
.B2(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_242),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_243),
.Y(n_267)
);

OR2x6_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_224),
.Y(n_244)
);

BUFx4f_ASAP7_75t_SL g251 ( 
.A(n_244),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_218),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_207),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_256),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_210),
.C(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.C(n_260),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_201),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_226),
.B1(n_237),
.B2(n_247),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_213),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_233),
.B1(n_243),
.B2(n_247),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_202),
.C(n_200),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_257),
.C(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_264),
.B(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_280),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_276),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_226),
.B1(n_232),
.B2(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_272),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_279),
.B1(n_283),
.B2(n_253),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_246),
.B1(n_240),
.B2(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_239),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_282),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_255),
.B(n_234),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_254),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_278),
.C(n_273),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_252),
.C(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_290),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_260),
.C(n_267),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_251),
.A3(n_255),
.B1(n_262),
.B2(n_253),
.C1(n_254),
.C2(n_243),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_292),
.A2(n_271),
.B(n_281),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_278),
.C(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_290),
.C(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_276),
.C(n_283),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_299),
.B(n_288),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_277),
.C(n_279),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_274),
.B1(n_268),
.B2(n_275),
.C(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_211),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_238),
.C(n_211),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_307),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_228),
.B(n_231),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_200),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_308),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_200),
.B(n_304),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.Y(n_318)
);


endmodule