module real_jpeg_30864_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_0),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_0),
.B(n_122),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_0),
.B(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_1),
.Y(n_122)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_1),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_2),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_25),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_2),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_2),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

AND2x4_ASAP7_75t_SL g97 ( 
.A(n_3),
.B(n_98),
.Y(n_97)
);

NAND2x1_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_122),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_4),
.B(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_8),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_8),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_8),
.B(n_119),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_8),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_9),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_10),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_10),
.B(n_96),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_15),
.B1(n_106),
.B2(n_111),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_R g143 ( 
.A(n_10),
.B(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_10),
.B(n_216),
.Y(n_215)
);

NAND2x1_ASAP7_75t_L g258 ( 
.A(n_10),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_10),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_13),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_13),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_13),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_13),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_13),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_15),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_15),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_16),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_17),
.B(n_175),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_149),
.CI(n_197),
.CON(n_18),
.SN(n_18)
);

HB1xp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.C(n_126),
.Y(n_20)
);

AOI221xp5_ASAP7_75t_L g199 ( 
.A1(n_21),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.C(n_203),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_21),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_21),
.B(n_200),
.Y(n_344)
);

XOR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_22),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_49),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_23),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_33),
.C(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_28),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_32),
.Y(n_141)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_32),
.Y(n_162)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_39),
.B(n_50),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_40),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_221)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_45),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_45),
.Y(n_306)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_48),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_48),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.C(n_59),
.Y(n_50)
);

XNOR2x1_ASAP7_75t_SL g209 ( 
.A(n_51),
.B(n_55),
.Y(n_209)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_59),
.B(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_89),
.B2(n_90),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_64),
.B(n_152),
.C(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_70),
.Y(n_322)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_84),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_79),
.B1(n_84),
.B2(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_87),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_88),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_95),
.C(n_100),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_93),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_126),
.Y(n_200)
);

XOR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_116),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_114),
.B2(n_115),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_114),
.C(n_116),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_121),
.C(n_123),
.Y(n_180)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_142),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_142),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_129),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.C(n_138),
.Y(n_129)
);

XNOR2x2_ASAP7_75t_L g234 ( 
.A(n_130),
.B(n_235),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_131),
.B(n_132),
.Y(n_237)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_135),
.B(n_139),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_176),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_188),
.B1(n_189),
.B2(n_196),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_179),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_184),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_192),
.B(n_194),
.C(n_195),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_225),
.B(n_342),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_203),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_222),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_221),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_221),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_217),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_211),
.A2(n_212),
.B1(n_217),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_217),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AO21x2_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_246),
.B(n_341),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_228),
.B(n_230),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_232),
.B(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_234),
.B(n_236),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.C(n_242),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_242),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_245),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_335),
.B(n_340),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_286),
.B(n_334),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_278),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_278),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_264),
.B(n_277),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_251),
.B(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_261),
.C(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_268),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx4f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_284),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_284),
.C(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_299),
.B(n_333),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_297),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.C(n_295),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_289),
.A2(n_290),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_315),
.Y(n_332)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_290),
.B(n_314),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_295),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_316),
.B(n_330),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_301),
.A2(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_307),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_302),
.A2(n_303),
.B1(n_307),
.B2(n_308),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_302),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_323),
.B(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_338),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);


endmodule