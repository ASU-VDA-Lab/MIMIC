module fake_aes_11050_n_663 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_663);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_663;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g90 ( .A(n_80), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_88), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_87), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_23), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_24), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_45), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_72), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_57), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_75), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_11), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_29), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_59), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_14), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_19), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_21), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_84), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_24), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_55), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_50), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_60), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_31), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_22), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_77), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_85), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_64), .Y(n_117) );
CKINVDCx14_ASAP7_75t_R g118 ( .A(n_28), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_22), .Y(n_120) );
INVx2_ASAP7_75t_SL g121 ( .A(n_4), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_65), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_21), .Y(n_123) );
INVxp67_ASAP7_75t_SL g124 ( .A(n_37), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_5), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_23), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_54), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_81), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_5), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_34), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_127), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_121), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_121), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_127), .B(n_0), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVxp33_ASAP7_75t_SL g141 ( .A(n_93), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_96), .Y(n_142) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_96), .A2(n_130), .B(n_111), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_118), .B(n_1), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_106), .B(n_1), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_106), .B(n_2), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_125), .B(n_2), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_98), .B(n_3), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_101), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_99), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_101), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_125), .B(n_3), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_126), .Y(n_157) );
OAI22xp5_ASAP7_75t_SL g158 ( .A1(n_94), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_157), .B(n_126), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_134), .B(n_110), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_132), .B(n_107), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_134), .B(n_110), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_157), .B(n_129), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
INVxp67_ASAP7_75t_SL g167 ( .A(n_144), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_139), .B(n_129), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
AO22x2_ASAP7_75t_L g170 ( .A1(n_139), .A2(n_130), .B1(n_112), .B2(n_122), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_136), .B(n_111), .Y(n_172) );
INVxp67_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
AND2x6_ASAP7_75t_L g174 ( .A(n_145), .B(n_112), .Y(n_174) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_143), .B(n_114), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_136), .B(n_114), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx8_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
NAND3x1_ASAP7_75t_L g182 ( .A(n_139), .B(n_116), .C(n_117), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_144), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_131), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_137), .B(n_116), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_137), .B(n_117), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_132), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_145), .B(n_113), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
AND2x4_ASAP7_75t_SL g195 ( .A(n_147), .B(n_95), .Y(n_195) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_179), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_174), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_179), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_168), .B(n_147), .Y(n_201) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
OAI21xp33_ASAP7_75t_L g203 ( .A1(n_175), .A2(n_156), .B(n_154), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_195), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_174), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_166), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_170), .A2(n_147), .B1(n_153), .B2(n_156), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_174), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_187), .A2(n_143), .B(n_154), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_167), .B(n_141), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_174), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_168), .B(n_153), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_167), .B(n_153), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_170), .A2(n_133), .B1(n_158), .B2(n_146), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_174), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_173), .B(n_133), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_186), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_170), .A2(n_158), .B1(n_146), .B2(n_155), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_173), .B(n_105), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_174), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_169), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_191), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_175), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_178), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_170), .A2(n_159), .B1(n_155), .B2(n_150), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_181), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_175), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_187), .A2(n_159), .B(n_155), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_194), .B(n_159), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_170), .A2(n_150), .B1(n_149), .B2(n_135), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_194), .B(n_135), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_207), .A2(n_168), .B1(n_195), .B2(n_192), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_197), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_200), .B(n_195), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
INVx4_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
BUFx12f_ASAP7_75t_L g248 ( .A(n_201), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_199), .B(n_185), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_200), .Y(n_250) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_206), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_207), .A2(n_182), .B1(n_188), .B2(n_172), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_200), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_206), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_241), .A2(n_182), .B1(n_188), .B2(n_172), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_201), .A2(n_192), .B1(n_185), .B2(n_160), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_239), .A2(n_187), .B(n_162), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_217), .B(n_164), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_197), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_219), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_199), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_197), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_241), .A2(n_176), .B(n_187), .C(n_189), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_219), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_217), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_219), .Y(n_267) );
AOI21x1_ASAP7_75t_L g268 ( .A1(n_209), .A2(n_177), .B(n_183), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_198), .A2(n_163), .B(n_161), .C(n_189), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_206), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_211), .B(n_190), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_216), .A2(n_100), .B1(n_104), .B2(n_163), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_217), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_212), .A2(n_224), .B(n_227), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_196), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_201), .B(n_160), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_206), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_201), .B(n_160), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_228), .B(n_164), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_214), .B(n_193), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_210), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_197), .B(n_161), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_206), .Y(n_287) );
BUFx2_ASAP7_75t_SL g288 ( .A(n_197), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_222), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_248), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_255), .A2(n_214), .B1(n_236), .B2(n_202), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_262), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_243), .A2(n_221), .B1(n_216), .B2(n_229), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_264), .A2(n_218), .B(n_240), .C(n_215), .Y(n_294) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_272), .A2(n_221), .B(n_204), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_277), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_249), .B(n_204), .Y(n_297) );
OAI21x1_ASAP7_75t_SL g298 ( .A1(n_271), .A2(n_228), .B(n_225), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_255), .A2(n_214), .B1(n_202), .B2(n_229), .Y(n_299) );
BUFx10_ASAP7_75t_L g300 ( .A(n_245), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
O2A1O1Ixp5_ASAP7_75t_L g302 ( .A1(n_268), .A2(n_226), .B(n_212), .C(n_224), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_252), .A2(n_214), .B1(n_202), .B2(n_233), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_249), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_248), .B(n_233), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_271), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_248), .B(n_228), .Y(n_308) );
AND2x6_ASAP7_75t_L g309 ( .A(n_245), .B(n_208), .Y(n_309) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_284), .A2(n_203), .B(n_238), .C(n_234), .Y(n_310) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_252), .A2(n_203), .B(n_225), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_257), .A2(n_202), .B1(n_231), .B2(n_208), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_247), .Y(n_313) );
AO31x2_ASAP7_75t_L g314 ( .A1(n_284), .A2(n_234), .A3(n_238), .B(n_140), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_273), .A2(n_182), .B1(n_208), .B2(n_193), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_283), .A2(n_242), .B1(n_230), .B2(n_232), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_285), .A2(n_197), .B1(n_222), .B2(n_232), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_279), .A2(n_242), .B1(n_230), .B2(n_164), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_279), .B(n_223), .Y(n_320) );
OR2x6_ASAP7_75t_L g321 ( .A(n_245), .B(n_205), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_281), .A2(n_193), .B1(n_205), .B2(n_213), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_259), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_281), .A2(n_213), .B1(n_140), .B2(n_135), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_259), .A2(n_149), .B1(n_140), .B2(n_150), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_245), .A2(n_102), .B1(n_103), .B2(n_220), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_316), .B(n_259), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_293), .A2(n_289), .B1(n_282), .B2(n_226), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_306), .Y(n_330) );
BUFx4f_ASAP7_75t_SL g331 ( .A(n_296), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_295), .A2(n_269), .B1(n_258), .B2(n_289), .C(n_148), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_315), .A2(n_247), .B1(n_274), .B2(n_278), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_293), .A2(n_291), .B1(n_303), .B2(n_299), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_320), .A2(n_282), .B1(n_274), .B2(n_278), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_268), .B(n_276), .Y(n_336) );
AND2x6_ASAP7_75t_L g337 ( .A(n_317), .B(n_251), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_304), .A2(n_282), .B1(n_149), .B2(n_138), .C(n_142), .Y(n_338) );
HB1xp67_ASAP7_75t_SL g339 ( .A(n_290), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_307), .A2(n_282), .B1(n_123), .B2(n_120), .C1(n_138), .C2(n_142), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_319), .A2(n_138), .B1(n_142), .B2(n_261), .C(n_246), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_294), .A2(n_220), .B(n_224), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_320), .A2(n_247), .B1(n_253), .B2(n_266), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_292), .A2(n_247), .B1(n_265), .B2(n_267), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_319), .B(n_316), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_297), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
OAI33xp33_ASAP7_75t_L g350 ( .A1(n_312), .A2(n_119), .A3(n_122), .B1(n_177), .B2(n_183), .B3(n_128), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_326), .A2(n_275), .B1(n_250), .B2(n_266), .Y(n_351) );
AO31x2_ASAP7_75t_L g352 ( .A1(n_310), .A2(n_287), .A3(n_265), .B(n_267), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g353 ( .A1(n_325), .A2(n_246), .B1(n_261), .B2(n_119), .C(n_265), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_212), .B1(n_226), .B2(n_227), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_324), .A2(n_227), .B1(n_267), .B2(n_220), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_326), .B(n_286), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_286), .B1(n_275), .B2(n_250), .C(n_253), .Y(n_358) );
OAI222xp33_ASAP7_75t_L g359 ( .A1(n_334), .A2(n_305), .B1(n_308), .B2(n_327), .C1(n_313), .C2(n_321), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_346), .A2(n_311), .B1(n_322), .B2(n_310), .C(n_324), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_341), .B(n_314), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_341), .B(n_301), .Y(n_362) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_348), .B(n_305), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_352), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_337), .B(n_301), .Y(n_365) );
OAI21xp5_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_318), .B(n_313), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_323), .B1(n_308), .B2(n_305), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_348), .Y(n_368) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_354), .B(n_308), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_354), .B(n_301), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g371 ( .A1(n_340), .A2(n_321), .B1(n_124), .B2(n_115), .C(n_97), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_337), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_328), .B(n_301), .Y(n_373) );
AOI31xp33_ASAP7_75t_L g374 ( .A1(n_333), .A2(n_338), .A3(n_350), .B(n_345), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
NOR2x1_ASAP7_75t_L g376 ( .A(n_349), .B(n_288), .Y(n_376) );
OAI221xp5_ASAP7_75t_SL g377 ( .A1(n_347), .A2(n_321), .B1(n_7), .B2(n_8), .C(n_9), .Y(n_377) );
OAI33xp33_ASAP7_75t_L g378 ( .A1(n_330), .A2(n_165), .A3(n_171), .B1(n_180), .B2(n_10), .B3(n_11), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_335), .A2(n_275), .B1(n_250), .B2(n_266), .C(n_253), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_357), .A2(n_331), .B1(n_349), .B2(n_353), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_309), .B1(n_300), .B2(n_298), .C1(n_275), .C2(n_266), .Y(n_382) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_253), .B1(n_250), .B2(n_178), .C(n_263), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_352), .B(n_309), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_332), .A2(n_178), .B1(n_263), .B2(n_260), .C(n_244), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_337), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_339), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_352), .B(n_300), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_361), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_387), .B(n_344), .C(n_358), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_371), .B(n_6), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_362), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g394 ( .A1(n_371), .A2(n_351), .B(n_343), .C(n_165), .Y(n_394) );
OAI33xp33_ASAP7_75t_L g395 ( .A1(n_381), .A2(n_8), .A3(n_9), .B1(n_10), .B2(n_12), .B3(n_13), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_368), .B(n_352), .Y(n_396) );
AOI211xp5_ASAP7_75t_L g397 ( .A1(n_359), .A2(n_356), .B(n_165), .C(n_180), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g398 ( .A(n_377), .B(n_171), .C(n_180), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_362), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_374), .A2(n_336), .B(n_355), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_381), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_380), .A2(n_309), .B1(n_337), .B2(n_287), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_360), .A2(n_309), .B1(n_337), .B2(n_287), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_373), .B(n_336), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_387), .B(n_359), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_377), .B(n_367), .C(n_360), .D(n_388), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_388), .B(n_171), .C(n_13), .D(n_14), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_373), .B(n_12), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
AOI33xp33_ASAP7_75t_L g414 ( .A1(n_388), .A2(n_15), .A3(n_16), .B1(n_17), .B2(n_18), .B3(n_19), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_373), .B(n_15), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_363), .A2(n_220), .B1(n_256), .B2(n_280), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_363), .A2(n_309), .B(n_260), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_386), .Y(n_422) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_375), .B(n_251), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_376), .Y(n_424) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_384), .B(n_16), .C(n_17), .D(n_18), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_403), .Y(n_426) );
NAND2xp33_ASAP7_75t_SL g427 ( .A(n_412), .B(n_386), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_419), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_422), .B(n_384), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_417), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_389), .B(n_364), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_389), .B(n_369), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_424), .B(n_375), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_406), .B(n_375), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_390), .B(n_375), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_390), .B(n_372), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_419), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_417), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_400), .B(n_372), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_400), .B(n_369), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_393), .B(n_399), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_408), .B(n_374), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_424), .B(n_372), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_393), .B(n_365), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_399), .B(n_365), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_408), .B(n_366), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_406), .B(n_365), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_392), .B(n_382), .C(n_366), .D(n_383), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_416), .B(n_365), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_416), .B(n_365), .Y(n_451) );
AND3x1_ASAP7_75t_L g452 ( .A(n_409), .B(n_383), .C(n_385), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_401), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_385), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_407), .B(n_20), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_20), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_413), .B(n_382), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_401), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_414), .B(n_379), .C(n_181), .Y(n_460) );
AOI31xp33_ASAP7_75t_L g461 ( .A1(n_420), .A2(n_378), .A3(n_379), .B(n_244), .Y(n_461) );
OAI31xp33_ASAP7_75t_L g462 ( .A1(n_411), .A2(n_378), .A3(n_26), .B(n_27), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_396), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_402), .B(n_25), .Y(n_465) );
NOR2xp67_ASAP7_75t_SL g466 ( .A(n_425), .B(n_288), .Y(n_466) );
NOR2x1p5_ASAP7_75t_L g467 ( .A(n_410), .B(n_280), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_423), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_412), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_402), .B(n_415), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_423), .Y(n_471) );
INVxp67_ASAP7_75t_SL g472 ( .A(n_415), .Y(n_472) );
OAI31xp33_ASAP7_75t_L g473 ( .A1(n_394), .A2(n_25), .A3(n_26), .B(n_27), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_391), .B(n_28), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_405), .B(n_29), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_418), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_459), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_463), .B(n_404), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_430), .B(n_397), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_463), .B(n_421), .Y(n_481) );
NOR3xp33_ASAP7_75t_L g482 ( .A(n_475), .B(n_395), .C(n_398), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_464), .B(n_181), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_435), .B(n_181), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_459), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_428), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_426), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_428), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_435), .B(n_181), .Y(n_490) );
INVx6_ASAP7_75t_L g491 ( .A(n_468), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_429), .Y(n_492) );
INVxp33_ASAP7_75t_L g493 ( .A(n_467), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_475), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_464), .B(n_181), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_453), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_435), .B(n_181), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_442), .B(n_30), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_469), .B(n_32), .Y(n_500) );
INVxp67_ASAP7_75t_SL g501 ( .A(n_469), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_442), .B(n_33), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_445), .B(n_35), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_472), .B(n_450), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_472), .B(n_36), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_450), .B(n_38), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_443), .B(n_39), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_445), .B(n_40), .Y(n_508) );
AOI211xp5_ASAP7_75t_SL g509 ( .A1(n_461), .A2(n_42), .B(n_46), .C(n_47), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_446), .B(n_48), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_465), .B(n_49), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_453), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_451), .B(n_51), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_453), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_431), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_431), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_456), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_451), .B(n_52), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_465), .B(n_53), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_439), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_439), .Y(n_521) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_474), .A2(n_237), .B(n_58), .Y(n_522) );
AND3x2_ASAP7_75t_L g523 ( .A(n_462), .B(n_56), .C(n_61), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_433), .Y(n_524) );
AND2x4_ASAP7_75t_SL g525 ( .A(n_448), .B(n_437), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_470), .B(n_62), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_432), .B(n_63), .Y(n_528) );
NOR3xp33_ASAP7_75t_L g529 ( .A(n_460), .B(n_237), .C(n_235), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_458), .B(n_66), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_446), .B(n_67), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_470), .B(n_68), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_456), .Y(n_533) );
OAI322xp33_ASAP7_75t_L g534 ( .A1(n_494), .A2(n_474), .A3(n_441), .B1(n_455), .B2(n_457), .C1(n_447), .C2(n_440), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_478), .B(n_485), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_493), .B(n_449), .Y(n_536) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_482), .B(n_473), .C(n_462), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_504), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_525), .Y(n_539) );
INVx4_ASAP7_75t_L g540 ( .A(n_491), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_487), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_525), .B(n_448), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_523), .A2(n_473), .B(n_461), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g544 ( .A1(n_493), .A2(n_457), .B(n_455), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_501), .B(n_441), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_488), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_492), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_495), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_517), .Y(n_549) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_533), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_527), .B(n_448), .Y(n_551) );
XNOR2x1_ASAP7_75t_L g552 ( .A(n_481), .B(n_452), .Y(n_552) );
OAI221xp5_ASAP7_75t_L g553 ( .A1(n_480), .A2(n_427), .B1(n_452), .B2(n_460), .C(n_466), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_491), .B(n_471), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_509), .A2(n_466), .B(n_476), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_515), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_516), .B(n_447), .Y(n_557) );
XNOR2xp5_ASAP7_75t_L g558 ( .A(n_480), .B(n_448), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_491), .Y(n_559) );
XNOR2xp5_ASAP7_75t_L g560 ( .A(n_499), .B(n_458), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_497), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_499), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_502), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_529), .A2(n_430), .B1(n_476), .B2(n_454), .Y(n_566) );
AO22x2_ASAP7_75t_L g567 ( .A1(n_512), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_567) );
AOI32xp33_ASAP7_75t_L g568 ( .A1(n_502), .A2(n_468), .A3(n_471), .B1(n_454), .B2(n_436), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_503), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_514), .B(n_454), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_483), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_503), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_434), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_484), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_486), .B(n_477), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_526), .B(n_444), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_483), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_486), .B(n_477), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_489), .B(n_477), .Y(n_579) );
XOR2xp5_ASAP7_75t_L g580 ( .A(n_479), .B(n_69), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_526), .A2(n_280), .B(n_270), .C(n_256), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_496), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_508), .B(n_71), .Y(n_583) );
XNOR2x2_ASAP7_75t_L g584 ( .A(n_532), .B(n_73), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_496), .Y(n_585) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_507), .A2(n_74), .B(n_76), .C(n_78), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_508), .B(n_270), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_490), .B(n_79), .Y(n_589) );
XOR2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_82), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_490), .B(n_83), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_498), .B(n_86), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_513), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_510), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_518), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_89), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_531), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_531), .B(n_251), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_505), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_528), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_511), .A2(n_235), .B(n_237), .C(n_254), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_519), .Y(n_603) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_530), .A2(n_178), .B(n_254), .C(n_270), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_522), .B(n_254), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_522), .A2(n_254), .B1(n_220), .B2(n_178), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_524), .B(n_178), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_504), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_517), .B(n_220), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_529), .A2(n_235), .B(n_371), .C(n_475), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_494), .A2(n_235), .B1(n_158), .B2(n_392), .C1(n_465), .C2(n_480), .Y(n_612) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_540), .A2(n_539), .B1(n_543), .B2(n_553), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_559), .B(n_542), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_536), .A2(n_537), .B1(n_553), .B2(n_567), .C(n_534), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_535), .Y(n_616) );
XNOR2x1_ASAP7_75t_L g617 ( .A(n_552), .B(n_558), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_545), .B(n_570), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_535), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_567), .B(n_551), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_612), .A2(n_560), .B1(n_599), .B2(n_600), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_538), .A2(n_609), .B1(n_601), .B2(n_603), .Y(n_622) );
AOI311xp33_ASAP7_75t_L g623 ( .A1(n_550), .A2(n_595), .A3(n_593), .B(n_544), .C(n_597), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_572), .A2(n_594), .B1(n_569), .B2(n_576), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_611), .A2(n_555), .B(n_549), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_611), .A2(n_549), .B(n_586), .C(n_602), .Y(n_626) );
BUFx8_ASAP7_75t_L g627 ( .A(n_592), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_574), .A2(n_565), .B1(n_564), .B2(n_573), .Y(n_628) );
AOI221x1_ASAP7_75t_L g629 ( .A1(n_554), .A2(n_607), .B1(n_544), .B2(n_591), .C(n_589), .Y(n_629) );
AOI22xp5_ASAP7_75t_SL g630 ( .A1(n_583), .A2(n_580), .B1(n_590), .B2(n_584), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_568), .A2(n_566), .B1(n_610), .B2(n_581), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_570), .A2(n_582), .B1(n_585), .B2(n_571), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_615), .A2(n_606), .B(n_586), .C(n_596), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g634 ( .A1(n_613), .A2(n_588), .B(n_604), .C(n_602), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_625), .A2(n_557), .B1(n_546), .B2(n_547), .C(n_548), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_626), .B(n_608), .C(n_557), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_617), .A2(n_577), .B1(n_556), .B2(n_561), .Y(n_637) );
NOR2xp67_ASAP7_75t_L g638 ( .A(n_624), .B(n_587), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_616), .B(n_541), .Y(n_639) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_631), .B(n_605), .Y(n_640) );
NAND4xp25_ASAP7_75t_SL g641 ( .A(n_621), .B(n_579), .C(n_578), .D(n_575), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_620), .B(n_562), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_623), .A2(n_579), .B1(n_575), .B2(n_578), .C(n_563), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_637), .B(n_630), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_633), .B(n_622), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_643), .B(n_618), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_640), .A2(n_629), .B(n_628), .C(n_632), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_634), .B(n_614), .C(n_619), .D(n_598), .Y(n_648) );
XNOR2xp5_ASAP7_75t_L g649 ( .A(n_636), .B(n_627), .Y(n_649) );
INVxp67_ASAP7_75t_L g650 ( .A(n_639), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_649), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_645), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_646), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_650), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_654), .Y(n_655) );
AND3x4_ASAP7_75t_L g656 ( .A(n_652), .B(n_644), .C(n_638), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_651), .B(n_642), .Y(n_657) );
AOI22x1_ASAP7_75t_L g658 ( .A1(n_655), .A2(n_653), .B1(n_652), .B2(n_647), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_657), .Y(n_659) );
NOR2xp67_ASAP7_75t_SL g660 ( .A(n_659), .B(n_648), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_658), .Y(n_661) );
AOI22xp5_ASAP7_75t_SL g662 ( .A1(n_661), .A2(n_657), .B1(n_656), .B2(n_660), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_635), .B(n_641), .Y(n_663) );
endmodule