module fake_jpeg_28858_n_509 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_509);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_509;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_52),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_59),
.Y(n_154)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_20),
.B(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_68),
.Y(n_104)
);

NOR2xp67_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_7),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_65),
.B(n_83),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_20),
.B(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_70),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_74),
.Y(n_110)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_34),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_6),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_32),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_92),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_23),
.A2(n_14),
.B(n_6),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_0),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_102),
.B(n_111),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_40),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_49),
.B(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_51),
.B(n_35),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_113),
.B(n_28),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_35),
.B1(n_45),
.B2(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_45),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_61),
.A2(n_30),
.B1(n_43),
.B2(n_34),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_128),
.B1(n_144),
.B2(n_153),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_43),
.B1(n_34),
.B2(n_15),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_90),
.Y(n_178)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_95),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_143),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_75),
.A2(n_19),
.B1(n_18),
.B2(n_46),
.Y(n_144)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_155),
.A2(n_192),
.B1(n_196),
.B2(n_33),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_71),
.C(n_80),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_159),
.B(n_82),
.Y(n_225)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_162),
.A2(n_144),
.B1(n_125),
.B2(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_24),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_174),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_40),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_165),
.B(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_172),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_42),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_16),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_16),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_200),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_19),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_19),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_98),
.A2(n_31),
.B1(n_94),
.B2(n_33),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_142),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_82),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_195),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_98),
.A2(n_33),
.B1(n_15),
.B2(n_84),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_18),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_19),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_112),
.A2(n_33),
.B1(n_96),
.B2(n_97),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_141),
.Y(n_204)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_24),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_203),
.C(n_28),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_135),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_231),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_127),
.B1(n_122),
.B2(n_146),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_213),
.A2(n_214),
.B1(n_167),
.B2(n_198),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_127),
.B1(n_146),
.B2(n_147),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_226),
.B1(n_236),
.B2(n_237),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_157),
.A2(n_112),
.B1(n_129),
.B2(n_76),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_167),
.B1(n_133),
.B2(n_169),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_151),
.B1(n_149),
.B2(n_147),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_165),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_158),
.A2(n_141),
.B1(n_39),
.B2(n_23),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_234),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_160),
.A2(n_151),
.B1(n_149),
.B2(n_145),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_145),
.B1(n_137),
.B2(n_136),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_159),
.A2(n_137),
.B1(n_55),
.B2(n_66),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_239),
.A2(n_125),
.B1(n_168),
.B2(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_174),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_186),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_254),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_155),
.B(n_164),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_245),
.A2(n_255),
.B(n_271),
.Y(n_286)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_248),
.B(n_207),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_264),
.Y(n_281)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_251),
.A2(n_261),
.B(n_227),
.Y(n_299)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_253),
.Y(n_297)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_223),
.B(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_171),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_258),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_226),
.B1(n_236),
.B2(n_239),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_205),
.B(n_166),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_209),
.A2(n_185),
.B1(n_133),
.B2(n_181),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_172),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_265),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_187),
.B1(n_170),
.B2(n_197),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_206),
.B1(n_242),
.B2(n_221),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_231),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_181),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_276),
.B1(n_235),
.B2(n_217),
.Y(n_289)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_205),
.B(n_170),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_271),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_223),
.B(n_191),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_273),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_190),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_189),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_275),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_189),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_222),
.A2(n_179),
.B1(n_50),
.B2(n_139),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_179),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_279),
.B(n_233),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_248),
.C(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_313),
.C(n_268),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_304),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_206),
.B1(n_209),
.B2(n_213),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_288),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_272),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_289),
.A2(n_302),
.B1(n_310),
.B2(n_244),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_217),
.B(n_220),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_292),
.A2(n_133),
.B(n_244),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_267),
.B(n_257),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_238),
.B(n_227),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_300),
.A2(n_273),
.B(n_274),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_246),
.B1(n_259),
.B2(n_249),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_259),
.A2(n_220),
.B1(n_242),
.B2(n_221),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_266),
.A2(n_234),
.B1(n_238),
.B2(n_193),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_308),
.A2(n_312),
.B1(n_263),
.B2(n_269),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_311),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_234),
.B1(n_203),
.B2(n_161),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_258),
.B(n_177),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_246),
.A2(n_234),
.B1(n_177),
.B2(n_199),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_245),
.C(n_275),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_315),
.A2(n_319),
.B(n_324),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_243),
.C(n_265),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_320),
.B(n_329),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_296),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_262),
.Y(n_323)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_254),
.Y(n_324)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_326),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_299),
.A2(n_252),
.B1(n_278),
.B2(n_247),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_327),
.A2(n_297),
.B1(n_280),
.B2(n_303),
.Y(n_376)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_291),
.B(n_256),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_339),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_331),
.A2(n_344),
.B1(n_283),
.B2(n_310),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_247),
.B(n_276),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_336),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_23),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_333),
.B(n_343),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_254),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_298),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_260),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_338),
.B(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_284),
.A2(n_278),
.B(n_215),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_341),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_293),
.B(n_286),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_346),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_307),
.B(n_46),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_285),
.B(n_253),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.Y(n_354)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_334),
.B(n_306),
.CI(n_287),
.CON(n_350),
.SN(n_350)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_19),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_321),
.C(n_325),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_337),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_353),
.B(n_360),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_355),
.A2(n_322),
.B1(n_343),
.B2(n_339),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_331),
.A2(n_287),
.B1(n_304),
.B2(n_309),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_356),
.A2(n_361),
.B1(n_378),
.B2(n_338),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_318),
.A2(n_308),
.B1(n_312),
.B2(n_292),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_358),
.A2(n_376),
.B1(n_370),
.B2(n_367),
.Y(n_382)
);

AOI22x1_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_314),
.B1(n_289),
.B2(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_337),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_319),
.A2(n_298),
.B1(n_311),
.B2(n_306),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_290),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_369),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_368),
.B(n_361),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_294),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_314),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_370),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_374),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_333),
.B(n_46),
.Y(n_377)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_12),
.C(n_11),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_345),
.A2(n_340),
.B1(n_324),
.B2(n_315),
.Y(n_378)
);

OA22x2_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_215),
.B1(n_250),
.B2(n_253),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_380),
.A2(n_345),
.B(n_330),
.C(n_317),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_382),
.A2(n_407),
.B1(n_378),
.B2(n_356),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_391),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_384),
.A2(n_389),
.B1(n_398),
.B2(n_354),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_335),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_386),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_334),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_364),
.A2(n_321),
.B(n_341),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_387),
.A2(n_405),
.B(n_371),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_316),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_381),
.B(n_348),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_396),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_397),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_357),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_355),
.A2(n_138),
.B1(n_250),
.B2(n_53),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_399),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_372),
.A2(n_39),
.B1(n_87),
.B2(n_85),
.Y(n_400)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_400),
.Y(n_413)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_401),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_349),
.B(n_39),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_409),
.B1(n_373),
.B2(n_374),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_364),
.A2(n_354),
.B(n_366),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_79),
.C(n_92),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_397),
.C(n_386),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_358),
.A2(n_103),
.B1(n_81),
.B2(n_91),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_408),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_430),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_422),
.B1(n_425),
.B2(n_429),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_385),
.C(n_395),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_420),
.C(n_426),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_431),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_362),
.C(n_354),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_370),
.B1(n_369),
.B2(n_359),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_392),
.A2(n_369),
.B1(n_359),
.B2(n_366),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_403),
.C(n_387),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_427),
.A2(n_394),
.B(n_371),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_394),
.A2(n_380),
.B1(n_363),
.B2(n_365),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_350),
.Y(n_430)
);

FAx1_ASAP7_75t_SL g431 ( 
.A(n_403),
.B(n_388),
.CI(n_407),
.CON(n_431),
.SN(n_431)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_403),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_435),
.B(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_418),
.C(n_428),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_438),
.C(n_447),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_399),
.C(n_401),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_408),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_440),
.B(n_70),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_424),
.B(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_442),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_426),
.A2(n_383),
.B(n_380),
.Y(n_444)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

NAND2x1_ASAP7_75t_SL g446 ( 
.A(n_431),
.B(n_380),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_446),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_398),
.C(n_373),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_414),
.B(n_379),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_449),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_425),
.B(n_379),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_422),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_451),
.C(n_8),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_415),
.C(n_423),
.Y(n_451)
);

BUFx24_ASAP7_75t_SL g452 ( 
.A(n_433),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_452),
.B(n_437),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_434),
.A2(n_432),
.B(n_421),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_453),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_445),
.A2(n_413),
.B1(n_429),
.B2(n_416),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_459),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_390),
.B1(n_89),
.B2(n_78),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_456),
.A2(n_465),
.B1(n_466),
.B2(n_436),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_447),
.A2(n_52),
.B1(n_118),
.B2(n_3),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_461),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_8),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_8),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_462),
.A2(n_11),
.B(n_9),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_450),
.A2(n_8),
.B1(n_12),
.B2(n_3),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_449),
.B1(n_446),
.B2(n_448),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_9),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_477),
.Y(n_490)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_457),
.A2(n_468),
.B(n_463),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_476),
.B(n_482),
.Y(n_484)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_441),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_479),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_434),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_482),
.Y(n_492)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_435),
.C(n_22),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_481),
.C(n_465),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_464),
.C(n_466),
.Y(n_481)
);

INVx6_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_470),
.C(n_473),
.Y(n_494)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_484),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_476),
.A2(n_454),
.B(n_5),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_485),
.B(n_486),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_454),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_3),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_5),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_492),
.B(n_480),
.C(n_479),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_494),
.C(n_491),
.Y(n_501)
);

AOI21xp33_ASAP7_75t_L g495 ( 
.A1(n_492),
.A2(n_471),
.B(n_4),
.Y(n_495)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_495),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_497),
.A2(n_489),
.B(n_488),
.C(n_491),
.Y(n_499)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_499),
.A2(n_502),
.A3(n_496),
.B1(n_493),
.B2(n_2),
.C1(n_0),
.C2(n_44),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_501),
.A2(n_2),
.B(n_44),
.Y(n_504)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g502 ( 
.A1(n_498),
.A2(n_490),
.B(n_5),
.C(n_44),
.D(n_22),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_504),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_505),
.B(n_500),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_2),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_507),
.A2(n_2),
.B(n_44),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_44),
.Y(n_509)
);


endmodule