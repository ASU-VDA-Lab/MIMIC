module fake_jpeg_19839_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_21),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_29),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_21),
.B(n_20),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_36),
.C(n_40),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_31),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_19),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_20),
.B1(n_17),
.B2(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_0),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_19),
.B1(n_31),
.B2(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_39),
.B1(n_34),
.B2(n_20),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_32),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_71),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_17),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_65),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_67)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_68),
.B(n_77),
.Y(n_95)
);

NAND4xp25_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_20),
.C(n_21),
.D(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_39),
.C(n_34),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_81),
.B1(n_83),
.B2(n_87),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_16),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_47),
.B1(n_53),
.B2(n_52),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_81)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_21),
.B1(n_18),
.B2(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_18),
.B1(n_31),
.B2(n_28),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_99),
.B(n_49),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_51),
.B1(n_49),
.B2(n_82),
.Y(n_133)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_98),
.Y(n_117)
);

CKINVDCx9p33_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_70),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_63),
.A2(n_56),
.B(n_18),
.Y(n_100)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_100),
.B(n_112),
.CON(n_118),
.SN(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_18),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_105),
.B(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_13),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_79),
.A2(n_55),
.B1(n_53),
.B2(n_52),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_70),
.B1(n_60),
.B2(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_71),
.B(n_34),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_77),
.B(n_72),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_59),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_22),
.A3(n_31),
.B1(n_49),
.B2(n_51),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_67),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_129),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_67),
.B1(n_69),
.B2(n_85),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_119),
.B1(n_91),
.B2(n_106),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_67),
.B1(n_61),
.B2(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_120),
.A2(n_133),
.B1(n_97),
.B2(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_142),
.B(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_86),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_75),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_70),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_51),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_139),
.B(n_102),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_22),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_93),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_144),
.B(n_156),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_100),
.B(n_88),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_153),
.B1(n_117),
.B2(n_128),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_154),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_95),
.B(n_111),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_159),
.B1(n_167),
.B2(n_135),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_95),
.B1(n_96),
.B2(n_114),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_95),
.B(n_98),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_101),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_108),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_105),
.B1(n_89),
.B2(n_113),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_99),
.B(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_115),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_97),
.B1(n_74),
.B2(n_60),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_74),
.C(n_60),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_121),
.C(n_125),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_0),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_140),
.B(n_117),
.C(n_139),
.D(n_121),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_169),
.C(n_146),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_187),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_128),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_152),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_194),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_195),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_193),
.A2(n_196),
.B1(n_159),
.B2(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_22),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_162),
.B1(n_150),
.B2(n_143),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_201),
.C(n_202),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_210),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_154),
.C(n_148),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_166),
.C(n_170),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_183),
.B1(n_181),
.B2(n_188),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_150),
.C(n_151),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_165),
.B1(n_160),
.B2(n_167),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_189),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_160),
.B1(n_8),
.B2(n_2),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_82),
.C(n_7),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_184),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_199),
.A2(n_182),
.B1(n_192),
.B2(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_187),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_174),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_181),
.B1(n_172),
.B2(n_195),
.Y(n_223)
);

OAI321xp33_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_5),
.A3(n_14),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_15),
.B(n_9),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_229),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_11),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_206),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_3),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_213),
.A2(n_4),
.B1(n_9),
.B2(n_12),
.Y(n_231)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_1),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_236),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_201),
.C(n_209),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_243),
.C(n_226),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_209),
.C(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_228),
.Y(n_246)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_236),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_243),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_203),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_254),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_220),
.B(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_253),
.B(n_239),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_225),
.B1(n_227),
.B2(n_232),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_261),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_258),
.A2(n_247),
.B1(n_249),
.B2(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_263),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_233),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_250),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_267),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_1),
.A3(n_14),
.B1(n_15),
.B2(n_260),
.C1(n_263),
.C2(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_15),
.B(n_1),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_264),
.C(n_273),
.Y(n_274)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_274),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_276),
.B(n_275),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_271),
.Y(n_278)
);


endmodule