module fake_netlist_1_2583_n_1090 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1090);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1090;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_476;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_769;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_828;
wire n_767;
wire n_1063;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_262;
wire n_556;
wire n_601;
wire n_439;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_260;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1088;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_269;
INVx2_ASAP7_75t_L g246 ( .A(n_121), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_63), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_242), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_237), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_60), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_107), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_103), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_55), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_122), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_236), .B(n_219), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_18), .Y(n_257) );
NOR2xp67_ASAP7_75t_L g258 ( .A(n_134), .B(n_166), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_214), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_57), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_172), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_102), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_77), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_159), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_59), .Y(n_266) );
INVxp33_ASAP7_75t_L g267 ( .A(n_99), .Y(n_267) );
INVxp33_ASAP7_75t_SL g268 ( .A(n_53), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_131), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_111), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_113), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_157), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_57), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
INVxp67_ASAP7_75t_SL g275 ( .A(n_44), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_43), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_50), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_84), .Y(n_278) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_86), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_167), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_110), .Y(n_281) );
INVxp33_ASAP7_75t_L g282 ( .A(n_198), .Y(n_282) );
INVxp67_ASAP7_75t_L g283 ( .A(n_64), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_42), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_155), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_25), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_67), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_112), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_38), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_161), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_243), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_245), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_240), .Y(n_295) );
CKINVDCx14_ASAP7_75t_R g296 ( .A(n_48), .Y(n_296) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_241), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_105), .Y(n_298) );
INVxp67_ASAP7_75t_L g299 ( .A(n_127), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_197), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_217), .Y(n_301) );
INVxp33_ASAP7_75t_SL g302 ( .A(n_210), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_164), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_177), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_126), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_124), .Y(n_306) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_201), .Y(n_307) );
INVxp67_ASAP7_75t_SL g308 ( .A(n_141), .Y(n_308) );
INVxp33_ASAP7_75t_L g309 ( .A(n_66), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_220), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_211), .Y(n_311) );
INVxp33_ASAP7_75t_L g312 ( .A(n_59), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_117), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_185), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_52), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_128), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_139), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_176), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_151), .Y(n_319) );
BUFx2_ASAP7_75t_SL g320 ( .A(n_196), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_94), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_238), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_100), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_213), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_72), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_205), .Y(n_326) );
BUFx2_ASAP7_75t_SL g327 ( .A(n_163), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_106), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_223), .B(n_49), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_5), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_39), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_36), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_184), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_186), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_218), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_212), .Y(n_336) );
INVxp33_ASAP7_75t_SL g337 ( .A(n_26), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_76), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_18), .Y(n_339) );
INVxp33_ASAP7_75t_SL g340 ( .A(n_108), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_193), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_239), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_4), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_11), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_200), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_140), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_203), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_76), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_61), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_39), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_221), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_43), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_199), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_63), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_28), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_150), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_90), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_48), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_147), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_145), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_21), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_37), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_89), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_78), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_202), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_22), .Y(n_366) );
CKINVDCx14_ASAP7_75t_R g367 ( .A(n_104), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_0), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_189), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_45), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_55), .Y(n_371) );
INVxp33_ASAP7_75t_SL g372 ( .A(n_215), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_190), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_309), .B(n_0), .Y(n_374) );
OR2x6_ASAP7_75t_L g375 ( .A(n_320), .B(n_1), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_285), .B(n_1), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_265), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_265), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_269), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_247), .B(n_2), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_247), .B(n_2), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_269), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g384 ( .A(n_297), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_271), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_336), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_271), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_293), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_315), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_296), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_272), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_336), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_336), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_264), .B(n_3), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_336), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_267), .B(n_3), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_272), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_246), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_348), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_293), .Y(n_400) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_305), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_274), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_274), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_280), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_312), .B(n_4), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_378), .B(n_282), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_375), .A2(n_337), .B1(n_268), .B2(n_287), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_400), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_388), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_388), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_378), .B(n_277), .Y(n_412) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_381), .B(n_280), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_390), .B(n_250), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_390), .B(n_299), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_398), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_398), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_384), .B(n_250), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_384), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
BUFx4_ASAP7_75t_L g422 ( .A(n_377), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_381), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_375), .A2(n_337), .B1(n_268), .B2(n_287), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_379), .B(n_277), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_381), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_382), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_388), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_382), .B(n_251), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_392), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_380), .B(n_302), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_385), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_392), .Y(n_443) );
OR2x6_ASAP7_75t_L g444 ( .A(n_375), .B(n_320), .Y(n_444) );
BUFx4f_ASAP7_75t_L g445 ( .A(n_444), .Y(n_445) );
INVx5_ASAP7_75t_L g446 ( .A(n_444), .Y(n_446) );
BUFx8_ASAP7_75t_L g447 ( .A(n_422), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_407), .B(n_377), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_444), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_442), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_444), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_444), .B(n_375), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g453 ( .A(n_413), .B(n_248), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_407), .B(n_252), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_440), .B(n_406), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_423), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_428), .A2(n_375), .B1(n_405), .B2(n_374), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_442), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_416), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_416), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_422), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_412), .B(n_374), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_423), .A2(n_375), .B1(n_405), .B2(n_402), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
INVx1_ASAP7_75t_SL g475 ( .A(n_429), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_438), .B(n_375), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_425), .B(n_252), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_438), .Y(n_478) );
BUFx4f_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_421), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_426), .B(n_427), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_426), .B(n_385), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_427), .A2(n_385), .B1(n_402), .B2(n_387), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_430), .B(n_396), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_415), .B(n_399), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_432), .B(n_383), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_408), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_432), .B(n_295), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_419), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_436), .B(n_383), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_414), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_411), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_408), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_437), .B(n_295), .Y(n_499) );
INVx1_ASAP7_75t_SL g500 ( .A(n_437), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_441), .A2(n_394), .B1(n_404), .B2(n_397), .C(n_391), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_441), .B(n_402), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_433), .B(n_387), .Y(n_503) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_433), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_433), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_409), .B(n_391), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_409), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_418), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_418), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_424), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
AND3x1_ASAP7_75t_L g512 ( .A(n_431), .B(n_394), .C(n_397), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_431), .A2(n_403), .B1(n_404), .B2(n_388), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_461), .Y(n_514) );
BUFx12f_ASAP7_75t_L g515 ( .A(n_447), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_455), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_446), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_469), .B(n_403), .Y(n_519) );
BUFx2_ASAP7_75t_L g520 ( .A(n_455), .Y(n_520) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_455), .Y(n_521) );
BUFx8_ASAP7_75t_L g522 ( .A(n_452), .Y(n_522) );
BUFx4_ASAP7_75t_SL g523 ( .A(n_447), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_455), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_289), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_461), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_457), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_446), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_461), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_457), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_463), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_447), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_475), .B(n_396), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_457), .B(n_275), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_447), .Y(n_537) );
OAI21xp33_ASAP7_75t_L g538 ( .A1(n_472), .A2(n_357), .B(n_340), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_467), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_463), .Y(n_540) );
BUFx3_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_445), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_469), .B(n_289), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_465), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_448), .B(n_399), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_465), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_450), .A2(n_443), .B(n_431), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_474), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_445), .A2(n_311), .B1(n_270), .B2(n_276), .Y(n_552) );
AND2x4_ASAP7_75t_SL g553 ( .A(n_452), .B(n_338), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_467), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
INVx5_ASAP7_75t_L g558 ( .A(n_446), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_480), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_452), .B(n_279), .Y(n_560) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_451), .B(n_476), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_445), .A2(n_358), .B1(n_349), .B2(n_357), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_480), .Y(n_563) );
OAI222xp33_ASAP7_75t_L g564 ( .A1(n_460), .A2(n_454), .B1(n_355), .B2(n_371), .C1(n_332), .C2(n_475), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_495), .B(n_340), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_466), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_500), .A2(n_372), .B1(n_367), .B2(n_355), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_453), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_456), .B(n_332), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_450), .A2(n_443), .B(n_307), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_476), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_485), .B(n_371), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_466), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_485), .B(n_283), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_462), .A2(n_443), .B(n_281), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_485), .A2(n_266), .B1(n_273), .B2(n_264), .Y(n_576) );
BUFx2_ASAP7_75t_L g577 ( .A(n_449), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_500), .B(n_266), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_458), .B(n_273), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_470), .Y(n_580) );
O2A1O1Ixp5_ASAP7_75t_L g581 ( .A1(n_459), .A2(n_308), .B(n_314), .C(n_306), .Y(n_581) );
INVx5_ASAP7_75t_L g582 ( .A(n_464), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_512), .A2(n_284), .B1(n_286), .B2(n_278), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_470), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_512), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_484), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_458), .B(n_278), .Y(n_587) );
AND2x4_ASAP7_75t_SL g588 ( .A(n_458), .B(n_284), .Y(n_588) );
CKINVDCx6p67_ASAP7_75t_R g589 ( .A(n_477), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_464), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_458), .A2(n_254), .B1(n_261), .B2(n_257), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_473), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_459), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_484), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_493), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_490), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_479), .Y(n_597) );
BUFx2_ASAP7_75t_L g598 ( .A(n_479), .Y(n_598) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_464), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_546), .A2(n_479), .B1(n_486), .B2(n_478), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_552), .A2(n_479), .B1(n_501), .B2(n_499), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_579), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_519), .B(n_473), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_553), .A2(n_482), .B1(n_498), .B2(n_478), .Y(n_604) );
BUFx2_ASAP7_75t_SL g605 ( .A(n_558), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_519), .B(n_483), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g607 ( .A1(n_544), .A2(n_553), .B1(n_515), .B2(n_569), .C1(n_564), .C2(n_562), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_516), .Y(n_608) );
BUFx2_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_525), .B(n_473), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_533), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_585), .A2(n_482), .B1(n_502), .B2(n_462), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_579), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_540), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
AO31x2_ASAP7_75t_L g617 ( .A1(n_566), .A2(n_491), .A3(n_492), .B(n_487), .Y(n_617) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_525), .A2(n_491), .B(n_487), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_560), .A2(n_478), .B1(n_492), .B2(n_481), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_502), .B(n_494), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_560), .A2(n_478), .B1(n_488), .B2(n_505), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_538), .A2(n_506), .B1(n_503), .B2(n_513), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_579), .Y(n_623) );
INVx3_ASAP7_75t_L g624 ( .A(n_516), .Y(n_624) );
CKINVDCx16_ASAP7_75t_R g625 ( .A(n_515), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_587), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_544), .B(n_464), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_560), .A2(n_464), .B1(n_496), .B2(n_471), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_581), .B(n_401), .C(n_400), .Y(n_629) );
AND2x4_ASAP7_75t_L g630 ( .A(n_520), .B(n_464), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_540), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_587), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_583), .A2(n_364), .B1(n_366), .B2(n_362), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_560), .A2(n_471), .B1(n_504), .B2(n_496), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_514), .B(n_471), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_548), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_538), .A2(n_325), .B(n_331), .C(n_330), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_548), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_568), .A2(n_327), .B1(n_323), .B2(n_326), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_583), .B(n_401), .C(n_400), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_571), .A2(n_496), .B1(n_504), .B2(n_471), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_514), .B(n_471), .Y(n_643) );
INVxp33_ASAP7_75t_L g644 ( .A(n_555), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_551), .Y(n_645) );
OR2x6_ASAP7_75t_L g646 ( .A(n_520), .B(n_471), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_526), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_522), .A2(n_507), .B1(n_324), .B2(n_326), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_539), .B(n_362), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_556), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_543), .A2(n_504), .B1(n_496), .B2(n_507), .Y(n_652) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_537), .A2(n_366), .B1(n_368), .B2(n_364), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_530), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_543), .A2(n_504), .B1(n_496), .B2(n_327), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_537), .A2(n_370), .B1(n_368), .B2(n_323), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_556), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_561), .A2(n_504), .B1(n_496), .B2(n_339), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_557), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_578), .B(n_504), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_561), .A2(n_343), .B1(n_350), .B2(n_344), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_545), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_554), .A2(n_370), .B1(n_333), .B2(n_359), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_566), .A2(n_509), .B(n_510), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_575), .A2(n_511), .B(n_497), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_557), .Y(n_666) );
CKINVDCx11_ASAP7_75t_R g667 ( .A(n_523), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_576), .A2(n_352), .B(n_354), .C(n_251), .Y(n_668) );
INVx4_ASAP7_75t_L g669 ( .A(n_516), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_534), .Y(n_670) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_536), .B(n_288), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_547), .Y(n_672) );
OAI22x1_ASAP7_75t_L g673 ( .A1(n_576), .A2(n_356), .B1(n_363), .B2(n_288), .Y(n_673) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_567), .A2(n_360), .B1(n_317), .B2(n_305), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_536), .A2(n_577), .B1(n_521), .B2(n_527), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_559), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_516), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_563), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_547), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_516), .B(n_363), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_595), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_563), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_595), .A2(n_361), .B1(n_315), .B2(n_365), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g684 ( .A1(n_535), .A2(n_361), .B1(n_315), .B2(n_365), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_521), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_550), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_591), .A2(n_258), .B(n_256), .C(n_369), .Y(n_687) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_521), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_536), .A2(n_361), .B1(n_315), .B2(n_369), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_577), .A2(n_361), .B1(n_249), .B2(n_255), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_521), .B(n_511), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_527), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_565), .A2(n_322), .B1(n_304), .B2(n_310), .C(n_253), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_527), .A2(n_259), .B1(n_262), .B2(n_260), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_572), .B(n_5), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_604), .A2(n_588), .B1(n_550), .B2(n_578), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_665), .A2(n_584), .B(n_580), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_609), .B(n_574), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_667), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_613), .A2(n_596), .B(n_524), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_662), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g702 ( .A1(n_633), .A2(n_667), .B1(n_606), .B2(n_610), .C1(n_653), .C2(n_673), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_618), .A2(n_584), .B1(n_573), .B2(n_586), .C(n_594), .Y(n_703) );
OAI21xp5_ASAP7_75t_L g704 ( .A1(n_641), .A2(n_570), .B(n_594), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_620), .A2(n_549), .B(n_599), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_691), .A2(n_497), .B(n_489), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_669), .B(n_527), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_662), .Y(n_708) );
OAI322xp33_ASAP7_75t_L g709 ( .A1(n_693), .A2(n_329), .A3(n_263), .B1(n_373), .B2(n_290), .C1(n_291), .C2(n_292), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_686), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_673), .A2(n_542), .B1(n_532), .B2(n_531), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_650), .A2(n_542), .B1(n_532), .B2(n_531), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_625), .A2(n_597), .B1(n_542), .B2(n_532), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_686), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_611), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_621), .A2(n_532), .B1(n_531), .B2(n_598), .Y(n_716) );
OR2x2_ASAP7_75t_L g717 ( .A(n_650), .B(n_531), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_611), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_675), .A2(n_532), .B1(n_531), .B2(n_598), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_681), .Y(n_720) );
BUFx8_ASAP7_75t_L g721 ( .A(n_680), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_695), .A2(n_671), .B1(n_614), .B2(n_616), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_601), .A2(n_542), .B1(n_597), .B2(n_593), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_600), .B(n_589), .Y(n_724) );
INVxp67_ASAP7_75t_SL g725 ( .A(n_612), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_648), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_603), .B(n_589), .Y(n_727) );
OA21x2_ASAP7_75t_L g728 ( .A1(n_629), .A2(n_386), .B(n_376), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_695), .A2(n_542), .B1(n_592), .B2(n_597), .Y(n_729) );
AOI222xp33_ASAP7_75t_L g730 ( .A1(n_656), .A2(n_347), .B1(n_294), .B2(n_298), .C1(n_300), .C2(n_345), .Y(n_730) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_685), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_602), .A2(n_518), .B1(n_528), .B2(n_517), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_668), .A2(n_318), .B1(n_342), .B2(n_346), .C(n_351), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_661), .A2(n_517), .B1(n_518), .B2(n_528), .C(n_529), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_623), .A2(n_541), .B1(n_529), .B2(n_590), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_637), .A2(n_353), .B1(n_341), .B2(n_335), .C(n_334), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_654), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_612), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_644), .B(n_541), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g740 ( .A1(n_683), .A2(n_316), .B(n_321), .C(n_313), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_663), .A2(n_328), .B1(n_400), .B2(n_401), .C(n_301), .Y(n_741) );
AO31x2_ASAP7_75t_L g742 ( .A1(n_615), .A2(n_386), .A3(n_395), .B(n_376), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_669), .B(n_558), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_672), .B(n_679), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_687), .A2(n_401), .B1(n_400), .B2(n_281), .C(n_301), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_622), .A2(n_582), .B1(n_558), .B2(n_599), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_680), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_626), .A2(n_590), .B1(n_582), .B2(n_400), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_649), .A2(n_582), .B1(n_558), .B2(n_599), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_632), .A2(n_582), .B1(n_401), .B2(n_317), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_638), .B(n_558), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_615), .A2(n_636), .B(n_631), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_674), .A2(n_582), .B1(n_401), .B2(n_599), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_631), .A2(n_582), .B1(n_599), .B2(n_303), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_636), .A2(n_246), .B1(n_319), .B2(n_303), .Y(n_755) );
AO21x2_ASAP7_75t_L g756 ( .A1(n_684), .A2(n_386), .B(n_376), .Y(n_756) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_646), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g758 ( .A1(n_640), .A2(n_395), .B(n_389), .C(n_401), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_639), .A2(n_401), .B1(n_395), .B2(n_389), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_670), .B(n_6), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_639), .A2(n_389), .B1(n_392), .B2(n_393), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g762 ( .A1(n_619), .A2(n_389), .B1(n_497), .B2(n_489), .C(n_508), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_645), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_645), .A2(n_389), .B1(n_392), .B2(n_393), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_647), .B(n_6), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_608), .B(n_7), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_627), .A2(n_393), .B1(n_392), .B2(n_508), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_651), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_651), .A2(n_393), .B(n_508), .C(n_435), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_690), .A2(n_508), .B1(n_393), .B2(n_435), .C(n_439), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_617), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_689), .A2(n_393), .B1(n_439), .B2(n_435), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_694), .B(n_439), .C(n_435), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_660), .A2(n_439), .B1(n_9), .B2(n_10), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_657), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_659), .B(n_8), .Y(n_776) );
OA21x2_ASAP7_75t_L g777 ( .A1(n_659), .A2(n_439), .B(n_88), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_681), .A2(n_8), .B1(n_9), .B2(n_11), .C(n_12), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_666), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_605), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_666), .B(n_13), .Y(n_781) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_685), .B(n_14), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_608), .B(n_15), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_709), .A2(n_658), .B1(n_655), .B2(n_628), .C(n_634), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_726), .Y(n_785) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_717), .Y(n_786) );
OAI33xp33_ASAP7_75t_L g787 ( .A1(n_755), .A2(n_676), .A3(n_678), .B1(n_682), .B2(n_19), .B3(n_20), .Y(n_787) );
NOR3xp33_ASAP7_75t_L g788 ( .A(n_778), .B(n_677), .C(n_624), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_730), .B(n_677), .C(n_624), .Y(n_789) );
AOI221xp5_ASAP7_75t_L g790 ( .A1(n_698), .A2(n_676), .B1(n_635), .B2(n_643), .C(n_664), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_760), .B(n_635), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_715), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_696), .A2(n_646), .B1(n_691), .B2(n_630), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_702), .B(n_617), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_737), .Y(n_795) );
NAND4xp25_ASAP7_75t_L g796 ( .A(n_733), .B(n_642), .C(n_652), .D(n_692), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_779), .A2(n_692), .B(n_688), .C(n_685), .Y(n_797) );
BUFx3_ASAP7_75t_L g798 ( .A(n_780), .Y(n_798) );
AOI222xp33_ASAP7_75t_L g799 ( .A1(n_699), .A2(n_643), .B1(n_630), .B2(n_685), .C1(n_688), .C2(n_21), .Y(n_799) );
OR2x6_ASAP7_75t_L g800 ( .A(n_766), .B(n_646), .Y(n_800) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_725), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g802 ( .A1(n_736), .A2(n_688), .B1(n_685), .B2(n_691), .C(n_617), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_718), .Y(n_803) );
OAI222xp33_ASAP7_75t_L g804 ( .A1(n_712), .A2(n_722), .B1(n_711), .B2(n_782), .C1(n_783), .C2(n_766), .Y(n_804) );
BUFx3_ASAP7_75t_L g805 ( .A(n_743), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_721), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_738), .Y(n_807) );
AND2x4_ASAP7_75t_L g808 ( .A(n_743), .B(n_688), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_725), .A2(n_688), .B(n_646), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_740), .B(n_617), .C(n_16), .Y(n_810) );
OR2x2_ASAP7_75t_L g811 ( .A(n_739), .B(n_617), .Y(n_811) );
OAI33xp33_ASAP7_75t_L g812 ( .A1(n_771), .A2(n_16), .A3(n_17), .B1(n_20), .B2(n_22), .B3(n_23), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_711), .A2(n_17), .B(n_23), .Y(n_813) );
OAI221xp5_ASAP7_75t_SL g814 ( .A1(n_722), .A2(n_24), .B1(n_25), .B2(n_26), .C(n_27), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_701), .B(n_29), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_721), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_816) );
BUFx3_ASAP7_75t_L g817 ( .A(n_707), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_747), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_818) );
OR2x2_ASAP7_75t_L g819 ( .A(n_744), .B(n_32), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_763), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_745), .B(n_34), .C(n_35), .Y(n_821) );
INVx4_ASAP7_75t_SL g822 ( .A(n_713), .Y(n_822) );
OA222x2_ASAP7_75t_L g823 ( .A1(n_724), .A2(n_40), .B1(n_41), .B2(n_42), .C1(n_44), .C2(n_45), .Y(n_823) );
AO21x2_ASAP7_75t_L g824 ( .A1(n_769), .A2(n_41), .B(n_46), .Y(n_824) );
OAI211xp5_ASAP7_75t_SL g825 ( .A1(n_727), .A2(n_46), .B(n_47), .C(n_49), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_708), .Y(n_826) );
OR2x6_ASAP7_75t_L g827 ( .A(n_783), .B(n_782), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_710), .B(n_47), .Y(n_828) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_729), .A2(n_51), .B1(n_53), .B2(n_54), .C(n_56), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_768), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_714), .B(n_58), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_781), .Y(n_832) );
INVx4_ASAP7_75t_L g833 ( .A(n_707), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_775), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_776), .B(n_62), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_774), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_731), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g838 ( .A1(n_729), .A2(n_68), .B1(n_69), .B2(n_70), .C(n_71), .Y(n_838) );
AND2x4_ASAP7_75t_L g839 ( .A(n_757), .B(n_91), .Y(n_839) );
OAI211xp5_ASAP7_75t_L g840 ( .A1(n_699), .A2(n_68), .B(n_69), .C(n_70), .Y(n_840) );
OAI211xp5_ASAP7_75t_L g841 ( .A1(n_753), .A2(n_73), .B(n_74), .C(n_75), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_753), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_703), .A2(n_80), .B1(n_81), .B2(n_82), .Y(n_843) );
OAI33xp33_ASAP7_75t_L g844 ( .A1(n_765), .A2(n_83), .A3(n_84), .B1(n_85), .B2(n_86), .B3(n_87), .Y(n_844) );
OAI222xp33_ASAP7_75t_L g845 ( .A1(n_720), .A2(n_83), .B1(n_85), .B2(n_87), .C1(n_92), .C2(n_93), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_700), .A2(n_95), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_732), .A2(n_101), .B1(n_109), .B2(n_114), .Y(n_847) );
AOI211xp5_ASAP7_75t_L g848 ( .A1(n_734), .A2(n_115), .B(n_116), .C(n_118), .Y(n_848) );
OAI322xp33_ASAP7_75t_L g849 ( .A1(n_751), .A2(n_119), .A3(n_120), .B1(n_123), .B2(n_125), .C1(n_129), .C2(n_130), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_732), .A2(n_132), .B1(n_133), .B2(n_135), .Y(n_850) );
OAI31xp33_ASAP7_75t_L g851 ( .A1(n_716), .A2(n_136), .A3(n_137), .B(n_138), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_742), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_704), .A2(n_723), .B1(n_741), .B2(n_697), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_735), .A2(n_142), .B1(n_143), .B2(n_144), .C(n_146), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_749), .A2(n_148), .B1(n_149), .B2(n_152), .Y(n_855) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_750), .A2(n_153), .B1(n_154), .B2(n_156), .C(n_158), .Y(n_856) );
OAI31xp33_ASAP7_75t_L g857 ( .A1(n_758), .A2(n_160), .A3(n_162), .B(n_165), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_750), .A2(n_168), .B1(n_169), .B2(n_170), .C(n_171), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_731), .Y(n_859) );
OAI33xp33_ASAP7_75t_L g860 ( .A1(n_759), .A2(n_173), .A3(n_174), .B1(n_175), .B2(n_178), .B3(n_179), .Y(n_860) );
AOI211xp5_ASAP7_75t_L g861 ( .A1(n_719), .A2(n_180), .B(n_181), .C(n_182), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g862 ( .A1(n_752), .A2(n_187), .B1(n_188), .B2(n_191), .Y(n_862) );
BUFx2_ASAP7_75t_L g863 ( .A(n_731), .Y(n_863) );
AND2x2_ASAP7_75t_L g864 ( .A(n_706), .B(n_192), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_794), .A2(n_756), .B1(n_762), .B2(n_748), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_785), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_786), .B(n_731), .Y(n_867) );
INVxp67_ASAP7_75t_L g868 ( .A(n_806), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_826), .B(n_742), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_795), .Y(n_870) );
OAI31xp33_ASAP7_75t_L g871 ( .A1(n_840), .A2(n_764), .A3(n_761), .B(n_759), .Y(n_871) );
BUFx3_ASAP7_75t_L g872 ( .A(n_805), .Y(n_872) );
AND2x2_ASAP7_75t_SL g873 ( .A(n_839), .B(n_777), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_799), .A2(n_748), .B1(n_746), .B2(n_754), .Y(n_874) );
INVx4_ASAP7_75t_L g875 ( .A(n_800), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_823), .B(n_756), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_828), .B(n_767), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g878 ( .A(n_816), .B(n_767), .C(n_769), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_825), .A2(n_705), .B1(n_770), .B2(n_773), .Y(n_879) );
OR2x2_ASAP7_75t_L g880 ( .A(n_811), .B(n_728), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_808), .B(n_194), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_792), .B(n_728), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_792), .Y(n_883) );
AND2x4_ASAP7_75t_L g884 ( .A(n_808), .B(n_195), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_803), .B(n_807), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_803), .B(n_728), .Y(n_886) );
INVx2_ASAP7_75t_SL g887 ( .A(n_817), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_810), .A2(n_777), .B1(n_772), .B2(n_209), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_835), .B(n_206), .Y(n_889) );
NAND2xp5_ASAP7_75t_SL g890 ( .A(n_802), .B(n_208), .Y(n_890) );
BUFx3_ASAP7_75t_L g891 ( .A(n_817), .Y(n_891) );
INVx3_ASAP7_75t_SL g892 ( .A(n_798), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_832), .B(n_244), .Y(n_893) );
OR2x6_ASAP7_75t_L g894 ( .A(n_800), .B(n_216), .Y(n_894) );
NAND3xp33_ASAP7_75t_L g895 ( .A(n_814), .B(n_222), .C(n_224), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_819), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_815), .Y(n_897) );
AOI33xp33_ASAP7_75t_L g898 ( .A1(n_818), .A2(n_225), .A3(n_226), .B1(n_227), .B2(n_228), .B3(n_230), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_807), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_833), .B(n_231), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_820), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_820), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_830), .Y(n_903) );
OAI31xp33_ASAP7_75t_L g904 ( .A1(n_845), .A2(n_233), .A3(n_234), .B(n_235), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_830), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_834), .Y(n_906) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_801), .Y(n_907) );
INVx2_ASAP7_75t_L g908 ( .A(n_834), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_800), .B(n_808), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_831), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_839), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_790), .B(n_843), .Y(n_912) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_836), .A2(n_827), .B1(n_789), .B2(n_829), .Y(n_913) );
OAI33xp33_ASAP7_75t_L g914 ( .A1(n_862), .A2(n_793), .A3(n_850), .B1(n_847), .B2(n_821), .B3(n_852), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_837), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_837), .B(n_859), .Y(n_916) );
INVx3_ASAP7_75t_L g917 ( .A(n_827), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_841), .B(n_788), .C(n_838), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_859), .B(n_863), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_827), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_812), .A2(n_844), .B1(n_787), .B2(n_842), .Y(n_921) );
INVx5_ASAP7_75t_SL g922 ( .A(n_839), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_813), .Y(n_923) );
INVx1_ASAP7_75t_SL g924 ( .A(n_822), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_809), .B(n_813), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_824), .Y(n_926) );
INVx3_ASAP7_75t_L g927 ( .A(n_864), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_804), .A2(n_849), .B1(n_784), .B2(n_862), .C(n_860), .Y(n_928) );
INVxp67_ASAP7_75t_L g929 ( .A(n_824), .Y(n_929) );
AND2x4_ASAP7_75t_L g930 ( .A(n_822), .B(n_864), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_822), .Y(n_931) );
NAND4xp25_ASAP7_75t_L g932 ( .A(n_848), .B(n_853), .C(n_796), .D(n_861), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_853), .A2(n_854), .B1(n_858), .B2(n_851), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_797), .B(n_855), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_856), .B(n_857), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_846), .B(n_791), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_785), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_826), .B(n_771), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_866), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_870), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_938), .B(n_869), .Y(n_941) );
OAI33xp33_ASAP7_75t_L g942 ( .A1(n_896), .A2(n_868), .A3(n_913), .B1(n_937), .B2(n_897), .B3(n_910), .Y(n_942) );
AND3x2_ASAP7_75t_L g943 ( .A(n_876), .B(n_931), .C(n_930), .Y(n_943) );
INVx2_ASAP7_75t_SL g944 ( .A(n_907), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_869), .B(n_885), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_916), .B(n_927), .Y(n_946) );
INVx1_ASAP7_75t_SL g947 ( .A(n_892), .Y(n_947) );
OAI21xp5_ASAP7_75t_L g948 ( .A1(n_918), .A2(n_895), .B(n_921), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_899), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g950 ( .A1(n_922), .A2(n_912), .B1(n_936), .B2(n_894), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_901), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_922), .B(n_880), .Y(n_952) );
NOR2x1_ASAP7_75t_L g953 ( .A(n_894), .B(n_924), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_902), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_916), .B(n_927), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_927), .B(n_915), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_915), .B(n_883), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_883), .B(n_905), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_905), .B(n_906), .Y(n_959) );
BUFx2_ASAP7_75t_L g960 ( .A(n_891), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_903), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_914), .A2(n_875), .B1(n_930), .B2(n_877), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_887), .B(n_922), .Y(n_963) );
OR2x2_ASAP7_75t_L g964 ( .A(n_908), .B(n_867), .Y(n_964) );
OAI21xp5_ASAP7_75t_L g965 ( .A1(n_921), .A2(n_878), .B(n_904), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_926), .B(n_919), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_911), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_919), .Y(n_968) );
AND2x4_ASAP7_75t_L g969 ( .A(n_875), .B(n_930), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_872), .B(n_892), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_923), .Y(n_971) );
OR2x2_ASAP7_75t_L g972 ( .A(n_925), .B(n_909), .Y(n_972) );
AO21x1_ASAP7_75t_L g973 ( .A1(n_875), .A2(n_890), .B(n_926), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_929), .B(n_886), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_917), .B(n_920), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_882), .B(n_886), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_917), .Y(n_977) );
INVx2_ASAP7_75t_L g978 ( .A(n_882), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_917), .B(n_920), .Y(n_979) );
BUFx3_ASAP7_75t_L g980 ( .A(n_881), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_873), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_873), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_889), .B(n_893), .Y(n_983) );
NAND4xp25_ASAP7_75t_L g984 ( .A(n_928), .B(n_933), .C(n_865), .D(n_934), .Y(n_984) );
OAI21xp5_ASAP7_75t_L g985 ( .A1(n_933), .A2(n_898), .B(n_890), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_934), .B(n_865), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_881), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_881), .B(n_884), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_900), .B(n_884), .Y(n_989) );
NAND4xp25_ASAP7_75t_L g990 ( .A(n_888), .B(n_874), .C(n_898), .D(n_935), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_884), .Y(n_991) );
AND2x4_ASAP7_75t_L g992 ( .A(n_888), .B(n_879), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_879), .B(n_871), .Y(n_993) );
NAND4xp25_ASAP7_75t_L g994 ( .A(n_876), .B(n_607), .C(n_816), .D(n_932), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_951), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_944), .Y(n_996) );
INVx3_ASAP7_75t_L g997 ( .A(n_969), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_939), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_940), .Y(n_999) );
XOR2xp5_ASAP7_75t_L g1000 ( .A(n_994), .B(n_984), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_951), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_954), .Y(n_1002) );
NOR3xp33_ASAP7_75t_L g1003 ( .A(n_948), .B(n_965), .C(n_942), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_971), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_978), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_941), .B(n_945), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_949), .Y(n_1007) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_960), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_961), .Y(n_1009) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_969), .B(n_955), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_945), .B(n_986), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_957), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_944), .B(n_968), .Y(n_1013) );
INVx1_ASAP7_75t_SL g1014 ( .A(n_947), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_970), .Y(n_1015) );
OAI21x1_ASAP7_75t_SL g1016 ( .A1(n_953), .A2(n_973), .B(n_989), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_976), .B(n_946), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_976), .B(n_946), .Y(n_1018) );
NOR3xp33_ASAP7_75t_L g1019 ( .A(n_990), .B(n_985), .C(n_993), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_967), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_964), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_958), .Y(n_1022) );
AOI32xp33_ASAP7_75t_L g1023 ( .A1(n_988), .A2(n_962), .A3(n_969), .B1(n_980), .B2(n_992), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_950), .A2(n_993), .B1(n_988), .B2(n_991), .Y(n_1024) );
XOR2xp5_ASAP7_75t_L g1025 ( .A(n_972), .B(n_952), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_972), .B(n_964), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_966), .B(n_956), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_957), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_1000), .B(n_943), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1006), .B(n_982), .Y(n_1030) );
AND2x4_ASAP7_75t_SL g1031 ( .A(n_1010), .B(n_979), .Y(n_1031) );
NAND2xp5_ASAP7_75t_SL g1032 ( .A(n_1016), .B(n_973), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_1019), .A2(n_983), .B1(n_992), .B2(n_987), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_995), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1011), .B(n_974), .Y(n_1035) );
OAI211xp5_ASAP7_75t_L g1036 ( .A1(n_1000), .A2(n_1003), .B(n_1023), .C(n_1024), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_995), .Y(n_1037) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_1014), .B(n_963), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1006), .B(n_974), .Y(n_1039) );
OAI22x1_ASAP7_75t_L g1040 ( .A1(n_1025), .A2(n_982), .B1(n_981), .B2(n_952), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1021), .B(n_959), .Y(n_1041) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_1008), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1001), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_1025), .A2(n_975), .B1(n_981), .B2(n_979), .Y(n_1044) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_997), .B(n_977), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1002), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1026), .Y(n_1047) );
NOR2xp67_ASAP7_75t_SL g1048 ( .A(n_1008), .B(n_996), .Y(n_1048) );
XNOR2xp5_ASAP7_75t_L g1049 ( .A(n_1010), .B(n_1015), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1026), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_998), .Y(n_1051) );
XOR2x2_ASAP7_75t_L g1052 ( .A(n_1017), .B(n_1018), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1027), .B(n_1012), .Y(n_1053) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_1005), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_1013), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_999), .Y(n_1056) );
XOR2x2_ASAP7_75t_SL g1057 ( .A(n_1016), .B(n_1020), .Y(n_1057) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_1028), .B(n_1022), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_1022), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_1004), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1007), .Y(n_1061) );
CKINVDCx16_ASAP7_75t_R g1062 ( .A(n_1055), .Y(n_1062) );
NOR2xp33_ASAP7_75t_L g1063 ( .A(n_1029), .B(n_1036), .Y(n_1063) );
AOI321xp33_ASAP7_75t_L g1064 ( .A1(n_1033), .A2(n_1044), .A3(n_1032), .B1(n_1038), .B2(n_1047), .C(n_1050), .Y(n_1064) );
INVx2_ASAP7_75t_SL g1065 ( .A(n_1049), .Y(n_1065) );
AOI21xp33_ASAP7_75t_L g1066 ( .A1(n_1040), .A2(n_1056), .B(n_1051), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1030), .Y(n_1067) );
NAND3xp33_ASAP7_75t_SL g1068 ( .A(n_1057), .B(n_1055), .C(n_1059), .Y(n_1068) );
AOI21xp5_ASAP7_75t_L g1069 ( .A1(n_1040), .A2(n_1052), .B(n_1031), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1030), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1067), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_1070), .B(n_1041), .Y(n_1072) );
AOI221xp5_ASAP7_75t_L g1073 ( .A1(n_1063), .A2(n_1059), .B1(n_1048), .B2(n_1058), .C(n_1042), .Y(n_1073) );
O2A1O1Ixp33_ASAP7_75t_L g1074 ( .A1(n_1068), .A2(n_1042), .B(n_1035), .C(n_1054), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1065), .Y(n_1075) );
OAI221xp5_ASAP7_75t_L g1076 ( .A1(n_1064), .A2(n_1048), .B1(n_1054), .B2(n_1039), .C(n_1061), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1075), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_1076), .A2(n_1069), .B1(n_1066), .B2(n_1062), .Y(n_1078) );
NOR3xp33_ASAP7_75t_L g1079 ( .A(n_1076), .B(n_1009), .C(n_1007), .Y(n_1079) );
XOR2x2_ASAP7_75t_L g1080 ( .A(n_1073), .B(n_1053), .Y(n_1080) );
NAND3xp33_ASAP7_75t_SL g1081 ( .A(n_1078), .B(n_1074), .C(n_1071), .Y(n_1081) );
HB1xp67_ASAP7_75t_L g1082 ( .A(n_1077), .Y(n_1082) );
O2A1O1Ixp33_ASAP7_75t_L g1083 ( .A1(n_1081), .A2(n_1079), .B(n_1080), .C(n_1072), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1082), .Y(n_1084) );
XOR2xp5_ASAP7_75t_L g1085 ( .A(n_1084), .B(n_1045), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1083), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1087 ( .A1(n_1086), .A2(n_1043), .B1(n_1046), .B2(n_1034), .C(n_1037), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_1085), .A2(n_1060), .B1(n_1043), .B2(n_1034), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1088), .Y(n_1089) );
AOI21xp5_ASAP7_75t_L g1090 ( .A1(n_1089), .A2(n_1087), .B(n_1060), .Y(n_1090) );
endmodule