module fake_jpeg_2027_n_80 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_1),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_30),
.B1(n_24),
.B2(n_26),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_45),
.B1(n_28),
.B2(n_34),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_2),
.C(n_3),
.Y(n_52)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_30),
.B1(n_24),
.B2(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_39),
.B1(n_43),
.B2(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_57),
.B1(n_7),
.B2(n_8),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_5),
.B(n_6),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_18),
.Y(n_64)
);

XNOR2x2_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_6),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_68),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_66),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_13),
.C(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_67),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_22),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_70),
.B1(n_63),
.B2(n_55),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_71),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_58),
.B(n_59),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_20),
.Y(n_80)
);


endmodule