module fake_jpeg_28069_n_202 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_25),
.Y(n_35)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_37)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_37),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_22),
.B1(n_25),
.B2(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_29),
.B1(n_26),
.B2(n_14),
.Y(n_71)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_22),
.B1(n_20),
.B2(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_55),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_28),
.B(n_30),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_30),
.B(n_28),
.C(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_31),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_53),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_27),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_24),
.B(n_19),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_46),
.B1(n_48),
.B2(n_29),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_31),
.B1(n_38),
.B2(n_19),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_85),
.B1(n_65),
.B2(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_79),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_44),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_40),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_40),
.B1(n_52),
.B2(n_26),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_82),
.B1(n_73),
.B2(n_62),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_26),
.B1(n_29),
.B2(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_88),
.B(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_12),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_24),
.C(n_12),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_67),
.C(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_106),
.B1(n_111),
.B2(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_105),
.B(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_104),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_58),
.B1(n_65),
.B2(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_24),
.B1(n_19),
.B2(n_12),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_24),
.C(n_10),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

XOR2x2_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_11),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_11),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_81),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_97),
.B(n_94),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_124),
.B(n_138),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_126),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_77),
.B1(n_10),
.B2(n_11),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_18),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_18),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_133),
.B(n_95),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_135),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_115),
.A2(n_10),
.B1(n_9),
.B2(n_7),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_110),
.B1(n_95),
.B2(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_100),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_149),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_112),
.C(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_145),
.C(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_117),
.C(n_98),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_153),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_120),
.B1(n_139),
.B2(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_159),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_123),
.C(n_118),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_145),
.C(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_132),
.B1(n_133),
.B2(n_131),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_144),
.B1(n_143),
.B2(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_169),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_R g169 ( 
.A(n_162),
.B(n_133),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_132),
.B1(n_149),
.B2(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_157),
.C(n_156),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_2),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_179),
.C(n_182),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_143),
.B(n_166),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_175),
.B(n_5),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_158),
.C(n_164),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_9),
.C(n_3),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_170),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_5),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_6),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_189),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_184),
.B1(n_185),
.B2(n_6),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_6),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_191),
.C(n_193),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_195),
.Y(n_202)
);


endmodule