module fake_jpeg_1838_n_228 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_228);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_0),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_61),
.B1(n_62),
.B2(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_95),
.B1(n_100),
.B2(n_85),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_62),
.B1(n_68),
.B2(n_78),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_54),
.B1(n_79),
.B2(n_66),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_103),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_81),
.B1(n_86),
.B2(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_118),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_83),
.B1(n_84),
.B2(n_74),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_63),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_76),
.B1(n_73),
.B2(n_82),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_92),
.A2(n_76),
.B1(n_65),
.B2(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_46),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_67),
.B1(n_56),
.B2(n_60),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_70),
.B1(n_75),
.B2(n_71),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_119),
.B1(n_77),
.B2(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_77),
.B1(n_71),
.B2(n_72),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_72),
.B1(n_63),
.B2(n_58),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_63),
.B(n_58),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_6),
.B(n_7),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_51),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_104),
.C(n_110),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_139),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_130),
.B(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_58),
.B(n_1),
.Y(n_130)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_44),
.C(n_42),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_3),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_121),
.B(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_141),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_162),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2x1_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_10),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_9),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_125),
.B(n_128),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_174),
.B(n_182),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_177),
.B(n_178),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_9),
.B(n_10),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_36),
.C(n_32),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_181),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_31),
.B(n_27),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_26),
.C(n_25),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_24),
.B(n_22),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_184),
.B(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_11),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_165),
.B(n_149),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_179),
.B(n_174),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_163),
.B1(n_157),
.B2(n_144),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_194),
.B1(n_147),
.B2(n_157),
.Y(n_206)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_196),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_144),
.B1(n_163),
.B2(n_173),
.Y(n_194)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_197),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_183),
.B1(n_147),
.B2(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_186),
.B1(n_182),
.B2(n_13),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_181),
.C(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_208),
.C(n_175),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_178),
.B(n_172),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_200),
.A2(n_195),
.B(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_163),
.B1(n_171),
.B2(n_187),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_214),
.B1(n_11),
.B2(n_12),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_185),
.B1(n_177),
.B2(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_207),
.B1(n_210),
.B2(n_209),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_220),
.B(n_218),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_221),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

AOI321xp33_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_219),
.A3(n_211),
.B1(n_18),
.B2(n_20),
.C(n_21),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_15),
.CI(n_16),
.CON(n_227),
.SN(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_219),
.Y(n_228)
);


endmodule