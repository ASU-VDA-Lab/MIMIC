module fake_jpeg_13531_n_347 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_50),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_19),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_39),
.B1(n_38),
.B2(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_30),
.B1(n_28),
.B2(n_31),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_60),
.A2(n_75),
.B1(n_90),
.B2(n_93),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_30),
.B(n_28),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_37),
.B(n_50),
.Y(n_106)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_85),
.Y(n_104)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_32),
.B1(n_24),
.B2(n_33),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_22),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_39),
.B1(n_38),
.B2(n_35),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_93),
.B1(n_75),
.B2(n_60),
.Y(n_97)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_22),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_39),
.B1(n_38),
.B2(n_32),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.C(n_37),
.Y(n_103)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_35),
.B1(n_39),
.B2(n_38),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_30),
.C(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_103),
.B1(n_126),
.B2(n_45),
.Y(n_149)
);

NOR2x1_ASAP7_75t_R g101 ( 
.A(n_67),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_46),
.B1(n_55),
.B2(n_31),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_111),
.B1(n_123),
.B2(n_44),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_112),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_65),
.B(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_118),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_31),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_57),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_66),
.B(n_25),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_25),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_122),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_78),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_132),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_52),
.B1(n_36),
.B2(n_35),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_73),
.B1(n_50),
.B2(n_81),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_90),
.A2(n_53),
.B1(n_45),
.B2(n_44),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_12),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_9),
.Y(n_167)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_53),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_88),
.C(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_50),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_1),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_153),
.B1(n_158),
.B2(n_1),
.Y(n_191)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_99),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_108),
.B1(n_115),
.B2(n_117),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_130),
.C(n_108),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_89),
.C(n_84),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_147),
.C(n_132),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_73),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_133),
.B1(n_118),
.B2(n_106),
.Y(n_172)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_45),
.B1(n_53),
.B2(n_74),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_88),
.B1(n_89),
.B2(n_84),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_162),
.B1(n_163),
.B2(n_131),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_107),
.B1(n_111),
.B2(n_104),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_35),
.B1(n_73),
.B2(n_2),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_12),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_178),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_174),
.B1(n_176),
.B2(n_186),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_98),
.B1(n_101),
.B2(n_100),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_164),
.A2(n_129),
.B1(n_131),
.B2(n_109),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_191),
.B1(n_4),
.B2(n_5),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_184),
.C(n_198),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_130),
.B1(n_99),
.B2(n_115),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_182),
.B(n_190),
.Y(n_221)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_117),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_145),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_197),
.B1(n_200),
.B2(n_136),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_196),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_8),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_16),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_9),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_7),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_138),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_151),
.A2(n_10),
.B1(n_13),
.B2(n_16),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_2),
.B(n_3),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_134),
.B(n_135),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_10),
.C(n_13),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_169),
.C(n_163),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_220),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_153),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_225),
.B(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_144),
.C(n_139),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_229),
.C(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_194),
.B(n_134),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_146),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_135),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_227),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_159),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_162),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_150),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_176),
.B(n_148),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_148),
.B1(n_136),
.B2(n_156),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_16),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_3),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_226),
.B1(n_227),
.B2(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_244),
.B1(n_231),
.B2(n_230),
.Y(n_269)
);

A2O1A1O1Ixp25_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_182),
.B(n_178),
.C(n_181),
.D(n_201),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_208),
.B(n_211),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_190),
.B(n_185),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_253),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_252),
.C(n_256),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_210),
.A2(n_186),
.B1(n_171),
.B2(n_175),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_171),
.C(n_193),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_218),
.B(n_211),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_211),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_200),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_206),
.C(n_215),
.Y(n_266)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_259),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_266),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_216),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_268),
.B(n_235),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_276),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_212),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_272),
.C(n_277),
.Y(n_286)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_217),
.C(n_193),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

XOR2x2_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_197),
.Y(n_275)
);

NOR3xp33_ASAP7_75t_SL g276 ( 
.A(n_240),
.B(n_230),
.C(n_183),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_183),
.C(n_173),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_205),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_278),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_173),
.B1(n_179),
.B2(n_192),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_269),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_291),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_256),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_235),
.CI(n_253),
.CON(n_293),
.SN(n_293)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_238),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_251),
.C(n_237),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_277),
.C(n_270),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_260),
.B1(n_251),
.B2(n_237),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_306),
.B1(n_293),
.B2(n_284),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_260),
.B(n_276),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_301),
.B(n_310),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_265),
.C(n_275),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_242),
.B(n_249),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_305),
.B(n_299),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_258),
.B1(n_246),
.B2(n_249),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_295),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_250),
.C(n_245),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_241),
.B1(n_246),
.B2(n_192),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_283),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_291),
.C(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_317),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_290),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_301),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_309),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_307),
.B1(n_303),
.B2(n_293),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_313),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_327),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_330),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_302),
.C(n_298),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_292),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_315),
.C(n_282),
.Y(n_332)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_315),
.B1(n_318),
.B2(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_335),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_324),
.A2(n_288),
.B1(n_294),
.B2(n_319),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_326),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_337),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_337),
.B(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_341),
.B(n_342),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_336),
.B1(n_339),
.B2(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_329),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_288),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_4),
.Y(n_347)
);


endmodule