module fake_jpeg_25145_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_42),
.Y(n_81)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_70),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_49),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_61),
.B1(n_50),
.B2(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_43),
.B1(n_55),
.B2(n_54),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_82),
.Y(n_85)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_58),
.Y(n_89)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_76),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_52),
.C(n_53),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_5),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_59),
.B1(n_57),
.B2(n_49),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_92),
.B1(n_98),
.B2(n_4),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_74),
.A2(n_57),
.B1(n_59),
.B2(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_73),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_104),
.A2(n_108),
.B(n_6),
.Y(n_116)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_27),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_112),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_92),
.B1(n_90),
.B2(n_86),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_113),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_121),
.B1(n_100),
.B2(n_117),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_99),
.A3(n_8),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_18),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_32),
.C(n_19),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_107),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_7),
.B(n_21),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.C(n_119),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_22),
.C(n_23),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_129),
.B1(n_121),
.B2(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_130),
.B(n_123),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_124),
.B(n_29),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_28),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_30),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_35),
.B(n_37),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_38),
.Y(n_136)
);


endmodule