module fake_jpeg_773_n_187 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_11),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_0),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_63),
.B1(n_48),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_48),
.B1(n_63),
.B2(n_61),
.Y(n_93)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_82),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_95),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_63),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_52),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_62),
.C(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_103),
.Y(n_108)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_55),
.B1(n_52),
.B2(n_60),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_53),
.B1(n_58),
.B2(n_75),
.Y(n_118)
);

NAND2x1_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_58),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_74),
.B(n_47),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_116),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_61),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_93),
.B1(n_86),
.B2(n_85),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_118),
.B1(n_18),
.B2(n_42),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_53),
.B(n_47),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_19),
.B1(n_45),
.B2(n_44),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_91),
.B1(n_94),
.B2(n_3),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_111),
.B1(n_105),
.B2(n_121),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_11),
.B(n_12),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_20),
.C(n_43),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_25),
.C(n_35),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_134),
.B1(n_141),
.B2(n_143),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_153),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_130),
.B(n_121),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_125),
.B(n_8),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_10),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_143),
.B1(n_134),
.B2(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_168),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_130),
.B1(n_142),
.B2(n_123),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_145),
.B1(n_152),
.B2(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_27),
.C(n_34),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_15),
.C(n_29),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_147),
.B1(n_159),
.B2(n_14),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_12),
.B1(n_13),
.B2(n_155),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_163),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_163),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_180),
.B(n_177),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_170),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_167),
.B(n_176),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_169),
.B(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_165),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_33),
.Y(n_187)
);


endmodule