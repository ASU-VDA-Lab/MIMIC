module fake_jpeg_3680_n_300 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_6),
.B(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_33),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_62),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_26),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_17),
.A2(n_15),
.B(n_14),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_41),
.C(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_67),
.Y(n_94)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_11),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_46),
.B(n_28),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_71),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_30),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_35),
.B1(n_40),
.B2(n_38),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_80),
.B(n_91),
.Y(n_133)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_43),
.B1(n_34),
.B2(n_29),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_104),
.B1(n_11),
.B2(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_40),
.B1(n_28),
.B2(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_103),
.B1(n_40),
.B2(n_32),
.Y(n_116)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_50),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_96),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_22),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_25),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_35),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_57),
.A2(n_40),
.B1(n_28),
.B2(n_36),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_43),
.B1(n_29),
.B2(n_32),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_48),
.B(n_26),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_52),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_107),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_48),
.B(n_30),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_79),
.C(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_115),
.B(n_124),
.C(n_128),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_129),
.B1(n_134),
.B2(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_40),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_130),
.B1(n_132),
.B2(n_139),
.Y(n_149)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_38),
.B(n_23),
.C(n_12),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_127),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_76),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_76),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_78),
.A2(n_38),
.B1(n_23),
.B2(n_12),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_77),
.A2(n_10),
.B1(n_9),
.B2(n_2),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_147),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_97),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_92),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_139)
);

INVx2_ASAP7_75t_R g141 ( 
.A(n_70),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_142),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_86),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_109),
.B1(n_81),
.B2(n_83),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_95),
.A2(n_109),
.B1(n_108),
.B2(n_90),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_102),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_74),
.Y(n_147)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_146),
.Y(n_201)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_108),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_97),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_175),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_177),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_129),
.B1(n_121),
.B2(n_135),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_81),
.B1(n_83),
.B2(n_89),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_89),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_172),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_70),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_102),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_180),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_110),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_110),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_119),
.B(n_133),
.C(n_115),
.D(n_140),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_186),
.B(n_207),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_119),
.B(n_115),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_133),
.C(n_126),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_198),
.C(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_120),
.B1(n_140),
.B2(n_134),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_120),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_163),
.C(n_156),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_124),
.B(n_114),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_199),
.A2(n_197),
.B(n_201),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_155),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_143),
.C(n_117),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_132),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_206),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_168),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_155),
.A2(n_127),
.B1(n_128),
.B2(n_141),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_169),
.B(n_149),
.C(n_177),
.D(n_160),
.Y(n_208)
);

AOI221xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_149),
.B1(n_160),
.B2(n_167),
.C(n_157),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_160),
.A2(n_141),
.B(n_148),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_153),
.B(n_180),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_148),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_212),
.C(n_150),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_152),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_111),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_157),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_214),
.B(n_219),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_216),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_150),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_229),
.C(n_236),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_152),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_227),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_225),
.B(n_226),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_230),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_206),
.B(n_209),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_162),
.B(n_165),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_173),
.C(n_174),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_151),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_151),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_238),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_164),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_164),
.C(n_111),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_183),
.A2(n_111),
.B(n_185),
.C(n_204),
.D(n_205),
.Y(n_237)
);

OA21x2_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_189),
.B(n_196),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_111),
.C(n_210),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_205),
.B(n_208),
.C(n_189),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_242),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_240),
.C(n_255),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_188),
.B1(n_202),
.B2(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_188),
.A3(n_190),
.B1(n_194),
.B2(n_223),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_235),
.B1(n_231),
.B2(n_223),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_220),
.B1(n_238),
.B2(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_214),
.A2(n_230),
.B1(n_219),
.B2(n_218),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_217),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_217),
.C(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_264),
.C(n_266),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_264),
.Y(n_280)
);

AOI321xp33_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_228),
.A3(n_236),
.B1(n_254),
.B2(n_250),
.C(n_239),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_261),
.B(n_267),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_228),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_256),
.C(n_241),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_241),
.C(n_253),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_240),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_252),
.B1(n_242),
.B2(n_258),
.Y(n_273)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_255),
.B(n_240),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_275),
.B(n_278),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_246),
.B(n_240),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_244),
.B1(n_248),
.B2(n_245),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_280),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_243),
.B(n_251),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_265),
.B(n_251),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_281),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_277),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_280),
.B(n_282),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_274),
.B(n_278),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g296 ( 
.A1(n_290),
.A2(n_283),
.B(n_286),
.C(n_288),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_292),
.B(n_294),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_287),
.C(n_281),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_263),
.B1(n_275),
.B2(n_260),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

AOI321xp33_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_291),
.A3(n_297),
.B1(n_293),
.B2(n_296),
.C(n_294),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);


endmodule