module fake_jpeg_3181_n_183 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_18),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_63),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_15),
.C(n_12),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_71),
.Y(n_88)
);

OR2x4_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_23),
.Y(n_100)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_70),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_12),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_27),
.B1(n_13),
.B2(n_21),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_40),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_32),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_86),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_79),
.B(n_84),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_13),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_27),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_32),
.Y(n_86)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_11),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_97),
.Y(n_116)
);

AO22x2_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_42),
.B1(n_40),
.B2(n_17),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_49),
.B(n_54),
.C(n_58),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_2),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_36),
.B1(n_17),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_101),
.A2(n_82),
.B1(n_94),
.B2(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_120),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_119),
.B1(n_96),
.B2(n_87),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_80),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_73),
.B(n_58),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_88),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_90),
.Y(n_125)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_54),
.B1(n_73),
.B2(n_6),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_90),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_133),
.C(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_100),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_77),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_119),
.B1(n_120),
.B2(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_117),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_91),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_110),
.B1(n_105),
.B2(n_106),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_148),
.B(n_135),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_115),
.B(n_111),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_142),
.B(n_133),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_123),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_147),
.C(n_139),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_124),
.B(n_126),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_159),
.Y(n_161)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_151),
.B(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_151),
.B1(n_152),
.B2(n_146),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_137),
.B1(n_111),
.B2(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_165),
.B(n_145),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_167),
.B(n_170),
.Y(n_174)
);

OAI322xp33_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_150),
.A3(n_158),
.B1(n_122),
.B2(n_144),
.C1(n_126),
.C2(n_127),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_162),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_163),
.B(n_164),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_173),
.B(n_161),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_175),
.B(n_176),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_89),
.A3(n_76),
.B1(n_75),
.B2(n_103),
.C1(n_6),
.C2(n_5),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_103),
.B(n_75),
.C(n_76),
.D(n_5),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_81),
.B1(n_80),
.B2(n_171),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_180),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_178),
.C(n_81),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_3),
.Y(n_183)
);


endmodule