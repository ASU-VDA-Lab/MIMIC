module real_aes_9004_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_385;
wire n_214;
wire n_275;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g464 ( .A(n_0), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_1), .A2(n_142), .B(n_146), .C(n_227), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_2), .A2(n_176), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g518 ( .A(n_3), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_4), .B(n_243), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_5), .A2(n_105), .B1(n_117), .B2(n_759), .Y(n_104) );
AOI21xp33_ASAP7_75t_L g483 ( .A1(n_6), .A2(n_176), .B(n_484), .Y(n_483) );
AND2x6_ASAP7_75t_L g142 ( .A(n_7), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g217 ( .A(n_8), .Y(n_217) );
INVx1_ASAP7_75t_L g110 ( .A(n_9), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_9), .B(n_42), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_10), .A2(n_175), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_11), .B(n_154), .Y(n_229) );
INVx1_ASAP7_75t_L g488 ( .A(n_12), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_13), .B(n_257), .Y(n_542) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
INVx1_ASAP7_75t_L g554 ( .A(n_15), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_16), .A2(n_152), .B(n_239), .C(n_241), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_17), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_18), .B(n_506), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_19), .B(n_176), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_20), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_21), .A2(n_257), .B(n_272), .C(n_274), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_22), .B(n_243), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_23), .B(n_154), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_24), .A2(n_184), .B(n_241), .C(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_25), .B(n_154), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_26), .Y(n_193) );
INVx1_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_28), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_29), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_30), .B(n_154), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_31), .A2(n_32), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_31), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_32), .Y(n_752) );
INVx1_ASAP7_75t_L g182 ( .A(n_33), .Y(n_182) );
INVx1_ASAP7_75t_L g497 ( .A(n_34), .Y(n_497) );
INVx2_ASAP7_75t_L g140 ( .A(n_35), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_36), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_37), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
INVxp67_ASAP7_75t_L g183 ( .A(n_38), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_39), .A2(n_146), .B(n_149), .C(n_157), .Y(n_145) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_40), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_142), .B(n_146), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_42), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g496 ( .A(n_43), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_44), .A2(n_201), .B(n_215), .C(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_45), .B(n_154), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_46), .A2(n_749), .B1(n_755), .B2(n_756), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_46), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_47), .A2(n_750), .B1(n_751), .B2(n_754), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_47), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_48), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_49), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_50), .B(n_458), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_51), .A2(n_462), .B1(n_469), .B2(n_757), .Y(n_468) );
INVx1_ASAP7_75t_L g270 ( .A(n_52), .Y(n_270) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_53), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_54), .B(n_176), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_55), .A2(n_146), .B1(n_274), .B2(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_56), .A2(n_71), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_56), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_57), .Y(n_515) );
CKINVDCx14_ASAP7_75t_R g213 ( .A(n_58), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_59), .A2(n_215), .B(n_260), .C(n_487), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_60), .Y(n_570) );
INVx1_ASAP7_75t_L g485 ( .A(n_61), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_62), .A2(n_91), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_62), .Y(n_457) );
INVx1_ASAP7_75t_L g143 ( .A(n_63), .Y(n_143) );
INVx1_ASAP7_75t_L g161 ( .A(n_64), .Y(n_161) );
INVx1_ASAP7_75t_SL g259 ( .A(n_65), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_66), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_67), .B(n_243), .Y(n_276) );
INVx1_ASAP7_75t_L g196 ( .A(n_68), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_SL g505 ( .A1(n_69), .A2(n_260), .B(n_506), .C(n_507), .Y(n_505) );
INVxp67_ASAP7_75t_L g508 ( .A(n_70), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_71), .Y(n_127) );
INVx1_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_73), .A2(n_176), .B(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_74), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_75), .A2(n_176), .B(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_76), .Y(n_500) );
INVx1_ASAP7_75t_L g564 ( .A(n_77), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_78), .A2(n_175), .B(n_177), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_79), .Y(n_144) );
INVx1_ASAP7_75t_L g237 ( .A(n_80), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_81), .A2(n_142), .B(n_146), .C(n_566), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_82), .A2(n_176), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g240 ( .A(n_83), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_84), .B(n_151), .Y(n_531) );
INVx2_ASAP7_75t_L g159 ( .A(n_85), .Y(n_159) );
INVx1_ASAP7_75t_L g228 ( .A(n_86), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_87), .B(n_506), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_88), .A2(n_142), .B(n_146), .C(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
OR2x2_ASAP7_75t_L g461 ( .A(n_89), .B(n_462), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_90), .A2(n_146), .B(n_195), .C(n_203), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_91), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_92), .B(n_158), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_93), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_94), .A2(n_142), .B(n_146), .C(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_95), .Y(n_546) );
INVx1_ASAP7_75t_L g504 ( .A(n_96), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_97), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_98), .B(n_151), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_99), .B(n_166), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_100), .B(n_166), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_101), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g273 ( .A(n_102), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_103), .A2(n_176), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g759 ( .A(n_107), .Y(n_759) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g471 ( .A(n_113), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_113), .Y(n_474) );
NOR2x2_ASAP7_75t_L g757 ( .A(n_113), .B(n_462), .Y(n_757) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_467), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_SL g758 ( .A(n_120), .Y(n_758) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_458), .B(n_466), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_129), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_SL g533 ( .A(n_126), .B(n_165), .Y(n_533) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
XOR2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_455), .Y(n_129) );
INVx2_ASAP7_75t_L g472 ( .A(n_130), .Y(n_472) );
OR4x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_345), .C(n_392), .D(n_432), .Y(n_130) );
NAND3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_291), .C(n_320), .Y(n_131) );
AOI211xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_206), .B(n_244), .C(n_284), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_133), .A2(n_304), .B(n_321), .C(n_325), .Y(n_320) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_135), .B(n_283), .Y(n_282) );
INVx3_ASAP7_75t_SL g287 ( .A(n_135), .Y(n_287) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_135), .Y(n_299) );
AND2x4_ASAP7_75t_L g303 ( .A(n_135), .B(n_251), .Y(n_303) );
AND2x2_ASAP7_75t_L g314 ( .A(n_135), .B(n_191), .Y(n_314) );
OR2x2_ASAP7_75t_L g338 ( .A(n_135), .B(n_247), .Y(n_338) );
AND2x2_ASAP7_75t_L g351 ( .A(n_135), .B(n_252), .Y(n_351) );
AND2x2_ASAP7_75t_L g391 ( .A(n_135), .B(n_377), .Y(n_391) );
AND2x2_ASAP7_75t_L g398 ( .A(n_135), .B(n_361), .Y(n_398) );
AND2x2_ASAP7_75t_L g428 ( .A(n_135), .B(n_169), .Y(n_428) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_163), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_145), .C(n_158), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_137), .A2(n_193), .B(n_194), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_137), .A2(n_225), .B(n_226), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_137), .A2(n_186), .B1(n_494), .B2(n_498), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_137), .A2(n_515), .B(n_516), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_137), .A2(n_564), .B(n_565), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
AND2x4_ASAP7_75t_L g176 ( .A(n_138), .B(n_142), .Y(n_176) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g156 ( .A(n_139), .Y(n_156) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g147 ( .A(n_140), .Y(n_147) );
INVx1_ASAP7_75t_L g275 ( .A(n_140), .Y(n_275) );
INVx1_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
INVx3_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
INVx1_ASAP7_75t_L g506 ( .A(n_141), .Y(n_506) );
BUFx3_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
INVx4_ASAP7_75t_SL g186 ( .A(n_142), .Y(n_186) );
INVx5_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g202 ( .A(n_147), .Y(n_202) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_147), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_153), .C(n_155), .Y(n_149) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_151), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_151), .A2(n_518), .B(n_519), .C(n_520), .Y(n_517) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_152), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_152), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_152), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g215 ( .A(n_154), .Y(n_215) );
INVx4_ASAP7_75t_L g257 ( .A(n_154), .Y(n_257) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_156), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_211), .B(n_218), .Y(n_210) );
INVx1_ASAP7_75t_L g223 ( .A(n_158), .Y(n_223) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_158), .A2(n_549), .B(n_555), .Y(n_548) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_L g167 ( .A(n_159), .B(n_160), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_165), .A2(n_192), .B(n_204), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_165), .B(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g243 ( .A(n_165), .Y(n_243) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_166), .Y(n_234) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_166), .A2(n_502), .B(n_509), .Y(n_501) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_168), .B(n_355), .Y(n_367) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_190), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_169), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_169), .B(n_190), .Y(n_305) );
BUFx3_ASAP7_75t_L g313 ( .A(n_169), .Y(n_313) );
OR2x2_ASAP7_75t_L g334 ( .A(n_169), .B(n_209), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_169), .B(n_355), .Y(n_445) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_174), .B(n_187), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_171), .A2(n_248), .B(n_249), .Y(n_247) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_171), .A2(n_563), .B(n_569), .Y(n_562) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g527 ( .A1(n_172), .A2(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_173), .A2(n_493), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_173), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_173), .A2(n_514), .B(n_521), .Y(n_513) );
INVx1_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_179), .B(n_180), .C(n_186), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g212 ( .A1(n_179), .A2(n_186), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_179), .A2(n_186), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_179), .A2(n_186), .B(n_255), .C(n_256), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g269 ( .A1(n_179), .A2(n_186), .B(n_270), .C(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g484 ( .A1(n_179), .A2(n_186), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_179), .A2(n_186), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_179), .A2(n_186), .B(n_551), .C(n_552), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_184), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_184), .B(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_184), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g198 ( .A(n_185), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_185), .A2(n_198), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g203 ( .A(n_186), .Y(n_203) );
INVx1_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_189), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_189), .A2(n_538), .B(n_545), .Y(n_537) );
AND2x2_ASAP7_75t_L g250 ( .A(n_190), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g298 ( .A(n_190), .Y(n_298) );
AND2x2_ASAP7_75t_L g361 ( .A(n_190), .B(n_252), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_190), .A2(n_364), .B1(n_366), .B2(n_368), .C(n_369), .Y(n_363) );
AND2x2_ASAP7_75t_L g377 ( .A(n_190), .B(n_247), .Y(n_377) );
AND2x2_ASAP7_75t_L g403 ( .A(n_190), .B(n_287), .Y(n_403) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g283 ( .A(n_191), .B(n_252), .Y(n_283) );
BUFx2_ASAP7_75t_L g417 ( .A(n_191), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_200), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_200), .B(n_228), .C(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_200), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_200), .A2(n_567), .B(n_568), .Y(n_566) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OAI32xp33_ASAP7_75t_L g383 ( .A1(n_207), .A2(n_344), .A3(n_358), .B1(n_384), .B2(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
AND2x2_ASAP7_75t_L g324 ( .A(n_208), .B(n_266), .Y(n_324) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g306 ( .A(n_209), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_209), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g378 ( .A(n_209), .B(n_266), .Y(n_378) );
AND2x2_ASAP7_75t_L g389 ( .A(n_209), .B(n_281), .Y(n_389) );
BUFx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g290 ( .A(n_210), .B(n_267), .Y(n_290) );
AND2x2_ASAP7_75t_L g294 ( .A(n_210), .B(n_267), .Y(n_294) );
AND2x2_ASAP7_75t_L g329 ( .A(n_210), .B(n_280), .Y(n_329) );
AND2x2_ASAP7_75t_L g336 ( .A(n_210), .B(n_232), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g341 ( .A1(n_210), .A2(n_287), .B(n_298), .C(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g395 ( .A(n_210), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_210), .B(n_221), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_219), .B(n_278), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_219), .B(n_294), .Y(n_384) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
OR2x2_ASAP7_75t_L g289 ( .A(n_220), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_232), .Y(n_220) );
AND2x2_ASAP7_75t_L g281 ( .A(n_221), .B(n_233), .Y(n_281) );
OR2x2_ASAP7_75t_L g296 ( .A(n_221), .B(n_233), .Y(n_296) );
AND2x2_ASAP7_75t_L g319 ( .A(n_221), .B(n_280), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_221), .Y(n_323) );
AND2x2_ASAP7_75t_L g342 ( .A(n_221), .B(n_279), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_221), .A2(n_307), .B1(n_353), .B2(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_221), .B(n_395), .Y(n_419) );
AND2x2_ASAP7_75t_L g434 ( .A(n_221), .B(n_294), .Y(n_434) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx3_ASAP7_75t_L g264 ( .A(n_222), .Y(n_264) );
AND2x2_ASAP7_75t_L g308 ( .A(n_222), .B(n_233), .Y(n_308) );
AND2x2_ASAP7_75t_L g310 ( .A(n_222), .B(n_266), .Y(n_310) );
AND3x2_ASAP7_75t_L g372 ( .A(n_222), .B(n_336), .C(n_373), .Y(n_372) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_230), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_223), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_223), .B(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_223), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g407 ( .A(n_232), .B(n_279), .Y(n_407) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g266 ( .A(n_233), .B(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_233), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_233), .B(n_278), .Y(n_340) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_233), .B(n_319), .C(n_395), .Y(n_447) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_242), .Y(n_233) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_234), .A2(n_253), .B(n_262), .Y(n_252) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_234), .A2(n_268), .B(n_276), .Y(n_267) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_243), .A2(n_483), .B(n_489), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_263), .B1(n_277), .B2(n_282), .Y(n_244) );
INVx1_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_247), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g359 ( .A(n_247), .Y(n_359) );
OAI31xp33_ASAP7_75t_L g375 ( .A1(n_250), .A2(n_376), .A3(n_377), .B(n_378), .Y(n_375) );
AND2x2_ASAP7_75t_L g400 ( .A(n_250), .B(n_287), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_250), .B(n_313), .Y(n_446) );
AND2x2_ASAP7_75t_L g355 ( .A(n_251), .B(n_287), .Y(n_355) );
AND2x2_ASAP7_75t_L g416 ( .A(n_251), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g286 ( .A(n_252), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g344 ( .A(n_252), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_261), .Y(n_543) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_264), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_265), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AOI221x1_ASAP7_75t_SL g332 ( .A1(n_266), .A2(n_333), .B1(n_335), .B2(n_337), .C(n_339), .Y(n_332) );
INVx2_ASAP7_75t_L g280 ( .A(n_267), .Y(n_280) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_267), .Y(n_374) );
INVx2_ASAP7_75t_L g520 ( .A(n_274), .Y(n_520) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g362 ( .A(n_277), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_278), .B(n_295), .Y(n_387) );
INVx1_ASAP7_75t_SL g450 ( .A(n_278), .Y(n_450) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g368 ( .A(n_281), .B(n_294), .Y(n_368) );
INVx1_ASAP7_75t_L g436 ( .A(n_282), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_282), .B(n_365), .Y(n_449) );
INVx2_ASAP7_75t_SL g288 ( .A(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g331 ( .A(n_283), .B(n_287), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_283), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_283), .B(n_358), .Y(n_385) );
AOI21xp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B(n_289), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_286), .B(n_358), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_286), .B(n_313), .Y(n_454) );
OR2x2_ASAP7_75t_L g326 ( .A(n_287), .B(n_305), .Y(n_326) );
AND2x2_ASAP7_75t_L g425 ( .A(n_287), .B(n_416), .Y(n_425) );
OAI22xp5_ASAP7_75t_SL g300 ( .A1(n_288), .A2(n_301), .B1(n_306), .B2(n_309), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_288), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g348 ( .A(n_290), .B(n_296), .Y(n_348) );
INVx1_ASAP7_75t_L g412 ( .A(n_290), .Y(n_412) );
AOI311xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_297), .A3(n_299), .B(n_300), .C(n_311), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_295), .A2(n_427), .B1(n_439), .B2(n_442), .C(n_444), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_295), .B(n_450), .Y(n_452) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_298), .A2(n_340), .B(n_341), .C(n_343), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_SL g408 ( .A1(n_302), .A2(n_304), .B(n_409), .C(n_410), .Y(n_408) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_303), .B(n_377), .Y(n_443) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_306), .A2(n_326), .B1(n_327), .B2(n_330), .C(n_332), .Y(n_325) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g328 ( .A(n_308), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g411 ( .A(n_308), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_312), .A2(n_370), .B(n_371), .C(n_375), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_313), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_313), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVxp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g335 ( .A(n_319), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_323), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g437 ( .A(n_326), .Y(n_437) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_329), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_329), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g441 ( .A(n_329), .Y(n_441) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g382 ( .A(n_331), .B(n_358), .Y(n_382) );
INVx1_ASAP7_75t_SL g376 ( .A(n_338), .Y(n_376) );
INVx1_ASAP7_75t_L g353 ( .A(n_344), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g345 ( .A(n_346), .B(n_363), .C(n_379), .Y(n_345) );
AOI322xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .A3(n_350), .B1(n_352), .B2(n_356), .C1(n_360), .C2(n_362), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g399 ( .A1(n_347), .A2(n_400), .B(n_401), .C(n_408), .Y(n_399) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_350), .A2(n_371), .B1(n_402), .B2(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g360 ( .A(n_358), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g397 ( .A(n_358), .B(n_398), .Y(n_397) );
AOI32xp33_ASAP7_75t_L g448 ( .A1(n_358), .A2(n_449), .A3(n_450), .B1(n_451), .B2(n_453), .Y(n_448) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g370 ( .A(n_361), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_361), .A2(n_414), .B1(n_418), .B2(n_420), .C(n_423), .Y(n_413) );
AND2x2_ASAP7_75t_L g427 ( .A(n_361), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g430 ( .A(n_365), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g440 ( .A(n_365), .B(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g431 ( .A(n_374), .B(n_395), .Y(n_431) );
AOI211xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B(n_383), .C(n_386), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_396), .B(n_399), .C(n_413), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_407), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g422 ( .A(n_419), .Y(n_422) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B(n_429), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_435), .B(n_438), .C(n_448), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_466), .A2(n_468), .B(n_758), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_748), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_473), .B2(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND3x1_ASAP7_75t_L g477 ( .A(n_478), .B(n_670), .C(n_715), .Y(n_477) );
NOR4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_593), .C(n_634), .D(n_651), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_510), .B(n_524), .C(n_556), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_490), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_481), .B(n_511), .Y(n_510) );
NOR4xp25_ASAP7_75t_L g617 ( .A(n_481), .B(n_611), .C(n_618), .D(n_624), .Y(n_617) );
AND2x2_ASAP7_75t_L g690 ( .A(n_481), .B(n_579), .Y(n_690) );
AND2x2_ASAP7_75t_L g709 ( .A(n_481), .B(n_655), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_481), .B(n_704), .Y(n_718) );
AND2x2_ASAP7_75t_L g731 ( .A(n_481), .B(n_523), .Y(n_731) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g576 ( .A(n_482), .Y(n_576) );
AND2x2_ASAP7_75t_L g583 ( .A(n_482), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g633 ( .A(n_482), .B(n_491), .Y(n_633) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_482), .B(n_579), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_482), .B(n_491), .Y(n_648) );
AND2x2_ASAP7_75t_L g657 ( .A(n_482), .B(n_582), .Y(n_657) );
BUFx2_ASAP7_75t_L g680 ( .A(n_482), .Y(n_680) );
AND2x2_ASAP7_75t_L g684 ( .A(n_482), .B(n_501), .Y(n_684) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
AND2x2_ASAP7_75t_L g523 ( .A(n_491), .B(n_501), .Y(n_523) );
BUFx2_ASAP7_75t_L g586 ( .A(n_491), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_491), .A2(n_619), .B1(n_621), .B2(n_622), .Y(n_618) );
OR2x2_ASAP7_75t_L g640 ( .A(n_491), .B(n_513), .Y(n_640) );
AND2x2_ASAP7_75t_L g704 ( .A(n_491), .B(n_582), .Y(n_704) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g572 ( .A(n_492), .B(n_513), .Y(n_572) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_501), .Y(n_579) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_492), .Y(n_621) );
OR2x2_ASAP7_75t_L g656 ( .A(n_492), .B(n_512), .Y(n_656) );
INVx1_ASAP7_75t_L g575 ( .A(n_501), .Y(n_575) );
INVx3_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
BUFx2_ASAP7_75t_L g608 ( .A(n_501), .Y(n_608) );
AND2x2_ASAP7_75t_L g641 ( .A(n_501), .B(n_576), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_510), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_512), .B(n_584), .Y(n_588) );
INVx1_ASAP7_75t_L g616 ( .A(n_512), .Y(n_616) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g582 ( .A(n_513), .Y(n_582) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
NAND2x1_ASAP7_75t_SL g524 ( .A(n_525), .B(n_534), .Y(n_524) );
AND2x2_ASAP7_75t_L g592 ( .A(n_525), .B(n_547), .Y(n_592) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_525), .Y(n_666) );
AND2x2_ASAP7_75t_L g693 ( .A(n_525), .B(n_613), .Y(n_693) );
AND2x2_ASAP7_75t_L g701 ( .A(n_525), .B(n_663), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_525), .B(n_559), .Y(n_728) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g560 ( .A(n_526), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g598 ( .A(n_526), .Y(n_598) );
INVx1_ASAP7_75t_L g604 ( .A(n_526), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_526), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_562), .Y(n_637) );
OR2x2_ASAP7_75t_L g675 ( .A(n_526), .B(n_630), .Y(n_675) );
AOI32xp33_ASAP7_75t_L g687 ( .A1(n_526), .A2(n_688), .A3(n_691), .B1(n_692), .B2(n_693), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_526), .B(n_663), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_526), .B(n_623), .Y(n_738) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_533), .Y(n_526) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g649 ( .A(n_535), .B(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_547), .Y(n_535) );
INVx1_ASAP7_75t_L g611 ( .A(n_536), .Y(n_611) );
AND2x2_ASAP7_75t_L g613 ( .A(n_536), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_536), .B(n_561), .Y(n_630) );
AND2x2_ASAP7_75t_L g663 ( .A(n_536), .B(n_639), .Y(n_663) );
AND2x2_ASAP7_75t_L g700 ( .A(n_536), .B(n_562), .Y(n_700) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g559 ( .A(n_537), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_537), .B(n_561), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_537), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g638 ( .A(n_537), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_544), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_543), .Y(n_540) );
INVx2_ASAP7_75t_L g614 ( .A(n_547), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_547), .B(n_561), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_547), .B(n_605), .Y(n_686) );
INVx1_ASAP7_75t_L g708 ( .A(n_547), .Y(n_708) );
INVx1_ASAP7_75t_L g725 ( .A(n_547), .Y(n_725) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g578 ( .A(n_548), .B(n_561), .Y(n_578) );
AND2x2_ASAP7_75t_L g600 ( .A(n_548), .B(n_562), .Y(n_600) );
INVx1_ASAP7_75t_L g639 ( .A(n_548), .Y(n_639) );
AOI221x1_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_571), .B1(n_577), .B2(n_579), .C(n_580), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_557), .A2(n_644), .B1(n_711), .B2(n_712), .Y(n_710) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g602 ( .A(n_558), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g697 ( .A(n_558), .B(n_577), .Y(n_697) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g653 ( .A(n_559), .B(n_578), .Y(n_653) );
INVx1_ASAP7_75t_L g665 ( .A(n_560), .Y(n_665) );
AND2x2_ASAP7_75t_L g676 ( .A(n_560), .B(n_663), .Y(n_676) );
AND2x2_ASAP7_75t_L g743 ( .A(n_560), .B(n_638), .Y(n_743) );
INVx2_ASAP7_75t_L g605 ( .A(n_561), .Y(n_605) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_572), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g695 ( .A(n_572), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_573), .B(n_656), .Y(n_659) );
INVx3_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_574), .A2(n_695), .B(n_740), .Y(n_739) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NOR2xp33_ASAP7_75t_SL g717 ( .A(n_577), .B(n_603), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_578), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g669 ( .A(n_578), .B(n_597), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_578), .B(n_604), .Y(n_746) );
AND2x2_ASAP7_75t_L g615 ( .A(n_579), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g682 ( .A(n_579), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B(n_589), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_582), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g631 ( .A(n_582), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g643 ( .A(n_582), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_582), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g667 ( .A(n_583), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_583), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_583), .B(n_586), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_586), .A2(n_625), .B(n_655), .C(n_657), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_586), .A2(n_673), .B1(n_676), .B2(n_677), .C(n_681), .Y(n_672) );
AND2x2_ASAP7_75t_L g668 ( .A(n_587), .B(n_621), .Y(n_668) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g628 ( .A(n_592), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g699 ( .A(n_592), .B(n_700), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_601), .C(n_626), .Y(n_593) );
NAND3xp33_ASAP7_75t_SL g712 ( .A(n_594), .B(n_713), .C(n_714), .Y(n_712) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_599), .Y(n_595) );
OR2x2_ASAP7_75t_L g685 ( .A(n_596), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .B1(n_609), .B2(n_615), .C(n_617), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_603), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_603), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g625 ( .A(n_608), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_608), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g745 ( .A(n_608), .B(n_656), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVxp67_ASAP7_75t_L g719 ( .A(n_611), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_613), .B(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g620 ( .A(n_614), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_616), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_616), .B(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_616), .B(n_683), .Y(n_722) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_620), .Y(n_646) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g736 ( .A(n_625), .B(n_656), .Y(n_736) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g714 ( .A(n_631), .Y(n_714) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI322xp33_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_640), .A3(n_641), .B1(n_642), .B2(n_645), .C1(n_647), .C2(n_649), .Y(n_634) );
OAI322xp33_ASAP7_75t_L g716 ( .A1(n_635), .A2(n_717), .A3(n_718), .B1(n_719), .B2(n_720), .C1(n_721), .C2(n_723), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx4_ASAP7_75t_L g650 ( .A(n_637), .Y(n_650) );
AND2x2_ASAP7_75t_L g711 ( .A(n_637), .B(n_663), .Y(n_711) );
AND2x2_ASAP7_75t_L g724 ( .A(n_637), .B(n_725), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_640), .Y(n_735) );
INVx1_ASAP7_75t_L g713 ( .A(n_641), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
OR2x2_ASAP7_75t_L g647 ( .A(n_643), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g730 ( .A(n_643), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_643), .B(n_684), .Y(n_741) );
OR2x2_ASAP7_75t_L g674 ( .A(n_646), .B(n_675), .Y(n_674) );
INVxp33_ASAP7_75t_L g691 ( .A(n_646), .Y(n_691) );
OAI221xp5_ASAP7_75t_SL g651 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_658), .C(n_660), .Y(n_651) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_650), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g734 ( .A(n_650), .Y(n_734) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVx3_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_657), .A2(n_682), .A3(n_699), .B1(n_701), .B2(n_702), .C1(n_705), .C2(n_709), .Y(n_698) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B1(n_668), .B2(n_669), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_694), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_672), .B(n_687), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_675), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NAND2xp33_ASAP7_75t_SL g692 ( .A(n_678), .B(n_689), .Y(n_692) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g732 ( .A1(n_680), .A2(n_733), .A3(n_735), .B1(n_736), .B2(n_737), .C1(n_739), .C2(n_742), .Y(n_732) );
AOI21xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_690), .B(n_738), .Y(n_747) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_696), .B(n_698), .C(n_710), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NOR4xp25_ASAP7_75t_L g715 ( .A(n_716), .B(n_726), .C(n_732), .D(n_744), .Y(n_715) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx14_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
OAI21xp5_ASAP7_75t_SL g744 ( .A1(n_745), .A2(n_746), .B(n_747), .Y(n_744) );
CKINVDCx16_ASAP7_75t_R g756 ( .A(n_749), .Y(n_756) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
endmodule