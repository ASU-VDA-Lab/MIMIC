module fake_jpeg_26653_n_248 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_24),
.B(n_32),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_52),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_18),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_22),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_44),
.B1(n_41),
.B2(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_24),
.B(n_34),
.C(n_30),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_19),
.Y(n_87)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_39),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_72),
.B1(n_73),
.B2(n_31),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_79),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_67),
.B1(n_84),
.B2(n_90),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_41),
.B1(n_43),
.B2(n_18),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_37),
.B1(n_30),
.B2(n_20),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_33),
.B1(n_35),
.B2(n_21),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_92),
.B1(n_21),
.B2(n_26),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_45),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_33),
.B1(n_35),
.B2(n_20),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_17),
.B(n_25),
.C(n_31),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_118),
.B(n_70),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_53),
.B1(n_38),
.B2(n_39),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_53),
.B1(n_38),
.B2(n_39),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_53),
.B1(n_39),
.B2(n_31),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_35),
.Y(n_109)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_80),
.B1(n_77),
.B2(n_74),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_26),
.B1(n_17),
.B2(n_33),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_112),
.A2(n_29),
.B1(n_51),
.B2(n_62),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

XOR2x1_ASAP7_75t_SL g118 ( 
.A(n_82),
.B(n_28),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_75),
.C(n_94),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_131),
.C(n_133),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_91),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_139),
.B(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_88),
.B1(n_80),
.B2(n_86),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_146),
.B1(n_106),
.B2(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_136),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_97),
.C(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_85),
.C(n_64),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_115),
.B1(n_100),
.B2(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_70),
.C(n_93),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_143),
.C(n_81),
.Y(n_166)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_114),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_60),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_108),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_80),
.B1(n_77),
.B2(n_74),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_100),
.B1(n_112),
.B2(n_104),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_29),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_153),
.B1(n_10),
.B2(n_12),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_95),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_2),
.B(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_152),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_155),
.B1(n_162),
.B2(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_144),
.B1(n_123),
.B2(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_95),
.B1(n_110),
.B2(n_102),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_163),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_129),
.A2(n_108),
.B(n_2),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_SL g182 ( 
.A1(n_161),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_123),
.A2(n_51),
.B1(n_29),
.B2(n_81),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_125),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_81),
.B(n_2),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_7),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_132),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_1),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_153),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_126),
.C(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_171),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_29),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_189),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_168),
.B(n_169),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_186),
.B(n_10),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_191),
.B1(n_160),
.B2(n_148),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_9),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_166),
.C(n_157),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_9),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_198),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_207),
.B(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_155),
.B1(n_148),
.B2(n_150),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_200),
.B1(n_162),
.B2(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_152),
.C(n_156),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.C(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_156),
.C(n_149),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

AOI21x1_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_160),
.B(n_181),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_215),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_174),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_216),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_158),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_151),
.B1(n_170),
.B2(n_189),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_195),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_227),
.C(n_229),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_214),
.B(n_210),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_188),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_202),
.B1(n_192),
.B2(n_198),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_175),
.C(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_227),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_232),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_221),
.A2(n_213),
.B(n_208),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_212),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_223),
.B(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.C(n_233),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_192),
.B(n_14),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_236),
.B1(n_14),
.B2(n_16),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_12),
.C(n_245),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_12),
.Y(n_248)
);


endmodule