module fake_jpeg_4049_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_33),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_34),
.B1(n_29),
.B2(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_30),
.B1(n_34),
.B2(n_41),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_23),
.B1(n_35),
.B2(n_18),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_20),
.Y(n_77)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_79),
.Y(n_108)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_22),
.B1(n_35),
.B2(n_19),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_17),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_17),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_26),
.Y(n_117)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_57),
.B1(n_66),
.B2(n_50),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_47),
.B1(n_63),
.B2(n_27),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_32),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_111),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_18),
.C(n_21),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_51),
.B1(n_72),
.B2(n_67),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_64),
.B1(n_63),
.B2(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_113),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_64),
.B1(n_27),
.B2(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_24),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_19),
.Y(n_148)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_126),
.B1(n_128),
.B2(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_55),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_73),
.B1(n_24),
.B2(n_22),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_42),
.B1(n_36),
.B2(n_37),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_55),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_79),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_153),
.B1(n_154),
.B2(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_136),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_144),
.C(n_147),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_146),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_124),
.Y(n_170)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_143),
.B1(n_149),
.B2(n_120),
.Y(n_175)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_36),
.C(n_37),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_32),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_117),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_97),
.B1(n_91),
.B2(n_90),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_97),
.C(n_96),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_101),
.A2(n_71),
.B1(n_21),
.B2(n_32),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_71),
.B1(n_96),
.B2(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_0),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_148),
.B1(n_119),
.B2(n_105),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_160),
.B(n_163),
.Y(n_194)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_166),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_171),
.B1(n_178),
.B2(n_154),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_167),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_179),
.C(n_180),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_172),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_182),
.B(n_176),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_124),
.B1(n_114),
.B2(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_176),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_108),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_137),
.B(n_152),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_158),
.B(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_108),
.B1(n_128),
.B2(n_110),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_115),
.B(n_110),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_131),
.B(n_120),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_115),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_134),
.C(n_16),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_187),
.A2(n_191),
.B1(n_201),
.B2(n_208),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_151),
.B1(n_145),
.B2(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_213),
.B1(n_186),
.B2(n_172),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_195),
.B(n_203),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_179),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_199),
.C(n_206),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_138),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_159),
.A2(n_105),
.B1(n_134),
.B2(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_211),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_163),
.A2(n_0),
.B(n_2),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_183),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_217),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_223),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_158),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_231),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_214),
.B1(n_200),
.B2(n_190),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_235),
.B1(n_198),
.B2(n_188),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_181),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_229),
.B(n_240),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_193),
.B(n_170),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_236),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_167),
.B1(n_170),
.B2(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_3),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_196),
.B(n_14),
.Y(n_241)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_234),
.A2(n_188),
.B1(n_193),
.B2(n_198),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_248),
.B1(n_262),
.B2(n_264),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_192),
.B(n_203),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_262),
.B(n_7),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_206),
.C(n_4),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_259),
.C(n_265),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_248)
);

AOI211xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_10),
.B(n_13),
.C(n_12),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_231),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_10),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_230),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_220),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_5),
.B(n_7),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_232),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_7),
.C(n_8),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_225),
.CI(n_218),
.CON(n_266),
.SN(n_266)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_277),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_242),
.CI(n_251),
.CON(n_288),
.SN(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_243),
.B(n_215),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_283),
.B1(n_248),
.B2(n_255),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_247),
.B(n_218),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_243),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_222),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_216),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_251),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_236),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_249),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_250),
.C(n_244),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_289),
.C(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_260),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_250),
.C(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_284),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_221),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_252),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_259),
.C(n_254),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_245),
.C(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_285),
.C(n_289),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_304),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_266),
.C(n_274),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_310),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_266),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_314),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_308),
.B(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_276),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_300),
.B1(n_267),
.B2(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_313),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_306),
.B1(n_310),
.B2(n_299),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_257),
.B1(n_255),
.B2(n_268),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_287),
.B(n_268),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_288),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_304),
.B(n_296),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_303),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_305),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_307),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_261),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_11),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_10),
.C(n_11),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_323),
.B(n_315),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_335),
.B(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_333),
.A2(n_326),
.B(n_12),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_12),
.B(n_13),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_338),
.B(n_336),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_8),
.C(n_9),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_14),
.B(n_8),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_8),
.B(n_9),
.Y(n_344)
);


endmodule