module fake_jpeg_13724_n_594 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_594);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_594;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_58),
.B(n_86),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_67),
.Y(n_120)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_38),
.B(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_20),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g171 ( 
.A(n_68),
.Y(n_171)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_39),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_89),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_87),
.Y(n_118)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_18),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_28),
.B(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_94),
.Y(n_119)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_29),
.B(n_0),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_30),
.B(n_49),
.Y(n_140)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_21),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_27),
.B(n_16),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_108),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_21),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_27),
.B(n_16),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_49),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_23),
.B1(n_53),
.B2(n_36),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_112),
.A2(n_121),
.B1(n_174),
.B2(n_34),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_64),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_113),
.B(n_159),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_53),
.B1(n_36),
.B2(n_47),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx5_ASAP7_75t_SL g235 ( 
.A(n_122),
.Y(n_235)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_92),
.A2(n_44),
.B1(n_47),
.B2(n_54),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_133),
.A2(n_153),
.B1(n_42),
.B2(n_31),
.Y(n_197)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_140),
.B(n_34),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_92),
.A2(n_44),
.B1(n_47),
.B2(n_54),
.Y(n_153)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_56),
.B(n_53),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_85),
.C(n_83),
.Y(n_206)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_79),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_84),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_34),
.Y(n_192)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_36),
.B1(n_34),
.B2(n_48),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_107),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_177),
.B(n_186),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_82),
.B1(n_91),
.B2(n_102),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_178),
.A2(n_207),
.B1(n_213),
.B2(n_217),
.Y(n_270)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_183),
.Y(n_295)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_184),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_130),
.B(n_95),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_189),
.B(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_210),
.C(n_216),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_88),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_196),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_197),
.A2(n_218),
.B1(n_236),
.B2(n_42),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_206),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_57),
.B1(n_62),
.B2(n_65),
.Y(n_199)
);

NAND2x1p5_ASAP7_75t_L g281 ( 
.A(n_199),
.B(n_175),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_135),
.B(n_32),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_204),
.Y(n_279)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_119),
.B(n_45),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_205),
.Y(n_284)
);

AO22x2_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_106),
.B1(n_105),
.B2(n_98),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_161),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_116),
.B1(n_141),
.B2(n_117),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_96),
.B1(n_75),
.B2(n_74),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_114),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_214),
.Y(n_264)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_124),
.B(n_30),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_147),
.A2(n_60),
.B1(n_72),
.B2(n_55),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_112),
.B1(n_121),
.B2(n_59),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_127),
.A2(n_63),
.B1(n_76),
.B2(n_33),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_223),
.A2(n_138),
.B1(n_168),
.B2(n_143),
.Y(n_286)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_33),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_137),
.B(n_45),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_42),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_146),
.B(n_69),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_166),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_80),
.Y(n_230)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_44),
.Y(n_232)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_233),
.Y(n_292)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_144),
.Y(n_234)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_116),
.A2(n_44),
.B1(n_48),
.B2(n_46),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_111),
.A2(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_31),
.C(n_25),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_240),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_111),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_282),
.C(n_296),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_249),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_254),
.A2(n_289),
.B1(n_217),
.B2(n_239),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_207),
.A2(n_141),
.B1(n_125),
.B2(n_149),
.Y(n_259)
);

CKINVDCx6p67_ASAP7_75t_R g308 ( 
.A(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_261),
.B(n_26),
.Y(n_310)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_207),
.B(n_199),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_262),
.B(n_281),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_155),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_265),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_155),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_251),
.B1(n_296),
.B2(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_186),
.B(n_147),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_278),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_138),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_199),
.B(n_125),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_286),
.A2(n_208),
.B1(n_26),
.B2(n_25),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_218),
.A2(n_123),
.B1(n_168),
.B2(n_143),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_206),
.B(n_123),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_291),
.B(n_293),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_199),
.B(n_150),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_235),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_235),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_220),
.B(n_149),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_304),
.Y(n_364)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_301),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_261),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_254),
.A2(n_263),
.B1(n_265),
.B2(n_293),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_306),
.A2(n_312),
.B1(n_327),
.B2(n_288),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_181),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_309),
.B(n_310),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_292),
.B(n_200),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_313),
.B(n_326),
.Y(n_394)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_185),
.B1(n_194),
.B2(n_209),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_316),
.A2(n_319),
.B1(n_1),
.B2(n_2),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_251),
.A2(n_200),
.B(n_205),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_317),
.A2(n_281),
.B(n_274),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_242),
.B(n_188),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_318),
.B(n_321),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_270),
.A2(n_184),
.B1(n_222),
.B2(n_187),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_322),
.B(n_332),
.Y(n_380)
);

AO22x1_ASAP7_75t_SL g323 ( 
.A1(n_262),
.A2(n_203),
.B1(n_215),
.B2(n_237),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_333),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_250),
.B(n_188),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_289),
.A2(n_151),
.B1(n_150),
.B2(n_201),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_251),
.A2(n_182),
.B(n_238),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_282),
.B(n_274),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_329),
.A2(n_340),
.B1(n_344),
.B2(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_271),
.B(n_211),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_330),
.B(n_341),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_243),
.B(n_279),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_278),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_342),
.Y(n_354)
);

MAJx2_ASAP7_75t_L g335 ( 
.A(n_260),
.B(n_228),
.C(n_182),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_335),
.B(n_255),
.C(n_285),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_267),
.B(n_211),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_336),
.Y(n_368)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

AND2x6_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_219),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_272),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_345),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_256),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_275),
.Y(n_345)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_347),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_391)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_176),
.Y(n_385)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_349),
.A2(n_240),
.B1(n_179),
.B2(n_283),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_325),
.A2(n_291),
.B1(n_281),
.B2(n_244),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_352),
.A2(n_361),
.B1(n_363),
.B2(n_388),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_371),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_345),
.Y(n_415)
);

AO32x1_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_268),
.A3(n_296),
.B1(n_276),
.B2(n_284),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_357),
.B(n_332),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_339),
.A2(n_325),
.B(n_302),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_359),
.A2(n_369),
.B(n_378),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_308),
.A2(n_286),
.B1(n_247),
.B2(n_288),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_362),
.A2(n_382),
.B1(n_383),
.B2(n_387),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_308),
.A2(n_269),
.B1(n_248),
.B2(n_273),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_302),
.A2(n_255),
.B(n_290),
.Y(n_369)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_246),
.C(n_283),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_373),
.B(n_381),
.C(n_390),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_180),
.B(n_183),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_300),
.B(n_180),
.C(n_221),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_306),
.A2(n_248),
.B1(n_273),
.B2(n_196),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_333),
.A2(n_46),
.B1(n_43),
.B2(n_31),
.Y(n_383)
);

OAI32xp33_ASAP7_75t_L g384 ( 
.A1(n_324),
.A2(n_43),
.A3(n_26),
.B1(n_25),
.B2(n_229),
.Y(n_384)
);

XOR2x2_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_323),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_300),
.A2(n_176),
.B1(n_2),
.B2(n_3),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_311),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_389),
.A2(n_311),
.B1(n_305),
.B2(n_320),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_317),
.B(n_4),
.C(n_5),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_303),
.B(n_5),
.C(n_6),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_393),
.C(n_307),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_335),
.B(n_6),
.C(n_7),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_354),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_395),
.B(n_396),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_324),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_354),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_397),
.B(n_404),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_419),
.Y(n_437)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_380),
.Y(n_400)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_401),
.Y(n_440)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_386),
.Y(n_403)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_376),
.Y(n_404)
);

AO21x2_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_308),
.B(n_323),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_405),
.A2(n_409),
.B1(n_378),
.B2(n_357),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_362),
.A2(n_308),
.B1(n_319),
.B2(n_316),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_406),
.A2(n_361),
.B1(n_363),
.B2(n_356),
.Y(n_443)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_408),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_351),
.A2(n_341),
.B(n_298),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_411),
.A2(n_415),
.B(n_383),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_342),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_414),
.Y(n_441)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_360),
.B(n_348),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_364),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_421),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_321),
.Y(n_417)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_315),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_423),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_307),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_429),
.Y(n_444)
);

BUFx12_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_426),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_375),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_382),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_353),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_355),
.B(n_337),
.C(n_322),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_432),
.B(n_381),
.C(n_373),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_359),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_436),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_371),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_443),
.A2(n_460),
.B1(n_464),
.B2(n_430),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_447),
.A2(n_467),
.B(n_402),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_468),
.C(n_418),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_423),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_450),
.B(n_451),
.Y(n_485)
);

NOR4xp25_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_368),
.C(n_357),
.D(n_394),
.Y(n_451)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_426),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_456),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_352),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_434),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_405),
.A2(n_374),
.B1(n_393),
.B2(n_387),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_458),
.A2(n_462),
.B1(n_415),
.B2(n_420),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_426),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_400),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_388),
.B1(n_392),
.B2(n_370),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_415),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_427),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_405),
.A2(n_375),
.B1(n_394),
.B2(n_358),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_406),
.A2(n_379),
.B1(n_390),
.B2(n_365),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_384),
.Y(n_466)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_418),
.B(n_299),
.C(n_365),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_470),
.A2(n_473),
.B1(n_483),
.B2(n_386),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_405),
.B1(n_410),
.B2(n_402),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_471),
.A2(n_479),
.B1(n_480),
.B2(n_493),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_445),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_472),
.B(n_491),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_441),
.B(n_401),
.Y(n_474)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_474),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_476),
.B(n_482),
.C(n_487),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_467),
.A2(n_411),
.B(n_427),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_478),
.A2(n_466),
.B(n_461),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_463),
.A2(n_405),
.B1(n_410),
.B2(n_399),
.Y(n_479)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_399),
.C(n_425),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_462),
.A2(n_429),
.B1(n_419),
.B2(n_424),
.Y(n_483)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_486),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_428),
.C(n_398),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_329),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_488),
.B(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_490),
.Y(n_510)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_436),
.B(n_413),
.C(n_409),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_492),
.B(n_465),
.C(n_440),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_443),
.A2(n_407),
.B1(n_424),
.B2(n_403),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_439),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_494),
.A2(n_457),
.B1(n_455),
.B2(n_465),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_446),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_437),
.A2(n_407),
.B1(n_391),
.B2(n_379),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_496),
.A2(n_457),
.B1(n_455),
.B2(n_449),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_454),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_498),
.B(n_501),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_437),
.Y(n_501)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_452),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_507),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_458),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_511),
.B(n_513),
.C(n_517),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_512),
.A2(n_349),
.B(n_338),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_489),
.B(n_435),
.C(n_444),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_444),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_515),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_438),
.Y(n_515)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_489),
.B(n_440),
.C(n_464),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_460),
.C(n_449),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_517),
.C(n_513),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_469),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_519),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_474),
.Y(n_520)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_521),
.A2(n_490),
.B1(n_486),
.B2(n_483),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_522),
.A2(n_480),
.B1(n_471),
.B2(n_479),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_500),
.A2(n_485),
.B(n_477),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_532),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_481),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_503),
.A2(n_470),
.B1(n_484),
.B2(n_473),
.Y(n_527)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_527),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_528),
.B(n_541),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_529),
.B(n_514),
.Y(n_552)
);

A2O1A1O1Ixp25_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_484),
.B(n_478),
.C(n_491),
.D(n_494),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_530),
.A2(n_510),
.B(n_506),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_493),
.B1(n_496),
.B2(n_472),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_508),
.B(n_344),
.C(n_334),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_539),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g537 ( 
.A1(n_502),
.A2(n_386),
.B(n_301),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_521),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_538),
.B(n_509),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_508),
.B(n_346),
.C(n_340),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_314),
.C(n_7),
.Y(n_541)
);

FAx1_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_518),
.CI(n_501),
.CON(n_543),
.SN(n_543)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_543),
.A2(n_524),
.B(n_530),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_544),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_545),
.B(n_525),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_528),
.C(n_539),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_547),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_507),
.C(n_515),
.Y(n_547)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_551),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_552),
.B(n_535),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_499),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_553),
.A2(n_556),
.B(n_524),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_498),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_554),
.B(n_6),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_505),
.Y(n_556)
);

OAI321xp33_ASAP7_75t_L g557 ( 
.A1(n_536),
.A2(n_15),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C(n_13),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_557),
.A2(n_532),
.B1(n_529),
.B2(n_541),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_562),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g561 ( 
.A1(n_548),
.A2(n_533),
.B(n_534),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_563),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_531),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_567),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_571),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_546),
.B(n_531),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_555),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_569),
.B(n_549),
.C(n_559),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_572),
.B(n_578),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_579),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_570),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_550),
.Y(n_579)
);

AOI322xp5_ASAP7_75t_L g580 ( 
.A1(n_575),
.A2(n_550),
.A3(n_566),
.B1(n_558),
.B2(n_563),
.C1(n_560),
.C2(n_543),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_580),
.B(n_581),
.Y(n_585)
);

MAJx2_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_548),
.C(n_562),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_572),
.B(n_568),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_583),
.B(n_576),
.Y(n_586)
);

AO21x1_ASAP7_75t_L g589 ( 
.A1(n_586),
.A2(n_587),
.B(n_8),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_584),
.A2(n_573),
.B1(n_551),
.B2(n_574),
.Y(n_587)
);

AOI322xp5_ASAP7_75t_L g588 ( 
.A1(n_585),
.A2(n_582),
.A3(n_543),
.B1(n_571),
.B2(n_554),
.C1(n_8),
.C2(n_14),
.Y(n_588)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_588),
.B(n_589),
.C(n_8),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_587),
.B1(n_11),
.B2(n_14),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_591),
.A2(n_10),
.B(n_14),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_592),
.A2(n_10),
.B(n_15),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_15),
.Y(n_594)
);


endmodule