module fake_jpeg_13449_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_12),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_8),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_95),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_64),
.Y(n_203)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_28),
.B1(n_42),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_67),
.A2(n_109),
.B1(n_128),
.B2(n_29),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_83),
.Y(n_184)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_84),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_19),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_57),
.Y(n_130)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_88),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_89),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_31),
.B(n_9),
.Y(n_95)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_31),
.Y(n_96)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_26),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_52),
.Y(n_145)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_103),
.Y(n_185)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_104),
.Y(n_206)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_26),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_119),
.B(n_25),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_27),
.Y(n_120)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_27),
.Y(n_124)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_127),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_35),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_130),
.B(n_131),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_57),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_59),
.A2(n_56),
.B1(n_53),
.B2(n_52),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_134),
.A2(n_154),
.B1(n_158),
.B2(n_195),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_135),
.A2(n_178),
.B1(n_179),
.B2(n_208),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_58),
.B(n_48),
.C(n_49),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g295 ( 
.A1(n_136),
.A2(n_219),
.B1(n_2),
.B2(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_56),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_143),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_53),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_145),
.B(n_153),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_151),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_37),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_43),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_80),
.A2(n_47),
.B1(n_40),
.B2(n_21),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_43),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_155),
.B(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_21),
.B1(n_49),
.B2(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_51),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_160),
.B(n_174),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_71),
.B(n_51),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_85),
.A2(n_49),
.B1(n_21),
.B2(n_30),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_86),
.A2(n_33),
.B1(n_30),
.B2(n_38),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_93),
.A2(n_40),
.B(n_47),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_104),
.A2(n_47),
.B1(n_40),
.B2(n_33),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_76),
.B(n_38),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_211),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_123),
.B(n_33),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_91),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_63),
.A2(n_29),
.B1(n_35),
.B2(n_25),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_106),
.A2(n_110),
.B1(n_129),
.B2(n_111),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_126),
.B1(n_125),
.B2(n_77),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_112),
.B(n_29),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_64),
.B(n_17),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_2),
.Y(n_285)
);

HAxp5_ASAP7_75t_SL g219 ( 
.A(n_70),
.B(n_25),
.CON(n_219),
.SN(n_219)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_187),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_223),
.B(n_238),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_136),
.A2(n_66),
.B1(n_68),
.B2(n_74),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_224),
.A2(n_258),
.B1(n_270),
.B2(n_173),
.Y(n_309)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_227),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_140),
.B(n_0),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_297),
.Y(n_302)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_229),
.Y(n_352)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_231),
.Y(n_321)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_233),
.Y(n_328)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx8_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_145),
.B(n_107),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_240),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_187),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_241),
.A2(n_261),
.B1(n_278),
.B2(n_281),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_152),
.B(n_98),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_134),
.A2(n_155),
.B1(n_140),
.B2(n_75),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_247),
.A2(n_198),
.B1(n_180),
.B2(n_183),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_248),
.B(n_257),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_156),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_249),
.B(n_254),
.Y(n_338)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_159),
.B(n_89),
.Y(n_254)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_255),
.Y(n_342)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

INVx4_ASAP7_75t_SL g257 ( 
.A(n_219),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_209),
.A2(n_17),
.B1(n_15),
.B2(n_14),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_203),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_262),
.B(n_263),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_161),
.B(n_162),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_265),
.B(n_266),
.Y(n_349)
);

INVx4_ASAP7_75t_SL g266 ( 
.A(n_185),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVx11_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_268),
.Y(n_341)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_163),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_269),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_184),
.Y(n_271)
);

INVx13_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_273),
.Y(n_332)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_274),
.Y(n_354)
);

INVx6_ASAP7_75t_SL g275 ( 
.A(n_185),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_275),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_193),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_276),
.B(n_282),
.Y(n_323)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_164),
.B(n_1),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_286),
.C(n_290),
.Y(n_312)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_196),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_284),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_285),
.B(n_292),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_172),
.B(n_17),
.C(n_15),
.Y(n_286)
);

INVx11_ASAP7_75t_L g287 ( 
.A(n_137),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_214),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_165),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g290 ( 
.A(n_188),
.B(n_2),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_169),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_213),
.Y(n_294)
);

AO22x1_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_169),
.B1(n_186),
.B2(n_182),
.Y(n_343)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_201),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_132),
.B(n_11),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_216),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_147),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_195),
.B1(n_194),
.B2(n_173),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_303),
.A2(n_325),
.B1(n_275),
.B2(n_248),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g367 ( 
.A1(n_309),
.A2(n_310),
.B1(n_358),
.B2(n_326),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_234),
.A2(n_167),
.B1(n_166),
.B2(n_144),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_232),
.A2(n_142),
.B(n_171),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_294),
.B(n_298),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_202),
.C(n_191),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_351),
.C(n_357),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_167),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_350),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_279),
.A2(n_168),
.B1(n_199),
.B2(n_215),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_277),
.A2(n_183),
.B1(n_148),
.B2(n_166),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_326),
.A2(n_359),
.B1(n_261),
.B2(n_227),
.Y(n_381)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_237),
.B(n_199),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_333),
.B(n_266),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_344),
.B1(n_345),
.B2(n_253),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_343),
.A2(n_229),
.B(n_6),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_279),
.A2(n_148),
.B1(n_144),
.B2(n_198),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_234),
.A2(n_180),
.B1(n_215),
.B2(n_182),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_186),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_259),
.B(n_3),
.C(n_4),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_228),
.B(n_3),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_232),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_230),
.B(n_6),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_286),
.C(n_251),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_345),
.A2(n_270),
.B1(n_271),
.B2(n_257),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

OAI21xp33_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_232),
.B(n_245),
.Y(n_363)
);

OAI21xp33_ASAP7_75t_SL g425 ( 
.A1(n_363),
.A2(n_367),
.B(n_358),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_364),
.A2(n_371),
.B(n_375),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_323),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_388),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_312),
.B(n_248),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_374),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_368),
.Y(n_432)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_344),
.A2(n_295),
.B1(n_280),
.B2(n_264),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_373),
.B1(n_376),
.B2(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_333),
.A2(n_280),
.B1(n_264),
.B2(n_283),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_334),
.A2(n_260),
.B(n_284),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_333),
.A2(n_291),
.B1(n_281),
.B2(n_265),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_378),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_312),
.B(n_226),
.C(n_299),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_379),
.B(n_380),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_250),
.C(n_272),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_341),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_309),
.A2(n_236),
.B1(n_255),
.B2(n_243),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_246),
.C(n_231),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_383),
.B(n_387),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_316),
.A2(n_235),
.B1(n_274),
.B2(n_256),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_386),
.A2(n_407),
.B(n_324),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_287),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_233),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_307),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_390),
.Y(n_430)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_314),
.A2(n_289),
.B(n_267),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_391),
.A2(n_349),
.B(n_354),
.Y(n_431)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_392),
.B(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_399),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_278),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_397),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_244),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_302),
.B(n_268),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_402),
.C(n_403),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_225),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_304),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_339),
.A2(n_6),
.B1(n_7),
.B2(n_322),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_302),
.B(n_6),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_7),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_320),
.A2(n_7),
.B1(n_343),
.B2(n_315),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_404),
.A2(n_354),
.B1(n_330),
.B2(n_313),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_320),
.B(n_318),
.C(n_331),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_405),
.B(n_406),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_323),
.B(n_351),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_343),
.A2(n_349),
.B1(n_335),
.B2(n_341),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_SL g462 ( 
.A1(n_412),
.A2(n_376),
.B1(n_401),
.B2(n_367),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_370),
.A2(n_359),
.B1(n_340),
.B2(n_306),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_414),
.A2(n_418),
.B1(n_421),
.B2(n_424),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_396),
.B(n_332),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_420),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_364),
.A2(n_407),
.B1(n_394),
.B2(n_392),
.Y(n_418)
);

AO22x1_ASAP7_75t_SL g420 ( 
.A1(n_400),
.A2(n_329),
.B1(n_327),
.B2(n_324),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_368),
.A2(n_332),
.B1(n_306),
.B2(n_346),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_397),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_436),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_423),
.B(n_431),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_342),
.B1(n_337),
.B2(n_317),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_425),
.A2(n_386),
.B(n_395),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_337),
.B1(n_342),
.B2(n_317),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_427),
.A2(n_437),
.B1(n_442),
.B2(n_445),
.Y(n_468)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_386),
.B(n_404),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_440),
.B(n_371),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_406),
.B(n_330),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_381),
.A2(n_336),
.B1(n_313),
.B2(n_348),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_375),
.A2(n_348),
.B(n_321),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_393),
.A2(n_336),
.B1(n_329),
.B2(n_327),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_431),
.B(n_411),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_373),
.A2(n_321),
.B1(n_319),
.B2(n_353),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_447),
.A2(n_452),
.B(n_481),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_430),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_456),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_429),
.B(n_366),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g510 ( 
.A(n_451),
.B(n_469),
.Y(n_510)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_379),
.C(n_387),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_460),
.C(n_477),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_430),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_433),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_463),
.Y(n_496)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_439),
.B(n_398),
.C(n_361),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_461),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_462),
.A2(n_476),
.B1(n_426),
.B2(n_424),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_417),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_391),
.B(n_399),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_464),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_465),
.B(n_466),
.Y(n_507)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_428),
.B(n_361),
.CI(n_374),
.CON(n_466),
.SN(n_466)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_419),
.B(n_405),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_408),
.B(n_352),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_446),
.C(n_301),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_416),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_472),
.Y(n_512)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_441),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_475),
.Y(n_505)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_432),
.A2(n_367),
.B1(n_380),
.B2(n_383),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_403),
.C(n_402),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_478),
.A2(n_434),
.B(n_410),
.Y(n_485)
);

OA22x2_ASAP7_75t_L g479 ( 
.A1(n_422),
.A2(n_367),
.B1(n_377),
.B2(n_378),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_479),
.B(n_480),
.Y(n_509)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_423),
.A2(n_384),
.B(n_328),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_419),
.B(n_304),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_440),
.C(n_444),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_415),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_484),
.B(n_489),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_485),
.A2(n_481),
.B(n_479),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_457),
.A2(n_418),
.B1(n_414),
.B2(n_421),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_486),
.A2(n_493),
.B1(n_502),
.B2(n_514),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_415),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_472),
.A2(n_432),
.B1(n_412),
.B2(n_437),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_491),
.A2(n_495),
.B1(n_511),
.B2(n_468),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_436),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_494),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_443),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_459),
.A2(n_443),
.B1(n_427),
.B2(n_428),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_500),
.C(n_503),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_435),
.C(n_409),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_450),
.A2(n_411),
.B1(n_426),
.B2(n_445),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_435),
.C(n_409),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_435),
.C(n_442),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_449),
.C(n_476),
.Y(n_525)
);

XOR2x1_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_434),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_506),
.B(n_455),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_516),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_459),
.A2(n_420),
.B1(n_353),
.B2(n_328),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_450),
.A2(n_420),
.B1(n_319),
.B2(n_301),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_467),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_456),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_517),
.B(n_529),
.Y(n_546)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_520),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_478),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_521),
.B(n_522),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_452),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_525),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_455),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_528),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_505),
.Y(n_527)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_527),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_489),
.B(n_466),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_488),
.B(n_448),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_507),
.B(n_496),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_530),
.B(n_448),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_447),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_533),
.C(n_537),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_470),
.C(n_464),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_534),
.A2(n_483),
.B1(n_499),
.B2(n_461),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_463),
.Y(n_535)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_535),
.Y(n_563)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_505),
.Y(n_536)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_536),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_510),
.B(n_470),
.C(n_479),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_510),
.B(n_479),
.C(n_420),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_539),
.C(n_540),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_500),
.B(n_479),
.C(n_480),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_503),
.C(n_498),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_544),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_475),
.C(n_474),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_497),
.C(n_485),
.Y(n_564)
);

XOR2x2_ASAP7_75t_L g544 ( 
.A(n_513),
.B(n_458),
.Y(n_544)
);

FAx1_ASAP7_75t_SL g545 ( 
.A(n_506),
.B(n_468),
.CI(n_453),
.CON(n_545),
.SN(n_545)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_545),
.A2(n_538),
.B1(n_486),
.B2(n_537),
.Y(n_551)
);

CKINVDCx14_ASAP7_75t_R g578 ( 
.A(n_547),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_533),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_541),
.A2(n_493),
.B1(n_502),
.B2(n_501),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_553),
.A2(n_556),
.B1(n_566),
.B2(n_569),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_543),
.A2(n_509),
.B1(n_511),
.B2(n_513),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_554),
.A2(n_557),
.B1(n_545),
.B2(n_490),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_539),
.A2(n_514),
.B1(n_509),
.B2(n_515),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_527),
.A2(n_509),
.B1(n_497),
.B2(n_505),
.Y(n_557)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_542),
.Y(n_559)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_559),
.Y(n_577)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_560),
.Y(n_587)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_561),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_564),
.B(n_532),
.Y(n_571)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_544),
.Y(n_568)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_568),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_525),
.A2(n_473),
.B1(n_490),
.B2(n_301),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_560),
.Y(n_570)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_570),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_571),
.B(n_581),
.Y(n_590)
);

XNOR2x1_ASAP7_75t_L g604 ( 
.A(n_572),
.B(n_580),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_558),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_585),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_550),
.B(n_526),
.C(n_559),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_575),
.B(n_583),
.Y(n_597)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_546),
.A2(n_522),
.B(n_521),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_582),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_554),
.A2(n_545),
.B1(n_523),
.B2(n_540),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_562),
.B(n_518),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_518),
.C(n_523),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_528),
.B1(n_519),
.B2(n_355),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_552),
.A2(n_519),
.B(n_355),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_548),
.B(n_562),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_553),
.A2(n_355),
.B1(n_556),
.B2(n_565),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_588),
.B(n_569),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_575),
.B(n_549),
.C(n_555),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_595),
.C(n_596),
.Y(n_606)
);

INVx11_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_592),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_580),
.A2(n_568),
.B(n_561),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_593),
.A2(n_599),
.B(n_603),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_549),
.C(n_555),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_567),
.C(n_564),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_576),
.A2(n_558),
.B(n_563),
.Y(n_599)
);

AOI22x1_ASAP7_75t_L g610 ( 
.A1(n_600),
.A2(n_573),
.B1(n_574),
.B2(n_581),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_584),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_557),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_584),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_576),
.A2(n_567),
.B(n_588),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_597),
.B(n_587),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_608),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_591),
.B(n_595),
.C(n_597),
.Y(n_608)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_609),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_610),
.B(n_613),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_593),
.A2(n_574),
.B(n_586),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_612),
.B(n_614),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_590),
.A2(n_585),
.B(n_572),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_596),
.B(n_582),
.C(n_604),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_598),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_604),
.B(n_601),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_616),
.B(n_617),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_590),
.B(n_592),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_606),
.B(n_603),
.C(n_602),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_624),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_608),
.A2(n_589),
.B(n_594),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_611),
.A2(n_609),
.B(n_606),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_626),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_589),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_627),
.B(n_599),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_628),
.A2(n_633),
.B(n_634),
.Y(n_635)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_612),
.C(n_594),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_625),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_632),
.A2(n_618),
.B(n_621),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_623),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_622),
.A2(n_615),
.B(n_611),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_629),
.A2(n_622),
.B(n_620),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_636),
.Y(n_640)
);

AO21x1_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_638),
.B(n_630),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_639),
.A2(n_635),
.B(n_610),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_641),
.B(n_640),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_SL g643 ( 
.A1(n_642),
.A2(n_616),
.B1(n_613),
.B2(n_598),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_600),
.Y(n_644)
);


endmodule