module real_jpeg_1867_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_148)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_68),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_68),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_4),
.B(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_40),
.C(n_55),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_4),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_4),
.B(n_54),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_27),
.C(n_45),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_33),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_50),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_168),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_69),
.B1(n_71),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_82),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_82),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_82),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_49),
.B1(n_58),
.B2(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_69),
.B1(n_71),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_12),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_129),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_129),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_14),
.A2(n_62),
.B1(n_69),
.B2(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_14),
.A2(n_40),
.B1(n_42),
.B2(n_62),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_62),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_16),
.A2(n_30),
.B1(n_40),
.B2(n_42),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_131),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_110),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.C(n_65),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_22),
.A2(n_23),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_24),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_26),
.A2(n_33),
.B1(n_98),
.B2(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_32),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_27),
.B(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_31),
.A2(n_32),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_31),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_31),
.A2(n_32),
.B1(n_148),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_31),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_31),
.A2(n_32),
.B1(n_193),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_32),
.A2(n_147),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_32),
.B(n_162),
.Y(n_195)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_33),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_33),
.A2(n_161),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_38),
.A2(n_43),
.B1(n_50),
.B2(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_40),
.B(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_43),
.A2(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_43),
.B(n_154),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_47),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_47),
.A2(n_175),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_47),
.A2(n_87),
.B1(n_151),
.B2(n_201),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_50),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_51),
.B(n_65),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_52),
.A2(n_63),
.B1(n_64),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_52),
.A2(n_63),
.B1(n_141),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_52),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_52),
.A2(n_172),
.B(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_53),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_54),
.B(n_126),
.Y(n_234)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_58),
.B(n_158),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_58),
.B(n_76),
.Y(n_182)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI32xp33_ASAP7_75t_L g180 ( 
.A1(n_59),
.A2(n_69),
.A3(n_75),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_61),
.A2(n_63),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_63),
.A2(n_125),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_72),
.B(n_79),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_73),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_69),
.A2(n_72),
.B(n_168),
.C(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_69),
.B(n_168),
.Y(n_169)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_74),
.A2(n_103),
.B(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_80),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_92),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_90),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_87),
.A2(n_153),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_106),
.B2(n_109),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_105),
.B1(n_107),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_98),
.A2(n_168),
.B(n_195),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_116),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_111),
.B(n_114),
.Y(n_279)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_116),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.C(n_127),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_117),
.A2(n_118),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_119),
.B(n_121),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_120),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_276),
.B(n_280),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_245),
.B(n_273),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_187),
.B(n_244),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_138),
.B(n_163),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.C(n_155),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_139),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_149),
.B(n_155),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_164),
.B(n_178),
.C(n_186),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_176),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_165),
.B(n_171),
.C(n_173),
.Y(n_258)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_179),
.B(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_239),
.B(n_243),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_228),
.B(n_238),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_210),
.B(n_227),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_204),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_204),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_196),
.B1(n_202),
.B2(n_203),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_199),
.C(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_221),
.B(n_226),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_216),
.B(n_220),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_219),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_224),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_230),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_259),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_259),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_257),
.C(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_251),
.C(n_255),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_272),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_266),
.C(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);


endmodule