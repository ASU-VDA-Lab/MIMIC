module real_jpeg_15912_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_11;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_1),
.A2(n_31),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_146),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_5),
.A2(n_104),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_7),
.A2(n_15),
.B1(n_33),
.B2(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_7),
.B(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_137),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_111),
.B(n_136),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_48),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_13),
.B(n_48),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_21),
.B1(n_32),
.B2(n_37),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_15),
.A2(n_22),
.B1(n_124),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_38),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_18),
.Y(n_143)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_20),
.Y(n_125)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_20),
.Y(n_128)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_20),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_41),
.Y(n_153)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_73),
.B1(n_109),
.B2(n_110),
.Y(n_48)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_49),
.B(n_110),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.A3(n_55),
.B1(n_58),
.B2(n_65),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_52),
.A2(n_79),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_90),
.B1(n_94),
.B2(n_97),
.Y(n_89)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_59),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_59),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_80),
.B1(n_98),
.B2(n_107),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_80),
.A2(n_98),
.B1(n_107),
.B2(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_129),
.B(n_135),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_134),
.Y(n_135)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_173),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_141),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_154),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_162),
.B1(n_163),
.B2(n_172),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);


endmodule