module fake_jpeg_23663_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_18),
.A2(n_1),
.B(n_2),
.Y(n_34)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_5),
.CI(n_6),
.CON(n_69),
.SN(n_69)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_40),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_2),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_42),
.C(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_3),
.B(n_4),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_4),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_47),
.B1(n_23),
.B2(n_17),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_16),
.B1(n_20),
.B2(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_15),
.B1(n_20),
.B2(n_24),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_57),
.B1(n_64),
.B2(n_69),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_23),
.B1(n_25),
.B2(n_19),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_71),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_91),
.B1(n_92),
.B2(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_77),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_56),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_82),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_79),
.B(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_33),
.B1(n_43),
.B2(n_39),
.Y(n_86)
);

AO22x1_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_65),
.B1(n_62),
.B2(n_50),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_17),
.B1(n_19),
.B2(n_30),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_36),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_32),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_61),
.C(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_30),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_27),
.B1(n_22),
.B2(n_7),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_68),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_106),
.B1(n_108),
.B2(n_97),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_68),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_111),
.B(n_89),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_90),
.B1(n_83),
.B2(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_110),
.B1(n_86),
.B2(n_71),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_54),
.C(n_51),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_79),
.B(n_78),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_45),
.B1(n_50),
.B2(n_27),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_27),
.B(n_22),
.C(n_8),
.D(n_9),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_86),
.A3(n_87),
.B1(n_81),
.B2(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_100),
.A2(n_72),
.B1(n_86),
.B2(n_75),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_125),
.B1(n_126),
.B2(n_99),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NOR4xp25_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_124),
.C(n_109),
.D(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_86),
.B1(n_89),
.B2(n_75),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_120),
.B(n_123),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_135),
.B1(n_114),
.B2(n_124),
.C(n_112),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_95),
.C(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_110),
.C(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_94),
.B1(n_93),
.B2(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_77),
.C(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_82),
.C(n_99),
.Y(n_134)
);

OAI21x1_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_123),
.B(n_113),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_27),
.CI(n_22),
.CON(n_145),
.SN(n_145)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_126),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_143),
.B1(n_145),
.B2(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_116),
.B(n_118),
.C(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_137),
.B1(n_131),
.B2(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_104),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_139),
.C(n_146),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_140),
.A3(n_146),
.B1(n_139),
.B2(n_144),
.C1(n_145),
.C2(n_104),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_156),
.C(n_150),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_144),
.B(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_12),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_10),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_154),
.B1(n_8),
.B2(n_9),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_5),
.C(n_8),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.Y(n_164)
);


endmodule