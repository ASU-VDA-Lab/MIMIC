module real_jpeg_13525_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_43),
.B1(n_59),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_2),
.A2(n_29),
.B1(n_37),
.B2(n_43),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_29),
.B1(n_37),
.B2(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_53),
.B1(n_59),
.B2(n_62),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_29),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_120)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_7),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_7),
.A2(n_29),
.B1(n_37),
.B2(n_68),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_9),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_64),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_9),
.B(n_112),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_62),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_99),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_45),
.B(n_49),
.C(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_9),
.B(n_105),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_33),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_85),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_62),
.B(n_178),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_64),
.B1(n_65),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_10),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_10),
.A2(n_59),
.B1(n_62),
.B2(n_109),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_109),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_29),
.B1(n_37),
.B2(n_109),
.Y(n_214)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_59),
.B1(n_62),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_78),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_29),
.B1(n_37),
.B2(n_78),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_13),
.A2(n_29),
.B1(n_37),
.B2(n_70),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_15),
.A2(n_29),
.B1(n_37),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_15),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_16),
.A2(n_36),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_131),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_113),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_21),
.B(n_113),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_22),
.A2(n_23),
.B1(n_80),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_54),
.B2(n_55),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_56),
.C(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_26),
.B(n_40),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_27),
.A2(n_32),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_28),
.A2(n_33),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_28),
.A2(n_33),
.B(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_28),
.A2(n_33),
.B1(n_95),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_33),
.B1(n_157),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_28),
.A2(n_33),
.B1(n_181),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_28),
.A2(n_33),
.B1(n_99),
.B2(n_214),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_28),
.A2(n_33),
.B1(n_207),
.B2(n_214),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_29),
.B(n_216),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_37),
.A2(n_50),
.B(n_99),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_42),
.A2(n_47),
.B1(n_85),
.B2(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_45),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_44),
.A2(n_62),
.A3(n_75),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_45),
.B(n_74),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_46),
.A2(n_51),
.B1(n_172),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_47),
.A2(n_84),
.B1(n_85),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_47),
.A2(n_85),
.B1(n_145),
.B2(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_47),
.A2(n_85),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_47),
.A2(n_85),
.B1(n_193),
.B2(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_71),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_69),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_57),
.A2(n_58),
.B1(n_108),
.B2(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_62),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_61),
.A3(n_64),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_62),
.Y(n_97)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_65),
.B(n_99),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_73),
.B1(n_79),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_72),
.A2(n_73),
.B1(n_102),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_72),
.A2(n_73),
.B1(n_153),
.B2(n_228),
.Y(n_227)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_73),
.Y(n_105)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_80),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_90),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_91),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.C(n_106),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_98),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_100),
.B(n_106),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_103),
.A2(n_105),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_119),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_164),
.B(n_242),
.C(n_247),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_158),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_135),
.B(n_158),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.C(n_150),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_136),
.A2(n_137),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_142),
.C(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_148),
.B(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_156),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_241),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_185),
.B(n_240),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_182),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_167),
.B(n_182),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_173),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_168),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_170),
.A2(n_173),
.B1(n_174),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_234),
.B(n_239),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_223),
.B(n_233),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_203),
.B(n_222),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_189),
.B(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_211),
.B(n_221),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_209),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_217),
.B(n_220),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_225),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_229),
.C(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);


endmodule