module fake_jpeg_14899_n_90 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_1),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_52),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_20),
.B1(n_32),
.B2(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_35),
.B1(n_6),
.B2(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_2),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_35),
.B1(n_40),
.B2(n_38),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_42),
.B1(n_45),
.B2(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_3),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.C(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_72),
.B1(n_11),
.B2(n_17),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_10),
.B(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_21),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_83),
.A2(n_82),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_27),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g89 ( 
.A(n_88),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_28),
.B(n_30),
.Y(n_90)
);


endmodule