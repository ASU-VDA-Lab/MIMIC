module fake_aes_10467_n_25 (n_1, n_2, n_4, n_3, n_5, n_0, n_25);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
AOI21x1_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_4), .B(n_5), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
OAI22x1_ASAP7_75t_L g8 ( .A1(n_1), .A2(n_2), .B1(n_4), .B2(n_3), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_0), .B(n_2), .Y(n_9) );
INVx5_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
BUFx4f_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
AOI21x1_ASAP7_75t_L g14 ( .A1(n_6), .A2(n_9), .B(n_8), .Y(n_14) );
INVx2_ASAP7_75t_SL g15 ( .A(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_11), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_15), .B(n_12), .Y(n_19) );
OAI221xp5_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_17), .B1(n_16), .B2(n_8), .C(n_14), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_18), .B(n_16), .Y(n_21) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_21), .B(n_10), .Y(n_22) );
AND2x2_ASAP7_75t_SL g23 ( .A(n_20), .B(n_10), .Y(n_23) );
OAI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_10), .B(n_22), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_24), .B(n_23), .Y(n_25) );
endmodule