module fake_jpeg_29978_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_0),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_32),
.B2(n_21),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_22),
.B1(n_21),
.B2(n_32),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_42),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

OR2x4_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_43),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_80),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_35),
.C(n_40),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_75),
.Y(n_110)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_34),
.B1(n_30),
.B2(n_18),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_58),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_30),
.B(n_27),
.Y(n_81)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_81),
.B(n_24),
.CI(n_33),
.CON(n_115),
.SN(n_115)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_63),
.B(n_19),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_16),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_10),
.B(n_13),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_119),
.B(n_103),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_33),
.B1(n_82),
.B2(n_68),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_29),
.B1(n_30),
.B2(n_25),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_111),
.B1(n_121),
.B2(n_73),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_26),
.B1(n_23),
.B2(n_27),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_118),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_87),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_71),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_132),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_80),
.B(n_86),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_129),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_84),
.C(n_86),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_130),
.C(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_23),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_135),
.Y(n_153)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

OR2x4_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_20),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_83),
.C(n_78),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_26),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_74),
.B1(n_78),
.B2(n_83),
.Y(n_136)
);

AO22x2_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_113),
.B1(n_101),
.B2(n_114),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_144),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_73),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_100),
.A2(n_67),
.B1(n_66),
.B2(n_4),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_123),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_67),
.B1(n_66),
.B2(n_4),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_158),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_100),
.C(n_115),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_130),
.C(n_122),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_112),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_143),
.B1(n_162),
.B2(n_158),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_125),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_145),
.C(n_151),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_171),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_141),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_169),
.B(n_170),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_129),
.C(n_106),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_147),
.B1(n_131),
.B2(n_146),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_182),
.C(n_183),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_181),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_163),
.C(n_131),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_148),
.B1(n_160),
.B2(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_185),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_163),
.B1(n_162),
.B2(n_108),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_142),
.B1(n_157),
.B2(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_107),
.B1(n_15),
.B2(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_2),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_174),
.A3(n_165),
.B1(n_175),
.B2(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_199),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_182),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_206),
.B1(n_107),
.B2(n_12),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_178),
.C(n_186),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_206),
.A2(n_197),
.B(n_193),
.C(n_107),
.Y(n_207)
);

AOI21x1_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_204),
.B(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_208),
.B(n_211),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_11),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C1(n_8),
.C2(n_2),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_213),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_3),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_207),
.C(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_3),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_8),
.C(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_8),
.Y(n_220)
);


endmodule