module fake_jpeg_22887_n_39 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx11_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_23),
.B1(n_19),
.B2(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_9),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.C(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_23),
.C(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_13),
.B2(n_15),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_10),
.CI(n_16),
.CON(n_38),
.SN(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_17),
.Y(n_39)
);


endmodule