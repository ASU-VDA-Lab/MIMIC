module real_aes_6725_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g165 ( .A1(n_0), .A2(n_166), .B(n_169), .C(n_173), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_1), .B(n_157), .Y(n_176) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_3), .B(n_167), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_4), .A2(n_130), .B(n_133), .C(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_5), .A2(n_125), .B(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_6), .A2(n_125), .B(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_7), .B(n_157), .Y(n_528) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_8), .A2(n_159), .B(n_231), .Y(n_230) );
AND2x6_ASAP7_75t_L g130 ( .A(n_9), .B(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_10), .A2(n_130), .B(n_133), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g488 ( .A(n_11), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_12), .B(n_39), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_13), .B(n_172), .Y(n_499) );
INVx1_ASAP7_75t_L g151 ( .A(n_14), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_15), .B(n_167), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_16), .A2(n_168), .B(n_508), .C(n_510), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_17), .B(n_157), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_18), .B(n_145), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_19), .A2(n_133), .B(n_136), .C(n_144), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_20), .A2(n_171), .B(n_239), .C(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_21), .B(n_172), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_22), .B(n_172), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_23), .Y(n_469) );
INVx1_ASAP7_75t_L g449 ( .A(n_24), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_25), .A2(n_133), .B(n_144), .C(n_234), .Y(n_233) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_26), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_27), .Y(n_495) );
INVx1_ASAP7_75t_L g463 ( .A(n_28), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_29), .A2(n_125), .B(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g128 ( .A(n_30), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_31), .A2(n_183), .B(n_184), .C(n_188), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_32), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_33), .A2(n_103), .B1(n_736), .B2(n_745), .C(n_749), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_33), .A2(n_754), .B1(n_759), .B2(n_760), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_33), .Y(n_759) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_34), .A2(n_171), .B(n_525), .C(n_527), .Y(n_524) );
INVxp67_ASAP7_75t_L g464 ( .A(n_35), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_36), .B(n_236), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_37), .A2(n_133), .B(n_144), .C(n_448), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g523 ( .A(n_38), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_40), .A2(n_173), .B(n_486), .C(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_41), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g252 ( .A(n_42), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_43), .B(n_167), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_44), .B(n_125), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_45), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_46), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_47), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_48), .A2(n_183), .B(n_188), .C(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g170 ( .A(n_49), .Y(n_170) );
INVx1_ASAP7_75t_L g214 ( .A(n_50), .Y(n_214) );
INVx1_ASAP7_75t_L g536 ( .A(n_51), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_52), .B(n_125), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_53), .Y(n_153) );
CKINVDCx14_ASAP7_75t_R g484 ( .A(n_54), .Y(n_484) );
INVx1_ASAP7_75t_L g131 ( .A(n_55), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_56), .B(n_125), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_57), .B(n_157), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_58), .A2(n_143), .B(n_199), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
INVx1_ASAP7_75t_SL g526 ( .A(n_60), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_61), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_62), .B(n_167), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_63), .B(n_157), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_64), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_65), .B(n_168), .Y(n_249) );
INVx1_ASAP7_75t_L g472 ( .A(n_66), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_67), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_68), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_69), .A2(n_133), .B(n_188), .C(n_197), .Y(n_196) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_70), .Y(n_223) );
INVx1_ASAP7_75t_L g740 ( .A(n_71), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_72), .A2(n_125), .B(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_73), .A2(n_94), .B1(n_757), .B2(n_758), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_73), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_74), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_75), .A2(n_125), .B(n_505), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_76), .A2(n_101), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_76), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_77), .A2(n_124), .B(n_459), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_78), .Y(n_446) );
INVx1_ASAP7_75t_L g506 ( .A(n_79), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_80), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_80), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_81), .B(n_141), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_82), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_83), .A2(n_125), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g509 ( .A(n_84), .Y(n_509) );
INVx2_ASAP7_75t_L g148 ( .A(n_85), .Y(n_148) );
INVx1_ASAP7_75t_L g498 ( .A(n_86), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_87), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_88), .B(n_172), .Y(n_250) );
OR2x2_ASAP7_75t_L g108 ( .A(n_89), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g438 ( .A(n_89), .Y(n_438) );
OR2x2_ASAP7_75t_L g744 ( .A(n_89), .B(n_734), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_90), .A2(n_133), .B(n_188), .C(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_91), .B(n_125), .Y(n_181) );
INVx1_ASAP7_75t_L g185 ( .A(n_92), .Y(n_185) );
INVxp67_ASAP7_75t_L g226 ( .A(n_93), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_94), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_95), .B(n_159), .Y(n_489) );
INVx1_ASAP7_75t_L g198 ( .A(n_96), .Y(n_198) );
INVx1_ASAP7_75t_L g245 ( .A(n_97), .Y(n_245) );
INVx2_ASAP7_75t_L g539 ( .A(n_98), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_99), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g216 ( .A(n_100), .B(n_147), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_101), .Y(n_723) );
OAI222xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_719), .B1(n_725), .B2(n_729), .C1(n_730), .C2(n_735), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_112), .B1(n_435), .B2(n_439), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_106), .A2(n_113), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g437 ( .A(n_109), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g734 ( .A(n_109), .Y(n_734) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_112), .A2(n_113), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_SL g113 ( .A(n_114), .B(n_390), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_325), .Y(n_114) );
NAND4xp25_ASAP7_75t_SL g115 ( .A(n_116), .B(n_270), .C(n_294), .D(n_317), .Y(n_115) );
AOI221xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_207), .B1(n_241), .B2(n_254), .C(n_257), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_177), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_119), .A2(n_155), .B1(n_208), .B2(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_119), .B(n_178), .Y(n_328) );
AND2x2_ASAP7_75t_L g347 ( .A(n_119), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_119), .B(n_331), .Y(n_417) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_155), .Y(n_119) );
AND2x2_ASAP7_75t_L g285 ( .A(n_120), .B(n_178), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_120), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g308 ( .A(n_120), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g313 ( .A(n_120), .B(n_156), .Y(n_313) );
INVx2_ASAP7_75t_L g345 ( .A(n_120), .Y(n_345) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_120), .Y(n_389) );
AND2x2_ASAP7_75t_L g406 ( .A(n_120), .B(n_283), .Y(n_406) );
INVx5_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g324 ( .A(n_121), .B(n_283), .Y(n_324) );
AND2x4_ASAP7_75t_L g338 ( .A(n_121), .B(n_155), .Y(n_338) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_121), .Y(n_342) );
AND2x2_ASAP7_75t_L g362 ( .A(n_121), .B(n_277), .Y(n_362) );
AND2x2_ASAP7_75t_L g412 ( .A(n_121), .B(n_179), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_121), .B(n_156), .Y(n_422) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_152), .Y(n_121) );
AOI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_132), .B(n_145), .Y(n_122) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_126), .B(n_130), .Y(n_246) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g143 ( .A(n_127), .Y(n_143) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
INVx1_ASAP7_75t_L g240 ( .A(n_128), .Y(n_240) );
INVx1_ASAP7_75t_L g135 ( .A(n_129), .Y(n_135) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
INVx3_ASAP7_75t_L g168 ( .A(n_129), .Y(n_168) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g236 ( .A(n_129), .Y(n_236) );
BUFx3_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
INVx4_ASAP7_75t_SL g175 ( .A(n_130), .Y(n_175) );
INVx5_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
AND2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx3_ASAP7_75t_L g174 ( .A(n_134), .Y(n_174) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_134), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B(n_142), .Y(n_136) );
INVx2_ASAP7_75t_L g141 ( .A(n_138), .Y(n_141) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx4_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_141), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_141), .A2(n_187), .B(n_214), .C(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_141), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
O2A1O1Ixp5_ASAP7_75t_L g497 ( .A1(n_141), .A2(n_474), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_142), .A2(n_167), .B(n_449), .C(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_143), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_146), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_147), .A2(n_181), .B(n_182), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_147), .A2(n_211), .B(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_147), .A2(n_246), .B(n_446), .C(n_447), .Y(n_445) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_147), .A2(n_482), .B(n_489), .Y(n_481) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_L g160 ( .A(n_148), .B(n_149), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_154), .A2(n_494), .B(n_500), .Y(n_493) );
AND2x2_ASAP7_75t_L g278 ( .A(n_155), .B(n_178), .Y(n_278) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_155), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_155), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g368 ( .A(n_155), .Y(n_368) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g256 ( .A(n_156), .B(n_193), .Y(n_256) );
AND2x2_ASAP7_75t_L g283 ( .A(n_156), .B(n_194), .Y(n_283) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_161), .B(n_176), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_158), .B(n_190), .Y(n_189) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_195), .B(n_205), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_158), .B(n_206), .Y(n_205) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_158), .A2(n_244), .B(n_251), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_158), .B(n_452), .Y(n_451) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_158), .A2(n_468), .B(n_475), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_158), .B(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_159), .A2(n_232), .B(n_233), .Y(n_231) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g253 ( .A(n_160), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B(n_165), .C(n_175), .Y(n_162) );
INVx2_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_164), .A2(n_175), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g459 ( .A1(n_164), .A2(n_175), .B(n_460), .C(n_461), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_164), .A2(n_175), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_164), .A2(n_175), .B(n_506), .C(n_507), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_164), .A2(n_175), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_164), .A2(n_175), .B(n_536), .C(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_167), .B(n_226), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_167), .A2(n_200), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_168), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_171), .B(n_526), .Y(n_525) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g486 ( .A(n_172), .Y(n_486) );
INVx2_ASAP7_75t_L g474 ( .A(n_173), .Y(n_474) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_174), .Y(n_187) );
INVx1_ASAP7_75t_L g510 ( .A(n_174), .Y(n_510) );
INVx1_ASAP7_75t_L g188 ( .A(n_175), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_177), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_191), .Y(n_177) );
OR2x2_ASAP7_75t_L g309 ( .A(n_178), .B(n_192), .Y(n_309) );
AND2x2_ASAP7_75t_L g346 ( .A(n_178), .B(n_256), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_178), .B(n_277), .Y(n_357) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_178), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_178), .B(n_313), .Y(n_430) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g255 ( .A(n_179), .Y(n_255) );
AND2x2_ASAP7_75t_L g264 ( .A(n_179), .B(n_192), .Y(n_264) );
AND2x2_ASAP7_75t_L g380 ( .A(n_179), .B(n_275), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_179), .B(n_313), .Y(n_402) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_189), .Y(n_179) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_192), .Y(n_348) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_193), .Y(n_300) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_201), .C(n_202), .Y(n_197) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_200), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_200), .B(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g527 ( .A(n_203), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_217), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_208), .B(n_290), .Y(n_409) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_209), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g261 ( .A(n_209), .B(n_262), .Y(n_261) );
INVx5_ASAP7_75t_SL g269 ( .A(n_209), .Y(n_269) );
OR2x2_ASAP7_75t_L g292 ( .A(n_209), .B(n_262), .Y(n_292) );
OR2x2_ASAP7_75t_L g302 ( .A(n_209), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g365 ( .A(n_209), .B(n_219), .Y(n_365) );
AND2x2_ASAP7_75t_SL g403 ( .A(n_209), .B(n_218), .Y(n_403) );
NOR4xp25_ASAP7_75t_L g424 ( .A(n_209), .B(n_345), .C(n_425), .D(n_426), .Y(n_424) );
AND2x2_ASAP7_75t_L g434 ( .A(n_209), .B(n_266), .Y(n_434) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_216), .Y(n_209) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g259 ( .A(n_218), .B(n_255), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_218), .B(n_261), .Y(n_428) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_228), .Y(n_218) );
OR2x2_ASAP7_75t_L g268 ( .A(n_219), .B(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_219), .B(n_243), .Y(n_287) );
INVxp67_ASAP7_75t_L g290 ( .A(n_219), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_219), .B(n_262), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_219), .B(n_229), .Y(n_356) );
AND2x2_ASAP7_75t_L g371 ( .A(n_219), .B(n_266), .Y(n_371) );
OR2x2_ASAP7_75t_L g400 ( .A(n_219), .B(n_229), .Y(n_400) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_227), .Y(n_219) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_220), .A2(n_504), .B(n_511), .Y(n_503) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_220), .A2(n_521), .B(n_528), .Y(n_520) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_220), .A2(n_534), .B(n_540), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_228), .B(n_305), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_228), .B(n_269), .Y(n_408) );
OR2x2_ASAP7_75t_L g429 ( .A(n_228), .B(n_306), .Y(n_429) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g242 ( .A(n_229), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g266 ( .A(n_229), .B(n_262), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_229), .B(n_243), .Y(n_281) );
AND2x2_ASAP7_75t_L g351 ( .A(n_229), .B(n_275), .Y(n_351) );
AND2x2_ASAP7_75t_L g385 ( .A(n_229), .B(n_269), .Y(n_385) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_230), .B(n_269), .Y(n_288) );
AND2x2_ASAP7_75t_L g316 ( .A(n_230), .B(n_243), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_237), .B(n_238), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_238), .A2(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_241), .B(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_242), .A2(n_331), .B1(n_367), .B2(n_384), .C(n_386), .Y(n_383) );
INVx5_ASAP7_75t_SL g262 ( .A(n_243), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_247), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_246), .A2(n_469), .B(n_470), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_246), .A2(n_495), .B(n_496), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g457 ( .A(n_253), .Y(n_457) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OAI33xp33_ASAP7_75t_L g282 ( .A1(n_255), .A2(n_283), .A3(n_284), .B1(n_286), .B2(n_289), .B3(n_293), .Y(n_282) );
OR2x2_ASAP7_75t_L g298 ( .A(n_255), .B(n_299), .Y(n_298) );
AOI322xp5_ASAP7_75t_L g407 ( .A1(n_255), .A2(n_324), .A3(n_331), .B1(n_408), .B2(n_409), .C1(n_410), .C2(n_413), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_255), .B(n_283), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_SL g431 ( .A1(n_255), .A2(n_283), .B(n_432), .C(n_434), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_256), .A2(n_271), .B1(n_276), .B2(n_279), .C(n_282), .Y(n_270) );
INVx1_ASAP7_75t_L g363 ( .A(n_256), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_256), .B(n_412), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B1(n_263), .B2(n_265), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g340 ( .A(n_261), .B(n_275), .Y(n_340) );
AND2x2_ASAP7_75t_L g398 ( .A(n_261), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g306 ( .A(n_262), .B(n_269), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_262), .B(n_275), .Y(n_334) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_264), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_264), .B(n_342), .Y(n_396) );
OAI321xp33_ASAP7_75t_L g415 ( .A1(n_264), .A2(n_337), .A3(n_416), .B1(n_417), .B2(n_418), .C(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g382 ( .A(n_265), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_266), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g321 ( .A(n_266), .B(n_269), .Y(n_321) );
AOI321xp33_ASAP7_75t_L g379 ( .A1(n_266), .A2(n_283), .A3(n_380), .B1(n_381), .B2(n_382), .C(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g296 ( .A(n_268), .B(n_281), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_269), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_269), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_269), .B(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g315 ( .A(n_273), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g280 ( .A(n_274), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g388 ( .A(n_275), .Y(n_388) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_278), .B(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g311 ( .A(n_283), .Y(n_311) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_285), .B(n_320), .Y(n_369) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
OR2x2_ASAP7_75t_L g333 ( .A(n_288), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g378 ( .A(n_288), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_289), .A2(n_336), .B1(n_339), .B2(n_341), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g433 ( .A(n_292), .B(n_356), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B1(n_301), .B2(n_307), .C(n_310), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx2_ASAP7_75t_L g331 ( .A(n_300), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_SL g377 ( .A(n_303), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_305), .B(n_355), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_305), .A2(n_373), .B(n_375), .Y(n_372) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g418 ( .A(n_306), .B(n_400), .Y(n_418) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g320 ( .A(n_309), .Y(n_320) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_314), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g364 ( .A(n_316), .B(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_L g426 ( .A(n_316), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_322), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_320), .B(n_338), .Y(n_374) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g395 ( .A(n_324), .Y(n_395) );
NAND5xp2_ASAP7_75t_L g325 ( .A(n_326), .B(n_343), .C(n_352), .D(n_372), .E(n_379), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B(n_332), .C(n_335), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_339), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g381 ( .A(n_341), .Y(n_381) );
OAI21xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_347), .B(n_349), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_344), .A2(n_398), .B1(n_401), .B2(n_403), .C(n_404), .Y(n_397) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
AOI321xp33_ASAP7_75t_L g352 ( .A1(n_345), .A2(n_353), .A3(n_357), .B1(n_358), .B2(n_364), .C(n_366), .Y(n_352) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g423 ( .A(n_357), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_359), .B(n_363), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g375 ( .A(n_360), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
NOR2xp67_ASAP7_75t_SL g387 ( .A(n_361), .B(n_368), .Y(n_387) );
AOI321xp33_ASAP7_75t_SL g419 ( .A1(n_364), .A2(n_420), .A3(n_421), .B1(n_422), .B2(n_423), .C(n_424), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_369), .C(n_370), .Y(n_366) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_377), .B(n_385), .Y(n_414) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .C(n_389), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_415), .C(n_427), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B(n_397), .C(n_407), .Y(n_391) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_395), .B(n_396), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_396), .A2(n_428), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g416 ( .A(n_398), .Y(n_416) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g420 ( .A(n_418), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
CKINVDCx14_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g728 ( .A(n_436), .Y(n_728) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_438), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g727 ( .A(n_439), .Y(n_727) );
OR4x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_609), .C(n_656), .D(n_696), .Y(n_439) );
NAND3xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_555), .C(n_584), .Y(n_440) );
AOI211xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_477), .B(n_512), .C(n_548), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g584 ( .A1(n_442), .A2(n_568), .B(n_585), .C(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_453), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_444), .B(n_547), .Y(n_546) );
INVx3_ASAP7_75t_SL g551 ( .A(n_444), .Y(n_551) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_444), .Y(n_563) );
AND2x4_ASAP7_75t_L g567 ( .A(n_444), .B(n_519), .Y(n_567) );
AND2x2_ASAP7_75t_L g578 ( .A(n_444), .B(n_467), .Y(n_578) );
OR2x2_ASAP7_75t_L g602 ( .A(n_444), .B(n_515), .Y(n_602) );
AND2x2_ASAP7_75t_L g615 ( .A(n_444), .B(n_520), .Y(n_615) );
AND2x2_ASAP7_75t_L g655 ( .A(n_444), .B(n_641), .Y(n_655) );
AND2x2_ASAP7_75t_L g662 ( .A(n_444), .B(n_625), .Y(n_662) );
AND2x2_ASAP7_75t_L g692 ( .A(n_444), .B(n_454), .Y(n_692) );
OR2x6_ASAP7_75t_L g444 ( .A(n_445), .B(n_451), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_453), .B(n_619), .Y(n_631) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_466), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_454), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g569 ( .A(n_454), .B(n_466), .Y(n_569) );
BUFx3_ASAP7_75t_L g577 ( .A(n_454), .Y(n_577) );
OR2x2_ASAP7_75t_L g598 ( .A(n_454), .B(n_480), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_454), .B(n_619), .Y(n_709) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B(n_465), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_456), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g516 ( .A(n_458), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_465), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_466), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g562 ( .A(n_466), .Y(n_562) );
AND2x2_ASAP7_75t_L g625 ( .A(n_466), .B(n_520), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_466), .A2(n_628), .B1(n_630), .B2(n_632), .C(n_633), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_466), .B(n_515), .Y(n_641) );
AND2x2_ASAP7_75t_L g667 ( .A(n_466), .B(n_551), .Y(n_667) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g547 ( .A(n_467), .B(n_520), .Y(n_547) );
BUFx2_ASAP7_75t_L g681 ( .A(n_467), .Y(n_681) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_478), .A2(n_608), .A3(n_622), .B1(n_648), .B2(n_649), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_490), .Y(n_478) );
AND2x2_ASAP7_75t_L g588 ( .A(n_479), .B(n_532), .Y(n_588) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR2x2_ASAP7_75t_L g570 ( .A(n_480), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_480), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g642 ( .A(n_480), .B(n_532), .Y(n_642) );
AND2x2_ASAP7_75t_L g653 ( .A(n_480), .B(n_545), .Y(n_653) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g554 ( .A(n_481), .B(n_533), .Y(n_554) );
AND2x2_ASAP7_75t_L g558 ( .A(n_481), .B(n_533), .Y(n_558) );
AND2x2_ASAP7_75t_L g593 ( .A(n_481), .B(n_544), .Y(n_593) );
AND2x2_ASAP7_75t_L g600 ( .A(n_481), .B(n_502), .Y(n_600) );
OAI211xp5_ASAP7_75t_L g605 ( .A1(n_481), .A2(n_551), .B(n_562), .C(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g659 ( .A(n_481), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_481), .B(n_492), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_490), .B(n_542), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_490), .B(n_558), .Y(n_648) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g553 ( .A(n_491), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
AND2x2_ASAP7_75t_L g545 ( .A(n_492), .B(n_503), .Y(n_545) );
OR2x2_ASAP7_75t_L g560 ( .A(n_492), .B(n_503), .Y(n_560) );
AND2x2_ASAP7_75t_L g583 ( .A(n_492), .B(n_544), .Y(n_583) );
INVx1_ASAP7_75t_L g587 ( .A(n_492), .Y(n_587) );
AND2x2_ASAP7_75t_L g606 ( .A(n_492), .B(n_543), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_492), .A2(n_571), .B1(n_617), .B2(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_492), .B(n_659), .Y(n_683) );
AND2x2_ASAP7_75t_L g698 ( .A(n_492), .B(n_558), .Y(n_698) );
INVx4_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx3_ASAP7_75t_L g530 ( .A(n_493), .Y(n_530) );
AND2x2_ASAP7_75t_L g572 ( .A(n_493), .B(n_503), .Y(n_572) );
AND2x2_ASAP7_75t_L g574 ( .A(n_493), .B(n_532), .Y(n_574) );
AND3x2_ASAP7_75t_L g636 ( .A(n_493), .B(n_600), .C(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g671 ( .A(n_502), .B(n_543), .Y(n_671) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g532 ( .A(n_503), .B(n_533), .Y(n_532) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_503), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_503), .B(n_542), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_503), .B(n_583), .C(n_659), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_529), .B1(n_541), .B2(n_546), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_515), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g623 ( .A(n_515), .Y(n_623) );
OAI31xp33_ASAP7_75t_L g639 ( .A1(n_518), .A2(n_640), .A3(n_641), .B(n_642), .Y(n_639) );
AND2x2_ASAP7_75t_L g664 ( .A(n_518), .B(n_551), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_518), .B(n_577), .Y(n_710) );
AND2x2_ASAP7_75t_L g619 ( .A(n_519), .B(n_551), .Y(n_619) );
AND2x2_ASAP7_75t_L g680 ( .A(n_519), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g550 ( .A(n_520), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g608 ( .A(n_520), .Y(n_608) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g629 ( .A(n_530), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_531), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AOI221x1_ASAP7_75t_SL g596 ( .A1(n_532), .A2(n_597), .B1(n_599), .B2(n_601), .C(n_603), .Y(n_596) );
INVx2_ASAP7_75t_L g544 ( .A(n_533), .Y(n_544) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_533), .Y(n_638) );
INVx1_ASAP7_75t_L g626 ( .A(n_541), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_542), .B(n_559), .Y(n_651) );
INVx1_ASAP7_75t_SL g714 ( .A(n_542), .Y(n_714) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g632 ( .A(n_545), .B(n_558), .Y(n_632) );
INVx1_ASAP7_75t_L g700 ( .A(n_546), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_546), .B(n_629), .Y(n_713) );
INVx2_ASAP7_75t_SL g552 ( .A(n_547), .Y(n_552) );
AND2x2_ASAP7_75t_L g595 ( .A(n_547), .B(n_551), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_547), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_547), .B(n_622), .Y(n_649) );
AOI21xp33_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_552), .B(n_553), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_550), .B(n_622), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_550), .B(n_577), .Y(n_718) );
OR2x2_ASAP7_75t_L g590 ( .A(n_551), .B(n_569), .Y(n_590) );
AND2x2_ASAP7_75t_L g689 ( .A(n_551), .B(n_680), .Y(n_689) );
OAI22xp5_ASAP7_75t_SL g564 ( .A1(n_552), .A2(n_565), .B1(n_570), .B2(n_573), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_552), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g612 ( .A(n_554), .B(n_560), .Y(n_612) );
INVx1_ASAP7_75t_L g676 ( .A(n_554), .Y(n_676) );
AOI311xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_561), .A3(n_563), .B(n_564), .C(n_575), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_559), .A2(n_691), .B1(n_703), .B2(n_706), .C(n_708), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_559), .B(n_714), .Y(n_716) );
INVx2_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g613 ( .A(n_561), .Y(n_613) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_562), .A2(n_604), .B(n_605), .C(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_SL g672 ( .A1(n_566), .A2(n_568), .B(n_673), .C(n_674), .Y(n_672) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_567), .B(n_641), .Y(n_707) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_570), .A2(n_590), .B1(n_591), .B2(n_594), .C(n_596), .Y(n_589) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g592 ( .A(n_572), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g675 ( .A(n_572), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_576), .A2(n_634), .B(n_635), .C(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_577), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_577), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g599 ( .A(n_583), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_587), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g701 ( .A(n_590), .Y(n_701) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_593), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_593), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g705 ( .A(n_593), .Y(n_705) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g646 ( .A(n_595), .B(n_622), .Y(n_646) );
INVx1_ASAP7_75t_SL g640 ( .A(n_602), .Y(n_640) );
INVx1_ASAP7_75t_L g617 ( .A(n_608), .Y(n_617) );
NAND3xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_627), .C(n_643), .Y(n_609) );
AOI322xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .A3(n_614), .B1(n_616), .B2(n_620), .C1(n_624), .C2(n_626), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_611), .A2(n_664), .B(n_665), .C(n_672), .Y(n_663) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_614), .A2(n_635), .B1(n_666), .B2(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_622), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g661 ( .A(n_622), .B(n_662), .Y(n_661) );
AOI32xp33_ASAP7_75t_L g712 ( .A1(n_622), .A2(n_713), .A3(n_714), .B1(n_715), .B2(n_717), .Y(n_712) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g634 ( .A(n_625), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_625), .A2(n_678), .B1(n_682), .B2(n_684), .C(n_687), .Y(n_677) );
AND2x2_ASAP7_75t_L g691 ( .A(n_625), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g694 ( .A(n_629), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g704 ( .A(n_629), .B(n_705), .Y(n_704) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g695 ( .A(n_638), .B(n_659), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B(n_647), .C(n_650), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_660), .B(n_663), .C(n_677), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_671), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g686 ( .A(n_683), .Y(n_686) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_693), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI211xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B(n_702), .C(n_712), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_698), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g729 ( .A(n_719), .Y(n_729) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_742), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_SL g748 ( .A(n_739), .Y(n_748) );
OA21x2_ASAP7_75t_L g746 ( .A1(n_741), .A2(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g769 ( .A(n_741), .Y(n_769) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
BUFx2_ASAP7_75t_L g747 ( .A(n_744), .Y(n_747) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_744), .Y(n_751) );
INVx2_ASAP7_75t_L g765 ( .A(n_744), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g767 ( .A(n_748), .B(n_768), .Y(n_767) );
O2A1O1Ixp33_ASAP7_75t_SL g749 ( .A1(n_750), .A2(n_752), .B(n_761), .C(n_766), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g760 ( .A(n_754), .Y(n_760) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx6p67_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
endmodule