module fake_jpeg_17304_n_349 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_0),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_19),
.B1(n_38),
.B2(n_37),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_36),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_54),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_38),
.B1(n_37),
.B2(n_26),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_22),
.B1(n_34),
.B2(n_27),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_38),
.B1(n_37),
.B2(n_31),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_31),
.B1(n_22),
.B2(n_21),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_30),
.B1(n_55),
.B2(n_34),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_87),
.Y(n_122)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_80),
.B(n_86),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_94),
.B1(n_56),
.B2(n_35),
.Y(n_137)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_105),
.B1(n_56),
.B2(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_85),
.B(n_96),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_70),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_51),
.B1(n_45),
.B2(n_43),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_74),
.B1(n_48),
.B2(n_47),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_40),
.B1(n_44),
.B2(n_28),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_68),
.A2(n_25),
.B1(n_36),
.B2(n_20),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_58),
.B(n_68),
.Y(n_118)
);

CKINVDCx6p67_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_25),
.B1(n_36),
.B2(n_20),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_58),
.B(n_27),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_63),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_18),
.Y(n_135)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_135),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_68),
.C(n_58),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_92),
.B(n_26),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_114),
.B(n_122),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_72),
.A3(n_75),
.B1(n_71),
.B2(n_67),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_122),
.B1(n_137),
.B2(n_123),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_127),
.B1(n_106),
.B2(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_142),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_74),
.B1(n_61),
.B2(n_56),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_49),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_89),
.C(n_23),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_97),
.B1(n_108),
.B2(n_111),
.Y(n_151)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_78),
.B(n_56),
.C(n_23),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_26),
.C(n_23),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_95),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_0),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_145),
.A2(n_158),
.B(n_167),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_147),
.B(n_152),
.Y(n_186)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_155),
.B1(n_160),
.B2(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_102),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_101),
.B1(n_106),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_156),
.B1(n_141),
.B2(n_133),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_137),
.B1(n_131),
.B2(n_122),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_106),
.B1(n_35),
.B2(n_33),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_23),
.C(n_26),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_144),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_169),
.B(n_138),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_118),
.B(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_174),
.B(n_157),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_148),
.B1(n_138),
.B2(n_125),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_181),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_141),
.B(n_134),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_112),
.B1(n_126),
.B2(n_128),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_163),
.B1(n_33),
.B2(n_32),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_190),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_144),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_166),
.C(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_132),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_139),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_196),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_139),
.B(n_112),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_33),
.B(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_128),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_152),
.B(n_120),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_9),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_116),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_217),
.Y(n_240)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_203),
.B(n_190),
.CI(n_177),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_208),
.C(n_215),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_183),
.B1(n_155),
.B2(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_160),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_192),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_164),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_209),
.B(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_151),
.B1(n_161),
.B2(n_165),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_148),
.B1(n_161),
.B2(n_113),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_113),
.B1(n_140),
.B2(n_116),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_140),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_171),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_163),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_194),
.B(n_196),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_219),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_32),
.C(n_29),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.C(n_226),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_11),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_29),
.C(n_20),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_10),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_175),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_212),
.B(n_202),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_170),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_249),
.C(n_250),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_199),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_242),
.B1(n_243),
.B2(n_246),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_248),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_189),
.B1(n_191),
.B2(n_186),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_186),
.B1(n_179),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_192),
.B1(n_188),
.B2(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_180),
.C(n_178),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_178),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_220),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_272),
.C(n_274),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_257),
.B(n_276),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_201),
.B1(n_205),
.B2(n_224),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_262),
.B1(n_269),
.B2(n_238),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_266),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_201),
.B1(n_221),
.B2(n_227),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_218),
.B(n_219),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_264),
.A2(n_231),
.B(n_239),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_252),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_226),
.B1(n_180),
.B2(n_2),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_237),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_180),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_9),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_229),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_244),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_SL g276 ( 
.A(n_233),
.B(n_12),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_250),
.C(n_249),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_285),
.C(n_287),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_290),
.B1(n_264),
.B2(n_260),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_256),
.B1(n_238),
.B2(n_261),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_268),
.B1(n_269),
.B2(n_265),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_251),
.C(n_239),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_237),
.C(n_244),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_273),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_292),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_276),
.B1(n_262),
.B2(n_257),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_245),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_295),
.B(n_18),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_12),
.B(n_17),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_281),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_297),
.A2(n_290),
.B(n_5),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_260),
.B1(n_271),
.B2(n_274),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_303),
.B1(n_304),
.B2(n_300),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_12),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_309),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_0),
.B(n_1),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_286),
.B(n_5),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_29),
.B1(n_18),
.B2(n_13),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_290),
.B1(n_15),
.B2(n_16),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_279),
.B1(n_281),
.B2(n_287),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_298),
.B1(n_308),
.B2(n_307),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_291),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_320),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_278),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_319),
.B1(n_305),
.B2(n_299),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_17),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_303),
.B(n_304),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g325 ( 
.A(n_320),
.B(n_308),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_319),
.B(n_313),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_314),
.A2(n_309),
.B1(n_15),
.B2(n_14),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_315),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_4),
.Y(n_341)
);

AOI21xp33_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_323),
.B(n_15),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_313),
.B(n_316),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_16),
.B(n_17),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_312),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_337),
.B(n_324),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_339),
.A2(n_340),
.B(n_341),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_334),
.A2(n_4),
.B(n_6),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_342),
.Y(n_345)
);

OAI321xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_331),
.A3(n_343),
.B1(n_7),
.B2(n_4),
.C(n_6),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_6),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_347),
.B(n_7),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_7),
.B(n_345),
.Y(n_349)
);


endmodule