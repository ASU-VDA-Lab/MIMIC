module fake_jpeg_28189_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_28),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_56),
.B(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_62),
.B1(n_30),
.B2(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_21),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_60),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_18),
.B1(n_24),
.B2(n_34),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_66),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_70),
.B1(n_61),
.B2(n_41),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_19),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_36),
.B1(n_43),
.B2(n_40),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_73),
.Y(n_93)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_23),
.B1(n_30),
.B2(n_26),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_44),
.B(n_41),
.C(n_35),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_80),
.B1(n_28),
.B2(n_1),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_44),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_32),
.C(n_33),
.Y(n_94)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_44),
.B1(n_35),
.B2(n_41),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_55),
.A3(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_98),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_33),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_32),
.B1(n_31),
.B2(n_28),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_16),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_6),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_67),
.B1(n_65),
.B2(n_83),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_76),
.B(n_65),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_123),
.B(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_119),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_126),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_89),
.B(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_131),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_133),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_75),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_139),
.Y(n_176)
);

BUFx4f_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_103),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_160),
.B(n_154),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_124),
.B1(n_131),
.B2(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_91),
.C(n_98),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_156),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_90),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_159),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_107),
.C(n_101),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_111),
.C(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_127),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_170),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_175),
.B1(n_142),
.B2(n_157),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_116),
.C(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_117),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_159),
.B1(n_143),
.B2(n_120),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_82),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_191),
.Y(n_196)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_156),
.B1(n_145),
.B2(n_140),
.C(n_146),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_146),
.B1(n_153),
.B2(n_73),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_185),
.B1(n_167),
.B2(n_178),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_141),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_141),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_162),
.B(n_176),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_72),
.B1(n_66),
.B2(n_88),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_63),
.B1(n_88),
.B2(n_15),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_187),
.B1(n_162),
.B2(n_172),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_166),
.B1(n_177),
.B2(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_201),
.C(n_202),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_164),
.B(n_171),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_176),
.B1(n_169),
.B2(n_63),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_188),
.C(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_190),
.C(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_186),
.C(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_201),
.Y(n_212)
);

OAI221xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_216),
.B1(n_209),
.B2(n_211),
.C(n_9),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_221),
.B(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.C(n_6),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_211),
.C(n_15),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_14),
.B(n_8),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_11),
.C(n_9),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);


endmodule