module real_aes_7133_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g515 ( .A(n_1), .Y(n_515) );
INVx1_ASAP7_75t_L g148 ( .A(n_2), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_3), .A2(n_38), .B1(n_173), .B2(n_461), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g180 ( .A1(n_4), .A2(n_164), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_5), .B(n_162), .Y(n_527) );
AND2x6_ASAP7_75t_L g141 ( .A(n_6), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_39), .Y(n_113) );
INVx1_ASAP7_75t_L g186 ( .A(n_9), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g133 ( .A(n_11), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_12), .B(n_154), .Y(n_470) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
INVx1_ASAP7_75t_L g509 ( .A(n_14), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_15), .B(n_129), .Y(n_498) );
AO32x2_ASAP7_75t_L g482 ( .A1(n_16), .A2(n_128), .A3(n_162), .B1(n_463), .B2(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_17), .B(n_173), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_18), .B(n_169), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_19), .B(n_129), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_20), .A2(n_49), .B1(n_173), .B2(n_461), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_21), .B(n_164), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_22), .A2(n_96), .B1(n_715), .B2(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_22), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_23), .A2(n_74), .B1(n_154), .B2(n_173), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_24), .B(n_173), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_25), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_26), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_28), .B(n_159), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_29), .B(n_152), .Y(n_151) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_30), .A2(n_101), .B1(n_114), .B2(n_722), .C1(n_728), .C2(n_737), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_30), .A2(n_87), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_30), .Y(n_731) );
INVx1_ASAP7_75t_L g201 ( .A(n_31), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_32), .B(n_159), .Y(n_454) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_33), .A2(n_116), .B1(n_713), .B2(n_714), .C1(n_717), .C2(n_719), .Y(n_115) );
INVx2_ASAP7_75t_L g139 ( .A(n_34), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_35), .B(n_173), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_36), .B(n_159), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_141), .B(n_144), .C(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g199 ( .A(n_40), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_41), .B(n_152), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_42), .B(n_173), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_43), .A2(n_84), .B1(n_221), .B2(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_44), .B(n_173), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_45), .B(n_173), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_46), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_47), .B(n_514), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_48), .B(n_164), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_50), .A2(n_59), .B1(n_154), .B2(n_173), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_51), .A2(n_144), .B1(n_154), .B2(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_52), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_53), .B(n_173), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g135 ( .A(n_54), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_55), .B(n_173), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_56), .A2(n_172), .B(n_184), .C(n_185), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_57), .Y(n_234) );
INVx1_ASAP7_75t_L g182 ( .A(n_58), .Y(n_182) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_61), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_62), .B(n_173), .Y(n_516) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_64), .Y(n_106) );
AO32x2_ASAP7_75t_L g458 ( .A1(n_65), .A2(n_162), .A3(n_237), .B1(n_459), .B2(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g534 ( .A(n_66), .Y(n_534) );
INVx1_ASAP7_75t_L g449 ( .A(n_67), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_SL g168 ( .A1(n_68), .A2(n_169), .B(n_170), .C(n_172), .Y(n_168) );
INVxp67_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_70), .B(n_154), .Y(n_450) );
INVx1_ASAP7_75t_L g105 ( .A(n_71), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_72), .Y(n_204) );
INVx1_ASAP7_75t_L g227 ( .A(n_73), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_75), .A2(n_141), .B(n_144), .C(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_76), .B(n_461), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_77), .B(n_154), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_78), .B(n_149), .Y(n_217) );
INVx2_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_80), .B(n_169), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_81), .B(n_154), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_82), .A2(n_141), .B(n_144), .C(n_147), .Y(n_143) );
OR2x2_ASAP7_75t_L g109 ( .A(n_83), .B(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g119 ( .A(n_83), .B(n_111), .Y(n_119) );
INVx2_ASAP7_75t_L g436 ( .A(n_83), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_85), .A2(n_99), .B1(n_154), .B2(n_155), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_86), .B(n_159), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_87), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_88), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_89), .A2(n_141), .B(n_144), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_90), .Y(n_247) );
INVx1_ASAP7_75t_L g167 ( .A(n_91), .Y(n_167) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_92), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_93), .B(n_149), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_94), .B(n_154), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_95), .B(n_162), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_96), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_98), .A2(n_164), .B(n_165), .Y(n_163) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_SL g727 ( .A(n_104), .Y(n_727) );
INVx1_ASAP7_75t_L g726 ( .A(n_106), .Y(n_726) );
OA21x2_ASAP7_75t_L g738 ( .A1(n_106), .A2(n_727), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_109), .Y(n_734) );
INVx2_ASAP7_75t_L g736 ( .A(n_109), .Y(n_736) );
BUFx2_ASAP7_75t_L g739 ( .A(n_109), .Y(n_739) );
NOR2x2_ASAP7_75t_L g721 ( .A(n_110), .B(n_436), .Y(n_721) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g435 ( .A(n_111), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_433), .B2(n_437), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g718 ( .A(n_118), .Y(n_718) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_121), .A2(n_433), .B1(n_438), .B2(n_718), .Y(n_717) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_121), .B(n_730), .Y(n_729) );
NAND2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_349), .Y(n_121) );
NOR5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_272), .C(n_304), .D(n_319), .E(n_336), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_188), .B(n_209), .C(n_260), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_125), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_125), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_126), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_126), .B(n_206), .Y(n_273) );
AND2x2_ASAP7_75t_L g314 ( .A(n_126), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_126), .B(n_283), .Y(n_318) );
OR2x2_ASAP7_75t_L g355 ( .A(n_126), .B(n_194), .Y(n_355) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g193 ( .A(n_127), .B(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g263 ( .A(n_127), .Y(n_263) );
OR2x2_ASAP7_75t_L g426 ( .A(n_127), .B(n_266), .Y(n_426) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B(n_156), .Y(n_127) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_128), .A2(n_195), .B(n_203), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_128), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g222 ( .A(n_128), .Y(n_222) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_130), .B(n_131), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_143), .Y(n_134) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_136), .A2(n_174), .B1(n_196), .B2(n_202), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_136), .A2(n_227), .B(n_228), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
AND2x4_ASAP7_75t_L g164 ( .A(n_137), .B(n_141), .Y(n_164) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g514 ( .A(n_138), .Y(n_514) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_140), .Y(n_198) );
INVx4_ASAP7_75t_SL g174 ( .A(n_141), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_141), .A2(n_448), .B(n_451), .Y(n_447) );
BUFx3_ASAP7_75t_L g463 ( .A(n_141), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_141), .A2(n_468), .B(n_472), .Y(n_467) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_141), .A2(n_508), .B(n_512), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_141), .A2(n_521), .B(n_524), .Y(n_520) );
INVx5_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
BUFx3_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
INVx1_ASAP7_75t_L g461 ( .A(n_145), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_151), .C(n_153), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_SL g448 ( .A1(n_149), .A2(n_172), .B(n_449), .C(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g485 ( .A(n_149), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_149), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_149), .A2(n_531), .B(n_532), .Y(n_530) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_150), .B(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_150), .B(n_186), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_150), .A2(n_152), .B1(n_460), .B2(n_462), .Y(n_459) );
INVx2_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx4_ASAP7_75t_L g243 ( .A(n_152), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_152), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_152), .A2(n_485), .B1(n_501), .B2(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_153), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_158), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_158), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g237 ( .A(n_159), .Y(n_237) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_159), .A2(n_447), .B(n_454), .Y(n_446) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_159), .A2(n_467), .B(n_475), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_160), .A2(n_329), .B1(n_330), .B2(n_333), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_160), .B(n_263), .Y(n_412) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_178), .Y(n_160) );
AND2x2_ASAP7_75t_L g208 ( .A(n_161), .B(n_194), .Y(n_208) );
AND2x2_ASAP7_75t_L g265 ( .A(n_161), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g270 ( .A(n_161), .Y(n_270) );
INVx3_ASAP7_75t_L g283 ( .A(n_161), .Y(n_283) );
OR2x2_ASAP7_75t_L g303 ( .A(n_161), .B(n_266), .Y(n_303) );
AND2x2_ASAP7_75t_L g322 ( .A(n_161), .B(n_179), .Y(n_322) );
BUFx2_ASAP7_75t_L g354 ( .A(n_161), .Y(n_354) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_175), .Y(n_161) );
INVx4_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_162), .A2(n_520), .B(n_527), .Y(n_519) );
BUFx2_ASAP7_75t_L g251 ( .A(n_164), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_174), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_166), .A2(n_174), .B(n_182), .C(n_183), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_166), .A2(n_174), .B(n_253), .C(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g471 ( .A(n_169), .Y(n_471) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_176), .A2(n_180), .B(n_187), .Y(n_179) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_177), .B(n_224), .Y(n_223) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_177), .B(n_463), .C(n_500), .Y(n_499) );
AO21x1_ASAP7_75t_L g589 ( .A1(n_177), .A2(n_500), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g269 ( .A(n_178), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
BUFx2_ASAP7_75t_L g192 ( .A(n_179), .Y(n_192) );
INVx2_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
OR2x2_ASAP7_75t_L g285 ( .A(n_179), .B(n_266), .Y(n_285) );
AND2x2_ASAP7_75t_L g315 ( .A(n_179), .B(n_194), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_179), .B(n_263), .Y(n_332) );
AND2x2_ASAP7_75t_L g372 ( .A(n_179), .B(n_283), .Y(n_372) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_179), .B(n_208), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_184), .A2(n_473), .B(n_474), .Y(n_472) );
O2A1O1Ixp5_ASAP7_75t_L g533 ( .A1(n_184), .A2(n_513), .B(n_534), .C(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp33_ASAP7_75t_SL g189 ( .A(n_190), .B(n_205), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_191), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_192), .A2(n_208), .B(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_192), .B(n_194), .Y(n_402) );
AND2x2_ASAP7_75t_L g338 ( .A(n_193), .B(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g266 ( .A(n_194), .Y(n_266) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_194), .Y(n_364) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g200 ( .A(n_198), .Y(n_200) );
INVx4_ASAP7_75t_L g255 ( .A(n_198), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_205), .B(n_263), .Y(n_431) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_206), .A2(n_374), .B1(n_375), .B2(n_380), .Y(n_373) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AND2x2_ASAP7_75t_L g264 ( .A(n_207), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g302 ( .A(n_207), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g339 ( .A(n_207), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_208), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g393 ( .A(n_208), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_235), .Y(n_210) );
INVx4_ASAP7_75t_L g279 ( .A(n_211), .Y(n_279) );
AND2x2_ASAP7_75t_L g357 ( .A(n_211), .B(n_324), .Y(n_357) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
INVx3_ASAP7_75t_L g276 ( .A(n_212), .Y(n_276) );
AND2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g294 ( .A(n_212), .Y(n_294) );
INVx2_ASAP7_75t_L g308 ( .A(n_212), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_212), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g365 ( .A(n_212), .B(n_360), .Y(n_365) );
AND2x2_ASAP7_75t_L g430 ( .A(n_212), .B(n_400), .Y(n_430) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_219), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
INVx1_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_222), .A2(n_507), .B(n_517), .Y(n_506) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_222), .A2(n_529), .B(n_536), .Y(n_528) );
AND2x2_ASAP7_75t_L g271 ( .A(n_225), .B(n_249), .Y(n_271) );
INVx2_ASAP7_75t_L g291 ( .A(n_225), .Y(n_291) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_233), .Y(n_225) );
INVx1_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
AND2x2_ASAP7_75t_L g342 ( .A(n_235), .B(n_290), .Y(n_342) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
INVx2_ASAP7_75t_L g281 ( .A(n_236), .Y(n_281) );
INVx1_ASAP7_75t_L g289 ( .A(n_236), .Y(n_289) );
AND2x2_ASAP7_75t_L g307 ( .A(n_236), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_236), .B(n_291), .Y(n_345) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
AND2x2_ASAP7_75t_L g324 ( .A(n_248), .B(n_281), .Y(n_324) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
AND2x2_ASAP7_75t_L g360 ( .A(n_249), .B(n_291), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_255), .A2(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g511 ( .A(n_255), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_267), .B(n_271), .Y(n_260) );
INVx1_ASAP7_75t_SL g305 ( .A(n_261), .Y(n_305) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_262), .B(n_269), .Y(n_362) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g311 ( .A(n_263), .B(n_266), .Y(n_311) );
AND2x2_ASAP7_75t_L g340 ( .A(n_263), .B(n_284), .Y(n_340) );
OR2x2_ASAP7_75t_L g343 ( .A(n_263), .B(n_303), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g407 ( .A1(n_264), .A2(n_356), .B1(n_408), .B2(n_409), .C1(n_411), .C2(n_413), .Y(n_407) );
BUFx2_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g310 ( .A(n_269), .B(n_311), .Y(n_310) );
INVx3_ASAP7_75t_SL g327 ( .A(n_269), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_269), .B(n_321), .Y(n_381) );
AND2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_276), .Y(n_316) );
INVx1_ASAP7_75t_L g335 ( .A(n_271), .Y(n_335) );
OAI221xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_274), .B1(n_278), .B2(n_282), .C(n_286), .Y(n_272) );
OR2x2_ASAP7_75t_L g344 ( .A(n_274), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g329 ( .A(n_276), .B(n_299), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_276), .B(n_289), .Y(n_369) );
AND2x2_ASAP7_75t_L g374 ( .A(n_276), .B(n_324), .Y(n_374) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_276), .Y(n_384) );
NAND2x1_ASAP7_75t_SL g395 ( .A(n_276), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g280 ( .A(n_277), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_277), .B(n_295), .Y(n_326) );
INVx1_ASAP7_75t_L g392 ( .A(n_277), .Y(n_392) );
INVx1_ASAP7_75t_L g367 ( .A(n_278), .Y(n_367) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g379 ( .A(n_279), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_279), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g396 ( .A(n_280), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_280), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g299 ( .A(n_281), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_281), .B(n_291), .Y(n_312) );
INVx1_ASAP7_75t_L g378 ( .A(n_281), .Y(n_378) );
INVx1_ASAP7_75t_L g399 ( .A(n_282), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI21xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_292), .B(n_301), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x2_ASAP7_75t_L g432 ( .A(n_288), .B(n_365), .Y(n_432) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g400 ( .A(n_289), .B(n_360), .Y(n_400) );
AOI32xp33_ASAP7_75t_L g313 ( .A1(n_290), .A2(n_296), .A3(n_314), .B1(n_316), .B2(n_317), .Y(n_313) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_290), .A2(n_322), .A3(n_405), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g295 ( .A(n_291), .Y(n_295) );
INVx1_ASAP7_75t_L g405 ( .A(n_291), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_297), .B2(n_298), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_293), .B(n_299), .Y(n_348) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_294), .B(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g297 ( .A(n_295), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_295), .B(n_324), .Y(n_414) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_303), .B(n_398), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_306), .B1(n_309), .B2(n_312), .C(n_313), .Y(n_304) );
OR2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g359 ( .A(n_307), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g363 ( .A(n_317), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B1(n_325), .B2(n_327), .C(n_328), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_322), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_322), .Y(n_427) );
INVx1_ASAP7_75t_L g421 ( .A(n_324), .Y(n_421) );
INVx1_ASAP7_75t_SL g356 ( .A(n_325), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_327), .B(n_355), .Y(n_417) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g398 ( .A(n_332), .Y(n_398) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_341), .B1(n_343), .B2(n_344), .C(n_346), .Y(n_336) );
NOR2xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_340), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_338), .A2(n_356), .B1(n_402), .B2(n_403), .Y(n_401) );
CKINVDCx14_ASAP7_75t_R g341 ( .A(n_342), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g420 ( .A1(n_343), .A2(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR3xp33_ASAP7_75t_SL g349 ( .A(n_350), .B(n_382), .C(n_406), .Y(n_349) );
NAND4xp25_ASAP7_75t_L g350 ( .A(n_351), .B(n_358), .C(n_366), .D(n_373), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
INVx3_ASAP7_75t_SL g423 ( .A(n_355), .Y(n_423) );
OR2x2_ASAP7_75t_L g428 ( .A(n_355), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_363), .B2(n_365), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_360), .B(n_378), .Y(n_419) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI21xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_368), .B(n_370), .Y(n_366) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_388), .C(n_401), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g416 ( .A(n_387), .Y(n_416) );
AOI222xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_393), .B1(n_394), .B2(n_397), .C1(n_399), .C2(n_400), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND4xp25_ASAP7_75t_SL g425 ( .A(n_398), .B(n_426), .C(n_427), .D(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_415), .C(n_424), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_424) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_634), .Y(n_438) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_583), .C(n_625), .Y(n_439) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_492), .B(n_537), .C(n_559), .Y(n_440) );
OAI211xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_455), .B(n_476), .C(n_487), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_443), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g646 ( .A(n_443), .B(n_563), .Y(n_646) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g548 ( .A(n_444), .B(n_479), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_444), .B(n_466), .Y(n_665) );
INVx1_ASAP7_75t_L g683 ( .A(n_444), .Y(n_683) );
AND2x2_ASAP7_75t_L g692 ( .A(n_444), .B(n_580), .Y(n_692) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g575 ( .A(n_445), .B(n_466), .Y(n_575) );
AND2x2_ASAP7_75t_L g633 ( .A(n_445), .B(n_580), .Y(n_633) );
INVx1_ASAP7_75t_L g677 ( .A(n_445), .Y(n_677) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g554 ( .A(n_446), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g562 ( .A(n_446), .Y(n_562) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_446), .Y(n_602) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_464), .Y(n_456) );
AND2x2_ASAP7_75t_L g541 ( .A(n_457), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g574 ( .A(n_457), .Y(n_574) );
OR2x2_ASAP7_75t_L g700 ( .A(n_457), .B(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_457), .B(n_466), .Y(n_704) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g479 ( .A(n_458), .Y(n_479) );
INVx1_ASAP7_75t_L g490 ( .A(n_458), .Y(n_490) );
AND2x2_ASAP7_75t_L g563 ( .A(n_458), .B(n_481), .Y(n_563) );
AND2x2_ASAP7_75t_L g603 ( .A(n_458), .B(n_482), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_463), .A2(n_530), .B(n_533), .Y(n_529) );
INVxp67_ASAP7_75t_L g645 ( .A(n_464), .Y(n_645) );
AND2x4_ASAP7_75t_L g670 ( .A(n_464), .B(n_563), .Y(n_670) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_465), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g480 ( .A(n_466), .B(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g549 ( .A(n_466), .B(n_482), .Y(n_549) );
INVx1_ASAP7_75t_L g555 ( .A(n_466), .Y(n_555) );
INVx2_ASAP7_75t_L g581 ( .A(n_466), .Y(n_581) );
AND2x2_ASAP7_75t_L g597 ( .A(n_466), .B(n_598), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_477), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g552 ( .A(n_479), .Y(n_552) );
AND2x2_ASAP7_75t_L g660 ( .A(n_479), .B(n_481), .Y(n_660) );
AND2x2_ASAP7_75t_L g577 ( .A(n_480), .B(n_562), .Y(n_577) );
AND2x2_ASAP7_75t_L g676 ( .A(n_480), .B(n_677), .Y(n_676) );
NOR2xp67_ASAP7_75t_L g598 ( .A(n_481), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g701 ( .A(n_481), .B(n_562), .Y(n_701) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx2_ASAP7_75t_L g491 ( .A(n_482), .Y(n_491) );
AND2x2_ASAP7_75t_L g580 ( .A(n_482), .B(n_581), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_485), .A2(n_513), .B(n_515), .C(n_516), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_485), .A2(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
AND2x2_ASAP7_75t_L g626 ( .A(n_489), .B(n_561), .Y(n_626) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_490), .B(n_562), .Y(n_611) );
INVx2_ASAP7_75t_L g610 ( .A(n_491), .Y(n_610) );
OAI222xp33_ASAP7_75t_L g614 ( .A1(n_491), .A2(n_554), .B1(n_615), .B2(n_617), .C1(n_618), .C2(n_621), .Y(n_614) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g539 ( .A(n_496), .Y(n_539) );
OR2x2_ASAP7_75t_L g650 ( .A(n_496), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g572 ( .A(n_497), .Y(n_572) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_497), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g629 ( .A(n_497), .B(n_543), .Y(n_629) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g590 ( .A(n_498), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_503), .A2(n_593), .B1(n_632), .B2(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_518), .Y(n_503) );
INVx3_ASAP7_75t_L g565 ( .A(n_504), .Y(n_565) );
OR2x2_ASAP7_75t_L g698 ( .A(n_504), .B(n_574), .Y(n_698) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g587 ( .A(n_505), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g595 ( .A(n_505), .B(n_543), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_505), .B(n_519), .Y(n_651) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g542 ( .A(n_506), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g546 ( .A(n_506), .B(n_519), .Y(n_546) );
AND2x2_ASAP7_75t_L g622 ( .A(n_506), .B(n_569), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_506), .B(n_528), .Y(n_662) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_518), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_518), .B(n_539), .Y(n_578) );
AND2x2_ASAP7_75t_L g582 ( .A(n_518), .B(n_572), .Y(n_582) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
INVx3_ASAP7_75t_L g543 ( .A(n_519), .Y(n_543) );
AND2x2_ASAP7_75t_L g568 ( .A(n_519), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g703 ( .A(n_519), .B(n_686), .Y(n_703) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
INVx2_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
AND2x2_ASAP7_75t_L g613 ( .A(n_528), .B(n_589), .Y(n_613) );
INVx1_ASAP7_75t_L g656 ( .A(n_528), .Y(n_656) );
OR2x2_ASAP7_75t_L g687 ( .A(n_528), .B(n_589), .Y(n_687) );
AND2x2_ASAP7_75t_L g707 ( .A(n_528), .B(n_543), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .B(n_544), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g545 ( .A(n_539), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_539), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g664 ( .A(n_541), .Y(n_664) );
INVx2_ASAP7_75t_SL g558 ( .A(n_542), .Y(n_558) );
AND2x2_ASAP7_75t_L g678 ( .A(n_542), .B(n_572), .Y(n_678) );
INVx2_ASAP7_75t_L g624 ( .A(n_543), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_543), .B(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B1(n_550), .B2(n_556), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_546), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g712 ( .A(n_546), .Y(n_712) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g637 ( .A(n_548), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_548), .B(n_580), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_549), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g653 ( .A(n_549), .B(n_602), .Y(n_653) );
INVx2_ASAP7_75t_L g709 ( .A(n_549), .Y(n_709) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
AND2x2_ASAP7_75t_L g579 ( .A(n_552), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_552), .B(n_597), .Y(n_630) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_554), .B(n_574), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g691 ( .A(n_557), .Y(n_691) );
O2A1O1Ixp33_ASAP7_75t_SL g641 ( .A1(n_558), .A2(n_642), .B(n_644), .C(n_647), .Y(n_641) );
OR2x2_ASAP7_75t_L g668 ( .A(n_558), .B(n_572), .Y(n_668) );
OAI221xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_564), .B1(n_566), .B2(n_573), .C(n_576), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_561), .B(n_610), .Y(n_617) );
AND2x2_ASAP7_75t_L g659 ( .A(n_561), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g695 ( .A(n_561), .Y(n_695) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
INVx1_ASAP7_75t_L g599 ( .A(n_562), .Y(n_599) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_565), .B(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g673 ( .A(n_565), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_565), .B(n_613), .Y(n_689) );
INVx2_ASAP7_75t_L g675 ( .A(n_566), .Y(n_675) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_570), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g616 ( .A(n_568), .B(n_587), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_568), .A2(n_584), .B(n_626), .C(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g594 ( .A(n_569), .B(n_589), .Y(n_594) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_573), .B(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g642 ( .A(n_574), .B(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_582), .Y(n_576) );
INVx1_ASAP7_75t_L g696 ( .A(n_578), .Y(n_696) );
INVx1_ASAP7_75t_L g643 ( .A(n_580), .Y(n_643) );
INVx1_ASAP7_75t_L g694 ( .A(n_582), .Y(n_694) );
AOI211xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_587), .B(n_591), .C(n_614), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g606 ( .A(n_586), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g657 ( .A(n_587), .Y(n_657) );
AND2x2_ASAP7_75t_L g706 ( .A(n_587), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B(n_604), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g620 ( .A(n_594), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_594), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g612 ( .A(n_595), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g688 ( .A(n_595), .Y(n_688) );
OAI32xp33_ASAP7_75t_L g699 ( .A1(n_595), .A2(n_647), .A3(n_654), .B1(n_695), .B2(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_597), .B(n_600), .Y(n_596) );
INVx1_ASAP7_75t_SL g667 ( .A(n_597), .Y(n_667) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g607 ( .A(n_603), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B(n_612), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_606), .A2(n_654), .B1(n_680), .B2(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_610), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g647 ( .A(n_613), .Y(n_647) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g640 ( .A(n_624), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_633), .A2(n_675), .B1(n_676), .B2(n_678), .C(n_679), .Y(n_674) );
NAND5xp2_ASAP7_75t_L g634 ( .A(n_635), .B(n_658), .C(n_674), .D(n_684), .E(n_702), .Y(n_634) );
AOI211xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_638), .B(n_641), .C(n_648), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g705 ( .A(n_642), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_654), .Y(n_648) );
INVx1_ASAP7_75t_SL g681 ( .A(n_651), .Y(n_681) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI322xp33_ASAP7_75t_L g663 ( .A1(n_654), .A2(n_664), .A3(n_665), .B1(n_666), .B2(n_667), .C1(n_668), .C2(n_669), .Y(n_663) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g666 ( .A(n_656), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_656), .B(n_681), .Y(n_680) );
AOI211xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_661), .B(n_663), .C(n_671), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_667), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g710 ( .A(n_677), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_692), .B1(n_693), .B2(n_697), .C(n_699), .Y(n_684) );
OAI211xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_688), .B(n_689), .C(n_690), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g711 ( .A(n_687), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .C(n_708), .Y(n_702) );
AOI21xp33_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_710), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
CKINVDCx6p67_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_733), .B(n_735), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
endmodule