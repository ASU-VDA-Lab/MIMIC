module fake_aes_8248_n_909 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_909);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_909;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_98), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_26), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_36), .B(n_7), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_88), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_100), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_51), .Y(n_118) );
INVx2_ASAP7_75t_SL g119 ( .A(n_67), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_29), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_12), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_34), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_4), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_106), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_109), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_93), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_94), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_15), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_30), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_1), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_2), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_60), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_16), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_75), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_35), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_68), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_89), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_96), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_6), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_78), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_33), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_104), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_15), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_54), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_55), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_1), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_46), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_38), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_73), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_137), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_111), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_129), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_119), .B(n_0), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_132), .B(n_0), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_137), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_112), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_123), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g168 ( .A(n_113), .B(n_18), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
INVx5_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_121), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_122), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_142), .B(n_3), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_121), .Y(n_177) );
INVx1_ASAP7_75t_SL g178 ( .A(n_155), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_175), .B(n_155), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_155), .B(n_134), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_175), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_155), .B(n_124), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_166), .B(n_131), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_174), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_177), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_169), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_177), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
NAND2xp33_ASAP7_75t_SL g196 ( .A(n_175), .B(n_122), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_156), .B(n_114), .Y(n_197) );
NAND2xp33_ASAP7_75t_SL g198 ( .A(n_175), .B(n_128), .Y(n_198) );
INVx5_ASAP7_75t_L g199 ( .A(n_164), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_166), .B(n_117), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_167), .B(n_143), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_169), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_171), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_167), .B(n_120), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_177), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_173), .B(n_147), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_174), .A2(n_140), .B1(n_128), .B2(n_149), .Y(n_208) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_173), .A2(n_153), .B(n_136), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_139), .B(n_151), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_177), .Y(n_211) );
BUFx6f_ASAP7_75t_SL g212 ( .A(n_169), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_177), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_170), .B(n_125), .Y(n_215) );
INVx8_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_160), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_170), .B(n_126), .Y(n_218) );
NOR2x1p5_ASAP7_75t_L g219 ( .A(n_159), .B(n_150), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_176), .B(n_138), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_170), .B(n_130), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_177), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_170), .B(n_145), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_191), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_183), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_213), .B(n_163), .Y(n_228) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_209), .A2(n_148), .B(n_115), .Y(n_229) );
INVx8_ASAP7_75t_L g230 ( .A(n_179), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_186), .B(n_163), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_208), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_179), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_178), .B(n_168), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g235 ( .A(n_212), .B(n_140), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_180), .B(n_171), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_183), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_192), .B(n_193), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_200), .B(n_165), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_179), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_201), .B(n_165), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_187), .B(n_146), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g245 ( .A1(n_179), .A2(n_141), .B1(n_144), .B2(n_149), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_185), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_185), .A2(n_171), .B(n_172), .Y(n_247) );
INVx8_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
NOR2xp67_ASAP7_75t_L g249 ( .A(n_195), .B(n_171), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_219), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_201), .B(n_152), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_191), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_204), .B(n_121), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_207), .Y(n_254) );
NOR2xp67_ASAP7_75t_SL g255 ( .A(n_212), .B(n_121), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_185), .A2(n_172), .B(n_162), .C(n_160), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_172), .B1(n_144), .B2(n_141), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_207), .B(n_172), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_197), .B(n_164), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_210), .B(n_164), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_225), .B(n_164), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_220), .B(n_160), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_203), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_189), .B(n_5), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_202), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_196), .A2(n_162), .B1(n_160), .B2(n_7), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_215), .B(n_160), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_209), .B(n_202), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_218), .B(n_160), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_203), .Y(n_271) );
NOR3xp33_ASAP7_75t_L g272 ( .A(n_196), .B(n_5), .C(n_6), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_222), .B(n_162), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_216), .B(n_162), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_198), .B(n_162), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_198), .B(n_162), .Y(n_276) );
INVxp33_ASAP7_75t_L g277 ( .A(n_189), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_205), .B(n_19), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_205), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_190), .A2(n_8), .B(n_9), .C(n_10), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_190), .B(n_20), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_212), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_182), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_221), .B(n_11), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_221), .B(n_11), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_181), .B(n_13), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_224), .B(n_13), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_224), .B(n_14), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_268), .A2(n_194), .B(n_214), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_230), .A2(n_194), .B1(n_214), .B2(n_211), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_254), .A2(n_206), .B(n_211), .C(n_184), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_230), .A2(n_206), .B1(n_188), .B2(n_184), .Y(n_292) );
OA22x2_ASAP7_75t_L g293 ( .A1(n_232), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_228), .B(n_17), .Y(n_294) );
NAND2x1p5_ASAP7_75t_L g295 ( .A(n_233), .B(n_199), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_240), .B(n_199), .Y(n_297) );
NOR2xp33_ASAP7_75t_R g298 ( .A(n_235), .B(n_21), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_243), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_231), .A2(n_188), .B(n_182), .C(n_199), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_241), .B(n_199), .Y(n_301) );
INVxp33_ASAP7_75t_SL g302 ( .A(n_257), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_240), .B(n_199), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_228), .B(n_181), .Y(n_304) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_181), .B(n_217), .Y(n_305) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_247), .A2(n_181), .B(n_217), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_227), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_230), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_241), .B(n_181), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g311 ( .A1(n_272), .A2(n_22), .B(n_23), .C(n_24), .Y(n_311) );
AOI21x1_ASAP7_75t_L g312 ( .A1(n_247), .A2(n_217), .B(n_27), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_257), .A2(n_217), .B1(n_28), .B2(n_31), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_251), .B(n_25), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_246), .A2(n_217), .B(n_37), .C(n_39), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_273), .A2(n_32), .B(n_41), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_241), .B(n_42), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_250), .B(n_43), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g319 ( .A1(n_246), .A2(n_45), .B1(n_47), .B2(n_48), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_258), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_261), .A2(n_49), .B(n_50), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_237), .Y(n_323) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_245), .Y(n_324) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_242), .B(n_52), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_271), .A2(n_53), .B(n_57), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_260), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_245), .A2(n_58), .B1(n_59), .B2(n_61), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_239), .A2(n_62), .B(n_63), .C(n_64), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_279), .A2(n_65), .B(n_66), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_269), .A2(n_69), .B(n_70), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_239), .B(n_110), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_248), .B(n_71), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_253), .A2(n_72), .B(n_74), .C(n_76), .Y(n_334) );
AO21x1_ASAP7_75t_L g335 ( .A1(n_286), .A2(n_77), .B(n_80), .Y(n_335) );
BUFx8_ASAP7_75t_L g336 ( .A(n_265), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g337 ( .A1(n_248), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_269), .A2(n_84), .B(n_86), .Y(n_338) );
AOI21x1_ASAP7_75t_L g339 ( .A1(n_236), .A2(n_87), .B(n_90), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_275), .A2(n_91), .B(n_92), .Y(n_340) );
BUFx12f_ASAP7_75t_L g341 ( .A(n_307), .Y(n_341) );
OAI21x1_ASAP7_75t_L g342 ( .A1(n_339), .A2(n_276), .B(n_278), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_307), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_308), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_312), .A2(n_281), .B(n_285), .Y(n_345) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_263), .B(n_253), .Y(n_346) );
OAI21x1_ASAP7_75t_SL g347 ( .A1(n_335), .A2(n_282), .B(n_267), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_289), .A2(n_283), .B(n_256), .Y(n_348) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_311), .B(n_272), .C(n_328), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_314), .A2(n_234), .B(n_226), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
NAND2x1_ASAP7_75t_L g352 ( .A(n_296), .B(n_242), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_332), .A2(n_266), .B(n_252), .Y(n_353) );
AO31x2_ASAP7_75t_L g354 ( .A1(n_315), .A2(n_280), .A3(n_287), .B(n_288), .Y(n_354) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_302), .A2(n_277), .B(n_244), .Y(n_355) );
AO21x1_ASAP7_75t_L g356 ( .A1(n_319), .A2(n_284), .B(n_229), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_329), .A2(n_229), .A3(n_262), .B(n_274), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_340), .A2(n_249), .B(n_259), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_323), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g360 ( .A1(n_320), .A2(n_264), .B(n_255), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_301), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_299), .B(n_242), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_313), .B(n_95), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_324), .B(n_97), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_325), .A2(n_99), .B(n_101), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_309), .B(n_102), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_297), .B(n_103), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_293), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_321), .B(n_105), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_294), .B(n_107), .C(n_108), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_304), .A2(n_291), .B(n_305), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_295), .B(n_318), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_325), .B(n_316), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_341), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_365), .Y(n_376) );
AO32x2_ASAP7_75t_L g377 ( .A1(n_356), .A2(n_337), .A3(n_298), .B1(n_338), .B2(n_331), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_369), .B(n_336), .Y(n_378) );
OAI21xp5_ASAP7_75t_L g379 ( .A1(n_349), .A2(n_292), .B(n_290), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_330), .B(n_326), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_359), .B(n_303), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_355), .A2(n_336), .B1(n_306), .B2(n_295), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_342), .A2(n_317), .B(n_322), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_351), .B(n_310), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_344), .A2(n_333), .B1(n_301), .B2(n_334), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_362), .B(n_367), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_361), .B(n_344), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_341), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_367), .B(n_364), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_342), .A2(n_372), .B(n_366), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_366), .A2(n_350), .B(n_356), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_373), .A2(n_361), .B1(n_360), .B2(n_343), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g395 ( .A(n_351), .B(n_343), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_346), .A2(n_348), .B(n_363), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_353), .A2(n_368), .B(n_363), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_347), .A2(n_368), .B1(n_358), .B2(n_371), .Y(n_400) );
OAI21x1_ASAP7_75t_L g401 ( .A1(n_352), .A2(n_358), .B(n_357), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_358), .A2(n_302), .B1(n_189), .B2(n_324), .Y(n_402) );
OA21x2_ASAP7_75t_L g403 ( .A1(n_357), .A2(n_356), .B(n_342), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_385), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_385), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_389), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_389), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_393), .A2(n_357), .B(n_354), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_389), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_392), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_396), .Y(n_416) );
OAI21x1_ASAP7_75t_L g417 ( .A1(n_393), .A2(n_357), .B(n_354), .Y(n_417) );
AO21x2_ASAP7_75t_L g418 ( .A1(n_397), .A2(n_354), .B(n_401), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_401), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_403), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
AO31x2_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_354), .A3(n_391), .B(n_396), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_383), .Y(n_424) );
INVx11_ASAP7_75t_L g425 ( .A(n_375), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_395), .Y(n_426) );
INVx4_ASAP7_75t_L g427 ( .A(n_383), .Y(n_427) );
AO21x2_ASAP7_75t_L g428 ( .A1(n_379), .A2(n_374), .B(n_399), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
OAI21x1_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_374), .B(n_380), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_395), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_384), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_386), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_402), .A2(n_388), .B1(n_398), .B2(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_380), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_386), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_377), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_390), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_378), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_377), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_387), .A2(n_302), .B1(n_369), .B2(n_324), .Y(n_446) );
OAI21x1_ASAP7_75t_L g447 ( .A1(n_377), .A2(n_393), .B(n_392), .Y(n_447) );
AOI21x1_ASAP7_75t_L g448 ( .A1(n_377), .A2(n_403), .B(n_356), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
BUFx2_ASAP7_75t_L g450 ( .A(n_416), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_405), .B(n_411), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_405), .B(n_411), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_419), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_416), .B(n_414), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_427), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_410), .B(n_414), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_421), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_410), .B(n_406), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_426), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_423), .B(n_406), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_421), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_421), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_431), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_425), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_431), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_423), .B(n_441), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_443), .B(n_435), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_423), .B(n_441), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_420), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_427), .Y(n_476) );
BUFx12f_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
AOI222xp33_ASAP7_75t_L g478 ( .A1(n_435), .A2(n_443), .B1(n_446), .B2(n_445), .C1(n_442), .C2(n_444), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_446), .A2(n_443), .B1(n_445), .B2(n_442), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_438), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_438), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_420), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_408), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_438), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_423), .B(n_441), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_433), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_427), .B(n_426), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_423), .B(n_443), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_409), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_439), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_426), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_426), .B(n_434), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_443), .B(n_425), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_442), .B(n_409), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_434), .B(n_436), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_422), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_422), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_442), .B(n_409), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_423), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_442), .B(n_413), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_413), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_423), .B(n_444), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_423), .B(n_418), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_440), .B(n_418), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_429), .Y(n_513) );
OR2x2_ASAP7_75t_SL g514 ( .A(n_436), .B(n_445), .Y(n_514) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_429), .B(n_432), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_429), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_432), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_418), .B(n_412), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_424), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_432), .B(n_418), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_424), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_418), .B(n_412), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_424), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_449), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_450), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_457), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_467), .A2(n_424), .B1(n_407), .B2(n_415), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_461), .B(n_424), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_489), .B(n_428), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_450), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_461), .B(n_412), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_501), .B(n_417), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_501), .B(n_417), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_452), .B(n_417), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_471), .B(n_428), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_501), .B(n_428), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_452), .B(n_448), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_476), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_449), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_457), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_454), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_460), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
AND2x4_ASAP7_75t_SL g546 ( .A(n_497), .B(n_495), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_501), .B(n_428), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_468), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_459), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_455), .B(n_463), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_451), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_455), .B(n_428), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_453), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_470), .B(n_448), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_470), .B(n_448), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_465), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_472), .B(n_447), .Y(n_559) );
INVx5_ASAP7_75t_L g560 ( .A(n_477), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_495), .B(n_447), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_502), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_503), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_489), .B(n_430), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g566 ( .A(n_477), .B(n_407), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_463), .B(n_447), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_478), .A2(n_407), .B(n_415), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_465), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_474), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_482), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_479), .B(n_472), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_482), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_467), .A2(n_415), .B1(n_430), .B2(n_437), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_513), .B(n_430), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_490), .B(n_492), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_487), .B(n_507), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_476), .B(n_491), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_483), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_459), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_490), .B(n_506), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_469), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_495), .B(n_509), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_487), .B(n_507), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_483), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_495), .B(n_516), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_469), .Y(n_587) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_464), .Y(n_588) );
BUFx2_ASAP7_75t_L g589 ( .A(n_516), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_464), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_473), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_473), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_516), .B(n_485), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_466), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_484), .B(n_493), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_476), .B(n_491), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_458), .B(n_462), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_484), .B(n_493), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_511), .B(n_458), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_511), .B(n_458), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_456), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_458), .B(n_510), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_498), .Y(n_603) );
INVx5_ASAP7_75t_L g604 ( .A(n_476), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_466), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_480), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_504), .B(n_508), .Y(n_607) );
INVx4_ASAP7_75t_L g608 ( .A(n_456), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_480), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_481), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_523), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_462), .B(n_517), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_510), .B(n_522), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_462), .B(n_517), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_481), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_515), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_515), .Y(n_617) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_486), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_486), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_515), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_518), .B(n_522), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_604), .B(n_491), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_621), .B(n_518), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_621), .B(n_520), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_594), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_524), .Y(n_626) );
OAI21xp5_ASAP7_75t_L g627 ( .A1(n_560), .A2(n_521), .B(n_456), .Y(n_627) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_608), .B(n_491), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_541), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_594), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_572), .A2(n_512), .B1(n_519), .B2(n_494), .C(n_499), .Y(n_631) );
BUFx2_ASAP7_75t_L g632 ( .A(n_608), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_605), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_605), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_551), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_596), .B(n_494), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_613), .B(n_494), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_556), .B(n_512), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_550), .B(n_514), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_546), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_556), .B(n_488), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_557), .B(n_488), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_599), .B(n_514), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_557), .B(n_496), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_559), .B(n_496), .Y(n_645) );
NOR2x1p5_ASAP7_75t_L g646 ( .A(n_608), .B(n_519), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_559), .B(n_499), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_532), .B(n_500), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_577), .B(n_500), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_596), .B(n_519), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_554), .B(n_505), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_589), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_584), .B(n_505), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_555), .B(n_603), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_600), .B(n_538), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_602), .B(n_576), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_547), .B(n_561), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_533), .B(n_534), .Y(n_658) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_568), .A2(n_581), .B1(n_536), .B2(n_531), .C(n_537), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_528), .B(n_567), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_526), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_607), .B(n_598), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_562), .Y(n_663) );
OR2x6_ASAP7_75t_L g664 ( .A(n_566), .B(n_578), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_563), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_583), .B(n_597), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_564), .Y(n_667) );
AND2x4_ASAP7_75t_SL g668 ( .A(n_616), .B(n_586), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_593), .B(n_548), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_548), .B(n_614), .Y(n_670) );
AND2x4_ASAP7_75t_SL g671 ( .A(n_612), .B(n_596), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_570), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_546), .B(n_525), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_525), .B(n_530), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_535), .B(n_539), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_595), .B(n_543), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_571), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_573), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_542), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_543), .B(n_580), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_545), .B(n_580), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_545), .B(n_549), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_588), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_588), .B(n_590), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_544), .B(n_582), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_579), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_578), .B(n_601), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
NAND2x1_ASAP7_75t_L g689 ( .A(n_540), .B(n_529), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_560), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_544), .B(n_582), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_530), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_531), .B(n_536), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_604), .B(n_540), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_552), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_611), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_617), .B(n_620), .Y(n_697) );
OR2x2_ASAP7_75t_L g698 ( .A(n_553), .B(n_587), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_552), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_604), .B(n_540), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_558), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_604), .B(n_591), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_558), .B(n_591), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_569), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_569), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_587), .B(n_592), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_592), .B(n_606), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_606), .B(n_609), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_609), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_575), .B(n_618), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_610), .B(n_615), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_610), .B(n_615), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_619), .B(n_565), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_560), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_619), .B(n_565), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_560), .B(n_574), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_574), .B(n_527), .Y(n_717) );
OAI221xp5_ASAP7_75t_SL g718 ( .A1(n_572), .A2(n_479), .B1(n_435), .B2(n_478), .C(n_402), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_524), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_646), .B(n_671), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_675), .B(n_638), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_675), .B(n_638), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_658), .B(n_660), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_624), .B(n_692), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_624), .B(n_649), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_649), .B(n_653), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_653), .B(n_623), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_658), .B(n_660), .Y(n_728) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_680), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_681), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_683), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_623), .B(n_682), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_676), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_662), .B(n_656), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_696), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_654), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_684), .Y(n_737) );
AND2x4_ASAP7_75t_L g738 ( .A(n_671), .B(n_628), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_682), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_686), .B(n_688), .Y(n_740) );
INVx2_ASAP7_75t_SL g741 ( .A(n_668), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_652), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_626), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_628), .B(n_668), .Y(n_744) );
INVx2_ASAP7_75t_SL g745 ( .A(n_714), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_629), .Y(n_746) );
OR2x2_ASAP7_75t_L g747 ( .A(n_637), .B(n_655), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_622), .A2(n_690), .B(n_632), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_666), .B(n_669), .Y(n_749) );
INVx1_ASAP7_75t_SL g750 ( .A(n_640), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_635), .Y(n_751) );
NAND2xp67_ASAP7_75t_SL g752 ( .A(n_717), .B(n_700), .Y(n_752) );
AND2x4_ASAP7_75t_L g753 ( .A(n_694), .B(n_636), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_641), .B(n_642), .Y(n_754) );
INVx2_ASAP7_75t_L g755 ( .A(n_710), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_714), .B(n_687), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_641), .B(n_642), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_710), .Y(n_758) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_710), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_670), .B(n_657), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_657), .B(n_655), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_673), .B(n_674), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_644), .B(n_719), .Y(n_763) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_664), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_698), .B(n_645), .Y(n_765) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_636), .B(n_697), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g767 ( .A1(n_664), .A2(n_639), .B1(n_622), .B2(n_643), .Y(n_767) );
AND2x4_ASAP7_75t_SL g768 ( .A(n_636), .B(n_694), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_644), .B(n_678), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_663), .B(n_665), .Y(n_770) );
INVxp67_ASAP7_75t_L g771 ( .A(n_693), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_647), .B(n_648), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_667), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_694), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_672), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_677), .Y(n_776) );
AND2x4_ASAP7_75t_SL g777 ( .A(n_664), .B(n_650), .Y(n_777) );
INVxp67_ASAP7_75t_SL g778 ( .A(n_702), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_648), .Y(n_779) );
INVx3_ASAP7_75t_L g780 ( .A(n_689), .Y(n_780) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_685), .Y(n_781) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_707), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_643), .B(n_650), .Y(n_783) );
OR2x6_ASAP7_75t_L g784 ( .A(n_627), .B(n_716), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_650), .B(n_713), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_717), .A2(n_631), .B1(n_715), .B2(n_713), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_651), .Y(n_787) );
AND2x4_ASAP7_75t_L g788 ( .A(n_715), .B(n_691), .Y(n_788) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_699), .B(n_704), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_740), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_764), .A2(n_718), .B1(n_659), .B2(n_708), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_789), .Y(n_792) );
AOI21xp33_ASAP7_75t_SL g793 ( .A1(n_767), .A2(n_701), .B(n_630), .Y(n_793) );
OAI21xp5_ASAP7_75t_SL g794 ( .A1(n_744), .A2(n_712), .B(n_711), .Y(n_794) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_748), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_729), .B(n_712), .Y(n_796) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_748), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_744), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_756), .A2(n_711), .B(n_706), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_740), .Y(n_800) );
AND2x2_ASAP7_75t_L g801 ( .A(n_788), .B(n_783), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_770), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_788), .B(n_703), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_723), .B(n_706), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_742), .A2(n_625), .B(n_630), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_782), .B(n_625), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_770), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_721), .B(n_633), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_721), .B(n_633), .Y(n_809) );
OAI21xp33_ASAP7_75t_L g810 ( .A1(n_786), .A2(n_634), .B(n_661), .Y(n_810) );
INVx2_ASAP7_75t_SL g811 ( .A(n_738), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_763), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_728), .B(n_634), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_771), .A2(n_679), .B1(n_695), .B2(n_705), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_722), .B(n_679), .Y(n_815) );
NAND2x1_ASAP7_75t_L g816 ( .A(n_738), .B(n_709), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_763), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_769), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_779), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_722), .B(n_709), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_769), .Y(n_821) );
AND2x2_ASAP7_75t_L g822 ( .A(n_762), .B(n_695), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_787), .B(n_705), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_733), .B(n_736), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_781), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_726), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_742), .B(n_771), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_727), .B(n_725), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_726), .Y(n_829) );
INVx2_ASAP7_75t_SL g830 ( .A(n_766), .Y(n_830) );
AO21x1_ASAP7_75t_SL g831 ( .A1(n_759), .A2(n_732), .B(n_754), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_727), .B(n_725), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_741), .A2(n_720), .B1(n_750), .B2(n_777), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_724), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_750), .B(n_734), .Y(n_835) );
INVx1_ASAP7_75t_SL g836 ( .A(n_768), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_790), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_793), .A2(n_720), .B(n_774), .C(n_753), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_833), .A2(n_745), .B(n_778), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_800), .Y(n_840) );
OR2x2_ASAP7_75t_L g841 ( .A(n_828), .B(n_732), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_802), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_807), .B(n_761), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_806), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_831), .B(n_753), .Y(n_845) );
NAND4xp25_ASAP7_75t_L g846 ( .A(n_791), .B(n_780), .C(n_752), .D(n_735), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_812), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_798), .A2(n_784), .B1(n_747), .B2(n_785), .Y(n_848) );
OAI31xp33_ASAP7_75t_L g849 ( .A1(n_795), .A2(n_780), .A3(n_749), .B(n_760), .Y(n_849) );
INVxp67_ASAP7_75t_L g850 ( .A(n_835), .Y(n_850) );
XNOR2x1_ASAP7_75t_L g851 ( .A(n_836), .B(n_784), .Y(n_851) );
BUFx6f_ASAP7_75t_L g852 ( .A(n_816), .Y(n_852) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_798), .A2(n_784), .B1(n_757), .B2(n_754), .Y(n_853) );
OAI22xp5_ASAP7_75t_SL g854 ( .A1(n_811), .A2(n_785), .B1(n_758), .B2(n_755), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_817), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_826), .B(n_724), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_818), .Y(n_857) );
NAND3xp33_ASAP7_75t_SL g858 ( .A(n_794), .B(n_757), .C(n_765), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_821), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_819), .Y(n_860) );
INVx1_ASAP7_75t_SL g861 ( .A(n_830), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_829), .B(n_834), .Y(n_862) );
OAI31xp33_ASAP7_75t_L g863 ( .A1(n_810), .A2(n_795), .A3(n_797), .B(n_798), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_823), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_844), .B(n_850), .Y(n_865) );
NAND2xp33_ASAP7_75t_L g866 ( .A(n_838), .B(n_811), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_864), .B(n_797), .Y(n_867) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_863), .B(n_827), .C(n_835), .D(n_799), .Y(n_868) );
OAI22xp5_ASAP7_75t_SL g869 ( .A1(n_854), .A2(n_830), .B1(n_827), .B2(n_792), .Y(n_869) );
AOI322xp5_ASAP7_75t_L g870 ( .A1(n_858), .A2(n_832), .A3(n_804), .B1(n_824), .B2(n_819), .C1(n_796), .C2(n_813), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_862), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g872 ( .A1(n_839), .A2(n_792), .B(n_825), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_861), .B(n_801), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_851), .A2(n_805), .B(n_825), .Y(n_874) );
O2A1O1Ixp33_ASAP7_75t_L g875 ( .A1(n_846), .A2(n_808), .B(n_809), .C(n_751), .Y(n_875) );
OAI211xp5_ASAP7_75t_SL g876 ( .A1(n_849), .A2(n_814), .B(n_820), .C(n_815), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_837), .Y(n_877) );
OAI21xp33_ASAP7_75t_L g878 ( .A1(n_853), .A2(n_730), .B(n_731), .Y(n_878) );
NOR3xp33_ASAP7_75t_L g879 ( .A(n_848), .B(n_854), .C(n_840), .Y(n_879) );
BUFx6f_ASAP7_75t_L g880 ( .A(n_865), .Y(n_880) );
AOI211xp5_ASAP7_75t_L g881 ( .A1(n_869), .A2(n_849), .B(n_852), .C(n_845), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g882 ( .A1(n_866), .A2(n_852), .B(n_842), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_868), .A2(n_852), .B(n_859), .Y(n_883) );
OA21x2_ASAP7_75t_L g884 ( .A1(n_872), .A2(n_860), .B(n_857), .Y(n_884) );
BUFx2_ASAP7_75t_L g885 ( .A(n_871), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_873), .B(n_841), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_877), .Y(n_887) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_882), .B(n_875), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_886), .B(n_870), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_881), .A2(n_874), .B1(n_879), .B2(n_867), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_885), .Y(n_891) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_880), .B(n_876), .C(n_878), .Y(n_892) );
AND2x4_ASAP7_75t_L g893 ( .A(n_891), .B(n_880), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_892), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_889), .B(n_880), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_893), .Y(n_896) );
NOR2xp67_ASAP7_75t_L g897 ( .A(n_894), .B(n_883), .Y(n_897) );
NOR2x1_ASAP7_75t_L g898 ( .A(n_895), .B(n_888), .Y(n_898) );
INVx3_ASAP7_75t_SL g899 ( .A(n_896), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_898), .B(n_890), .Y(n_900) );
AOI22x1_ASAP7_75t_L g901 ( .A1(n_899), .A2(n_897), .B1(n_887), .B2(n_884), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_900), .B(n_884), .Y(n_902) );
INVx2_ASAP7_75t_SL g903 ( .A(n_901), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_902), .B(n_855), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_903), .A2(n_847), .B1(n_856), .B2(n_843), .C(n_746), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_905), .A2(n_904), .B(n_803), .Y(n_906) );
OA21x2_ASAP7_75t_L g907 ( .A1(n_906), .A2(n_773), .B(n_776), .Y(n_907) );
AOI31xp33_ASAP7_75t_L g908 ( .A1(n_907), .A2(n_737), .A3(n_775), .B(n_743), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g909 ( .A1(n_908), .A2(n_822), .B1(n_772), .B2(n_739), .Y(n_909) );
endmodule