module fake_jpeg_17977_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_11),
.Y(n_32)
);

INVx8_ASAP7_75t_SL g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_25),
.B1(n_27),
.B2(n_20),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_21),
.C(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_26),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_0),
.Y(n_49)
);

XOR2x1_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_20),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_53),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_63),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_31),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_28),
.B1(n_17),
.B2(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_84),
.Y(n_93)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_82),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_18),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_48),
.C(n_50),
.Y(n_98)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_87),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_61),
.B1(n_59),
.B2(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_17),
.B1(n_19),
.B2(n_30),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_49),
.B1(n_64),
.B2(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_47),
.B1(n_29),
.B2(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_38),
.B1(n_33),
.B2(n_23),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_52),
.B1(n_51),
.B2(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_29),
.B1(n_19),
.B2(n_33),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_85),
.B1(n_61),
.B2(n_57),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_78),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_106),
.B(n_87),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_57),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_108),
.B(n_15),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_81),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_110),
.B1(n_90),
.B2(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_82),
.A2(n_11),
.B1(n_1),
.B2(n_3),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_23),
.CI(n_22),
.CON(n_109),
.SN(n_109)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_23),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_68),
.C(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_116),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_106),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_88),
.C(n_72),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_131),
.C(n_140),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_141),
.B(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_80),
.B1(n_70),
.B2(n_85),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_77),
.B(n_76),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_137),
.B(n_139),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_95),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_109),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_84),
.C(n_81),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_143),
.B(n_149),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_163),
.B(n_119),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_128),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_152),
.C(n_117),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_93),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_106),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_162),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_127),
.B1(n_128),
.B2(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_103),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_106),
.B(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_74),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_120),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_118),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_170),
.C(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_146),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_158),
.B1(n_165),
.B2(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_R g173 ( 
.A1(n_163),
.A2(n_92),
.B(n_141),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_181),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_154),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_123),
.B1(n_133),
.B2(n_135),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_188),
.B1(n_183),
.B2(n_175),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_67),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_187),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_147),
.B1(n_157),
.B2(n_165),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_169),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_200),
.B1(n_205),
.B2(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_206),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_164),
.B1(n_115),
.B2(n_80),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_164),
.C(n_102),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_178),
.C(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_89),
.B1(n_148),
.B2(n_130),
.Y(n_208)
);

AOI321xp33_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_167),
.A3(n_170),
.B1(n_186),
.B2(n_188),
.C(n_179),
.Y(n_209)
);

OAI21x1_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_197),
.B(n_199),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_215),
.C(n_196),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_178),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_189),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_172),
.C(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_219),
.C(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_194),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_184),
.C(n_174),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_174),
.B1(n_1),
.B2(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_220),
.B(n_205),
.Y(n_225)
);

AO22x2_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_21),
.B1(n_0),
.B2(n_5),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_224),
.A2(n_231),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_208),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_229),
.B(n_230),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_222),
.C(n_212),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_234),
.A2(n_221),
.B(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_217),
.B1(n_218),
.B2(n_0),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_241),
.B1(n_9),
.B2(n_10),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_21),
.B1(n_6),
.B2(n_7),
.Y(n_241)
);

AOI31xp33_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_4),
.A3(n_6),
.B(n_7),
.Y(n_243)
);

OAI21x1_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_4),
.B(n_7),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_232),
.B(n_6),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_9),
.B(n_12),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_251),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_8),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_12),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_240),
.C(n_10),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_16),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_254),
.B(n_255),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_238),
.C(n_11),
.Y(n_254)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_245),
.B(n_250),
.C(n_16),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_257),
.B(n_13),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_13),
.B(n_14),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_13),
.B(n_14),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_261),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule