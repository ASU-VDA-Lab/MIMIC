module real_jpeg_19567_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_341, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_341;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_0),
.A2(n_23),
.B1(n_26),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_121),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_121),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_1),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_14),
.B(n_48),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_119),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_94),
.B1(n_175),
.B2(n_176),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_1),
.B(n_76),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_30),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_1),
.A2(n_30),
.B(n_204),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_114),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_114),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_114),
.Y(n_193)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_4),
.Y(n_95)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_128),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_25),
.B1(n_42),
.B2(n_43),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_25),
.B1(n_47),
.B2(n_48),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_58),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_11),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_116),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_116),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_116),
.Y(n_254)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_338),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_82),
.B(n_336),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_20),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_21),
.A2(n_54),
.B(n_254),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_22),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_338)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_28),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_23),
.B(n_119),
.CON(n_118),
.SN(n_118)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_32),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_27),
.A2(n_34),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_30),
.Y(n_125)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_29),
.A2(n_35),
.B1(n_118),
.B2(n_125),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_29),
.A2(n_42),
.A3(n_66),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_30),
.A2(n_64),
.B(n_65),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_31),
.A2(n_55),
.B(n_59),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_34),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_37),
.B(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_74),
.C(n_78),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_38),
.A2(n_39),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_52),
.C(n_60),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_40),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_40),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_40),
.A2(n_60),
.B1(n_61),
.B2(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_46),
.B(n_50),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_41),
.A2(n_50),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_41),
.A2(n_46),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_41),
.A2(n_46),
.B1(n_171),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_41),
.A2(n_46),
.B1(n_193),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_41),
.A2(n_211),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_41),
.A2(n_46),
.B1(n_101),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_41),
.A2(n_109),
.B(n_246),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_43),
.A2(n_49),
.B(n_119),
.C(n_167),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_43),
.B(n_65),
.Y(n_205)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_46),
.B(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_47),
.B(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_51),
.B(n_110),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_52),
.A2(n_53),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_54),
.A2(n_59),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_54),
.A2(n_59),
.B1(n_134),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_54),
.A2(n_81),
.B(n_300),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_59),
.B(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_68),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_69),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_70),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_64),
.A2(n_70),
.B1(n_113),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_64),
.A2(n_70),
.B1(n_146),
.B2(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_64),
.B(n_73),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_64),
.A2(n_68),
.B(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_64),
.A2(n_70),
.B1(n_271),
.B2(n_292),
.Y(n_291)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_69),
.A2(n_77),
.B(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_69),
.A2(n_257),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_78),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_329),
.B(n_335),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_305),
.A3(n_324),
.B1(n_327),
.B2(n_328),
.C(n_341),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_284),
.B(n_304),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_262),
.B(n_283),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_151),
.B(n_236),
.C(n_261),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_139),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_88),
.B(n_139),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_122),
.B2(n_138),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_106),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_91),
.B(n_106),
.C(n_138),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_100),
.B2(n_105),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_92),
.B(n_105),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_94),
.A2(n_96),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_99),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_94),
.A2(n_161),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_94),
.A2(n_163),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_94),
.A2(n_95),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_119),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_98),
.A2(n_159),
.B(n_196),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_102),
.B(n_227),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_117),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_123),
.B(n_131),
.C(n_136),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_140),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_145),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_147),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_235),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_229),
.B(n_234),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_216),
.B(n_228),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_198),
.B(n_215),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_185),
.B(n_197),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_172),
.B(n_184),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_168),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_179),
.B(n_183),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_178),
.Y(n_183)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_187),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_196),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_206),
.B1(n_213),
.B2(n_214),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_201),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_207),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_218),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_225),
.C(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_237),
.B(n_238),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_259),
.B2(n_260),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_248),
.C(n_260),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_258),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_256),
.C(n_258),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_282),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_276),
.C(n_282),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_272),
.C(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_278),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_295),
.B(n_299),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_280),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_285),
.B(n_286),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_302),
.B2(n_303),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_289),
.B(n_294),
.C(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_292),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_307),
.C(n_316),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_293),
.B(n_307),
.CI(n_316),
.CON(n_326),
.SN(n_326)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_299),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_317),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_309),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_312),
.C(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_322),
.C(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_326),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);


endmodule