module fake_jpeg_10406_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx14_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_4),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_21),
.B(n_22),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_16),
.C(n_15),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_13),
.B(n_11),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.C(n_7),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_21),
.B(n_12),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_14),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_33),
.C(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_14),
.B2(n_9),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_8),
.B(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_3),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B(n_8),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_3),
.C(n_5),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_1),
.Y(n_40)
);


endmodule