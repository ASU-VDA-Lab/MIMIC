module fake_jpeg_11575_n_261 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_44),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_27),
.B(n_0),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_50),
.B(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_80),
.Y(n_104)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_3),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_20),
.B(n_3),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_30),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_24),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_72),
.Y(n_91)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_76),
.Y(n_118)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_5),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_13),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_26),
.B1(n_28),
.B2(n_41),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_84),
.A2(n_88),
.B1(n_96),
.B2(n_97),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_28),
.B1(n_41),
.B2(n_31),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_37),
.B1(n_32),
.B2(n_31),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_32),
.B1(n_38),
.B2(n_25),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_38),
.C(n_25),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_110),
.C(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_42),
.A2(n_24),
.B1(n_34),
.B2(n_19),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_104),
.B1(n_118),
.B2(n_54),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_104),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_19),
.B1(n_7),
.B2(n_9),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_19),
.B(n_48),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_59),
.C(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_126),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_7),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_130),
.B(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_152),
.Y(n_174)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_133),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_157),
.B(n_163),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_136),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_64),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_95),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_101),
.B(n_89),
.C(n_94),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_136),
.B(n_130),
.C(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_148),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_146),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_120),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_86),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_151),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_155),
.Y(n_185)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_86),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_111),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_157),
.B(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_164),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_87),
.B(n_119),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_128),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_148),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_171),
.B(n_188),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_162),
.B1(n_135),
.B2(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_180),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_162),
.B1(n_149),
.B2(n_165),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_158),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_157),
.B1(n_154),
.B2(n_160),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_147),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_132),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_172),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_142),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_201),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_208),
.B(n_166),
.Y(n_227)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_132),
.B(n_159),
.C(n_180),
.Y(n_207)
);

XNOR2x2_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_212),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_193),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_179),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_174),
.B(n_191),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_175),
.B1(n_182),
.B2(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_213),
.Y(n_223)
);

AOI221xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_183),
.B1(n_207),
.B2(n_196),
.C(n_176),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_169),
.B1(n_166),
.B2(n_192),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_212),
.B1(n_213),
.B2(n_203),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_176),
.B(n_197),
.C(n_181),
.D(n_202),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_227),
.A2(n_208),
.B(n_204),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_200),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_200),
.C(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_230),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_234),
.B1(n_236),
.B2(n_224),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_218),
.A2(n_194),
.B1(n_208),
.B2(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_237),
.B1(n_223),
.B2(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_194),
.C(n_188),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_240),
.A2(n_244),
.B(n_233),
.C(n_238),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_229),
.B1(n_228),
.B2(n_227),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_237),
.B(n_226),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_241),
.B(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_249),
.B1(n_241),
.B2(n_221),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_236),
.B1(n_222),
.B2(n_234),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_225),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_250),
.A2(n_252),
.B(n_168),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_251),
.A2(n_214),
.B1(n_221),
.B2(n_181),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_173),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_258),
.C(n_255),
.Y(n_260)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_260),
.B(n_173),
.CI(n_253),
.CON(n_261),
.SN(n_261)
);


endmodule