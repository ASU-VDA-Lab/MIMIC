module fake_netlist_1_9551_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_71), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_58), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_29), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_48), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_25), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_23), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_50), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_51), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_64), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_68), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_4), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_79), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_1), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
INVx2_ASAP7_75t_SL g97 ( .A(n_75), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_31), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_54), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_66), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_56), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_43), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_47), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_34), .Y(n_105) );
INVx2_ASAP7_75t_SL g106 ( .A(n_19), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
INVxp67_ASAP7_75t_SL g108 ( .A(n_15), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_33), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_61), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_57), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
NOR2xp67_ASAP7_75t_L g118 ( .A(n_52), .B(n_28), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_32), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_59), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_17), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_16), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_46), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_45), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_97), .B(n_1), .Y(n_126) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_80), .A2(n_35), .B(n_77), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_106), .B(n_2), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_113), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_81), .A2(n_36), .B(n_76), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_87), .B(n_3), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_108), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_86), .B(n_7), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_87), .B(n_8), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_111), .A2(n_121), .B1(n_102), .B2(n_117), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g142 ( .A1(n_92), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_97), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_112), .B(n_124), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_112), .B(n_9), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_81), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_101), .B(n_10), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_82), .B(n_41), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_94), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_95), .B(n_11), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_100), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_85), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_96), .B(n_11), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
BUFx8_ASAP7_75t_L g163 ( .A(n_98), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_143), .B(n_88), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_140), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_133), .A2(n_109), .B1(n_95), .B2(n_122), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_143), .B(n_110), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_129), .B(n_124), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_133), .B(n_137), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_133), .A2(n_109), .B1(n_122), .B2(n_107), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_134), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_152), .A2(n_107), .B1(n_116), .B2(n_117), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_163), .B(n_123), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_133), .A2(n_116), .B1(n_103), .B2(n_120), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_163), .B(n_89), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_143), .B(n_120), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_139), .B(n_103), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_152), .B(n_90), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_154), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_150), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_144), .B(n_114), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_135), .B(n_114), .Y(n_185) );
AND2x6_ASAP7_75t_L g186 ( .A(n_137), .B(n_105), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_131), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_163), .B(n_115), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_125), .B(n_105), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_137), .A2(n_99), .B1(n_98), .B2(n_93), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_125), .B(n_162), .Y(n_196) );
NAND2xp33_ASAP7_75t_L g197 ( .A(n_150), .B(n_99), .Y(n_197) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_150), .B(n_118), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_139), .A2(n_118), .B1(n_13), .B2(n_14), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_151), .B(n_12), .Y(n_200) );
AND3x2_ASAP7_75t_L g201 ( .A(n_156), .B(n_12), .C(n_13), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_157), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_146), .B(n_53), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_136), .B(n_18), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_129), .B(n_21), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_158), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_191), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_200), .B(n_157), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_179), .B(n_136), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_182), .B(n_148), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_179), .B(n_148), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_200), .B(n_128), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_182), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_196), .B(n_162), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_193), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
OR2x6_ASAP7_75t_L g223 ( .A(n_185), .B(n_135), .Y(n_223) );
INVx1_ASAP7_75t_SL g224 ( .A(n_187), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_178), .Y(n_225) );
BUFx12f_ASAP7_75t_L g226 ( .A(n_209), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_182), .B(n_160), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_203), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_178), .B(n_160), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_178), .B(n_159), .Y(n_231) );
AO22x1_ASAP7_75t_L g232 ( .A1(n_195), .A2(n_142), .B1(n_150), .B2(n_128), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_178), .B(n_146), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_185), .B(n_142), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_203), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_171), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_186), .B(n_159), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_169), .A2(n_153), .B1(n_147), .B2(n_150), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_145), .B(n_127), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_165), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_186), .B(n_153), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_169), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_186), .B(n_147), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_171), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_187), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_186), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_172), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_186), .B(n_145), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_165), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_164), .B(n_167), .Y(n_251) );
AND2x4_ASAP7_75t_L g252 ( .A(n_207), .B(n_170), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_186), .B(n_155), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_165), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_188), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_172), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_186), .B(n_155), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_173), .B(n_138), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_181), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_186), .A2(n_138), .B1(n_130), .B2(n_126), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_206), .B(n_141), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_169), .B(n_155), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_206), .B(n_140), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_175), .B(n_140), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_213), .A2(n_183), .B(n_192), .C(n_185), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_264), .A2(n_198), .B(n_183), .Y(n_269) );
XOR2xp5_ASAP7_75t_L g270 ( .A(n_260), .B(n_130), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_216), .A2(n_207), .B1(n_194), .B2(n_166), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_264), .A2(n_176), .B(n_174), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_252), .A2(n_202), .B1(n_199), .B2(n_185), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_215), .A2(n_192), .B(n_185), .C(n_168), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_229), .B(n_189), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_234), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_266), .A2(n_205), .B(n_204), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_218), .B(n_169), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_247), .B(n_181), .Y(n_281) );
NAND3xp33_ASAP7_75t_L g282 ( .A(n_239), .B(n_208), .C(n_205), .Y(n_282) );
AO32x2_ASAP7_75t_L g283 ( .A1(n_240), .A2(n_127), .A3(n_132), .B1(n_150), .B2(n_169), .Y(n_283) );
OAI22x1_ASAP7_75t_L g284 ( .A1(n_224), .A2(n_161), .B1(n_201), .B2(n_132), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_218), .B(n_169), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_252), .A2(n_204), .B1(n_169), .B2(n_190), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_211), .B(n_190), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_266), .A2(n_127), .B(n_132), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_225), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_249), .A2(n_127), .B(n_132), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_217), .B(n_184), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_218), .B(n_184), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_230), .A2(n_149), .B(n_188), .C(n_210), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_245), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_227), .A2(n_210), .B(n_188), .Y(n_296) );
NOR2xp33_ASAP7_75t_R g297 ( .A(n_226), .B(n_150), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_247), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_246), .B(n_210), .C(n_26), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_212), .Y(n_301) );
OAI22xp5_ASAP7_75t_SL g302 ( .A1(n_223), .A2(n_141), .B1(n_140), .B2(n_30), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_226), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_L g304 ( .A1(n_251), .A2(n_221), .B(n_222), .C(n_233), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_217), .B(n_243), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_267), .A2(n_141), .B(n_27), .C(n_37), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_252), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_227), .A2(n_141), .B(n_38), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_256), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_258), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_212), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_241), .Y(n_316) );
BUFx12f_ASAP7_75t_L g317 ( .A(n_223), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_269), .A2(n_239), .B(n_267), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_291), .A2(n_251), .B(n_214), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_268), .A2(n_262), .B(n_265), .C(n_244), .Y(n_320) );
AO31x2_ASAP7_75t_L g321 ( .A1(n_304), .A2(n_253), .A3(n_257), .B(n_238), .Y(n_321) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_276), .A2(n_242), .B(n_212), .Y(n_322) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_285), .B(n_235), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_275), .Y(n_324) );
AOI21xp5_ASAP7_75t_SL g325 ( .A1(n_304), .A2(n_263), .B(n_219), .Y(n_325) );
OAI22xp33_ASAP7_75t_L g326 ( .A1(n_273), .A2(n_235), .B1(n_223), .B2(n_214), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_271), .A2(n_235), .B1(n_219), .B2(n_228), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_288), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_289), .A2(n_241), .B(n_255), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_270), .A2(n_232), .B1(n_141), .B2(n_254), .C(n_250), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_278), .A2(n_263), .B(n_219), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_301), .B(n_263), .Y(n_332) );
OAI22x1_ASAP7_75t_L g333 ( .A1(n_303), .A2(n_255), .B1(n_254), .B2(n_250), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_SL g334 ( .A1(n_306), .A2(n_22), .B(n_40), .C(n_42), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_317), .A2(n_263), .B1(n_236), .B2(n_228), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_286), .A2(n_236), .B1(n_228), .B2(n_219), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_299), .A2(n_236), .B1(n_228), .B2(n_141), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_286), .A2(n_308), .B1(n_279), .B2(n_276), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_296), .A2(n_236), .B(n_49), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_274), .A2(n_44), .B(n_55), .C(n_60), .Y(n_342) );
A2O1A1Ixp33_ASAP7_75t_L g343 ( .A1(n_294), .A2(n_62), .B(n_63), .C(n_65), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_292), .A2(n_67), .B(n_69), .Y(n_344) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_300), .B(n_70), .C(n_72), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_275), .B(n_73), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_287), .A2(n_78), .B1(n_312), .B2(n_295), .Y(n_347) );
BUFx10_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_293), .A2(n_280), .B1(n_295), .B2(n_312), .Y(n_349) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_313), .A2(n_314), .B1(n_290), .B2(n_280), .C1(n_302), .C2(n_277), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_292), .A2(n_272), .B(n_282), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_277), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
OAI21xp33_ASAP7_75t_L g354 ( .A1(n_347), .A2(n_284), .B(n_297), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_323), .B(n_281), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_347), .A2(n_309), .B(n_311), .C(n_305), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_328), .B(n_298), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_348), .B(n_281), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_346), .B(n_298), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_341), .A2(n_316), .B(n_305), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_329), .A2(n_283), .B(n_297), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_348), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_283), .B1(n_311), .B2(n_350), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_319), .A2(n_283), .B(n_320), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_352), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_340), .B(n_283), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_322), .A2(n_327), .B1(n_335), .B2(n_330), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_346), .A2(n_332), .B1(n_333), .B2(n_324), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_325), .A2(n_351), .B(n_318), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g372 ( .A1(n_331), .A2(n_338), .B(n_342), .Y(n_372) );
INVxp33_ASAP7_75t_SL g373 ( .A(n_336), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_334), .A2(n_343), .B(n_345), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_324), .B(n_321), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_321), .B(n_352), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_321), .B(n_337), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_344), .A2(n_341), .B(n_329), .Y(n_378) );
AO31x2_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_319), .A3(n_304), .B(n_349), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_329), .A2(n_289), .B(n_351), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_380), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_353), .Y(n_383) );
NAND2xp33_ASAP7_75t_R g384 ( .A(n_360), .B(n_373), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_353), .Y(n_385) );
OAI31xp33_ASAP7_75t_L g386 ( .A1(n_373), .A2(n_354), .A3(n_358), .B(n_363), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_360), .B(n_367), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_360), .B(n_366), .Y(n_388) );
INVx5_ASAP7_75t_SL g389 ( .A(n_360), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_366), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_354), .B(n_359), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_381), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_381), .B(n_358), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_375), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_365), .A2(n_370), .B(n_378), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_363), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_359), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_376), .Y(n_398) );
AO21x2_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_377), .B(n_374), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_357), .B(n_369), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_366), .B(n_369), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_380), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_366), .B(n_371), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_362), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_368), .B(n_364), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
NAND2x1p5_ASAP7_75t_SL g415 ( .A(n_408), .B(n_355), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_389), .A2(n_363), .B1(n_356), .B2(n_355), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_393), .B(n_362), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_396), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_383), .B(n_361), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_386), .B(n_361), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_398), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_383), .B(n_378), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_393), .B(n_385), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_385), .B(n_392), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_382), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_392), .B(n_398), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_382), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_401), .B(n_402), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_400), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_400), .Y(n_435) );
OAI31xp33_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_403), .A3(n_386), .B(n_388), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_388), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_403), .B(n_402), .Y(n_440) );
AOI211xp5_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_401), .B(n_413), .C(n_388), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_413), .B(n_408), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_405), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_387), .B(n_408), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_405), .Y(n_445) );
AND2x4_ASAP7_75t_SL g446 ( .A(n_388), .B(n_409), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_410), .B(n_391), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_389), .A2(n_387), .B1(n_391), .B2(n_404), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_410), .B(n_389), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_410), .B(n_391), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_389), .A2(n_391), .B1(n_404), .B2(n_399), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
INVx4_ASAP7_75t_L g458 ( .A(n_421), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_428), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_423), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_425), .B(n_389), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_418), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_428), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_435), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_446), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_426), .B(n_409), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_435), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_422), .B(n_391), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_435), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_446), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_436), .A2(n_391), .B1(n_399), .B2(n_409), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_455), .B(n_399), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_399), .B1(n_409), .B2(n_395), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_417), .B(n_395), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_427), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_429), .B(n_395), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_422), .B(n_444), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_417), .B(n_395), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_416), .B(n_384), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_432), .B(n_395), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_432), .B(n_411), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_444), .B(n_411), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_414), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_414), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_440), .B(n_390), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_440), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_446), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_430), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_431), .B(n_390), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_442), .B(n_390), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_430), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_455), .B(n_390), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_442), .B(n_390), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_457), .B(n_390), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_457), .B(n_449), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_449), .B(n_448), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_433), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_433), .B(n_434), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_434), .B(n_443), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_439), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_448), .B(n_453), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_451), .B(n_453), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_451), .B(n_431), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_424), .Y(n_512) );
OR2x6_ASAP7_75t_L g513 ( .A(n_452), .B(n_416), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_437), .B(n_441), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_438), .B(n_445), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_459), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_501), .B(n_456), .Y(n_517) );
NOR2xp67_ASAP7_75t_SL g518 ( .A(n_468), .B(n_437), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_492), .A2(n_441), .B1(n_415), .B2(n_454), .C(n_450), .Y(n_519) );
INVx1_ASAP7_75t_SL g520 ( .A(n_464), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_483), .B(n_415), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_461), .Y(n_522) );
OR2x6_ASAP7_75t_L g523 ( .A(n_468), .B(n_513), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_467), .B(n_469), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_459), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_438), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_501), .B(n_438), .Y(n_527) );
INVx4_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_475), .Y(n_530) );
INVxp67_ASAP7_75t_SL g531 ( .A(n_459), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_489), .B(n_439), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_480), .B(n_454), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_474), .Y(n_534) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_485), .B(n_420), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_490), .B(n_445), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_502), .B(n_452), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_483), .B(n_447), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_511), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_460), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_495), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_470), .B(n_415), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_462), .B(n_424), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_458), .B(n_419), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_480), .B(n_445), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_458), .B(n_447), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_481), .B(n_447), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_458), .B(n_419), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_481), .B(n_505), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_484), .B(n_486), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_484), .B(n_486), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_515), .B(n_487), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_505), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_476), .A2(n_479), .B1(n_513), .B2(n_514), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_504), .B(n_509), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_510), .B(n_487), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_510), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_497), .B(n_508), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_515), .B(n_478), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_493), .A2(n_463), .B(n_472), .C(n_488), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_478), .B(n_482), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_493), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_513), .B(n_512), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_503), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_491), .B(n_503), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_478), .B(n_512), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_553), .B(n_513), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_553), .B(n_472), .Y(n_571) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_528), .A2(n_494), .B1(n_466), .B2(n_471), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_554), .B(n_500), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_534), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_554), .B(n_491), .Y(n_575) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_528), .B(n_465), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_540), .B(n_466), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_522), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_528), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_564), .B(n_533), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_529), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_564), .B(n_498), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_541), .Y(n_584) );
OA211x2_ASAP7_75t_L g585 ( .A1(n_557), .A2(n_499), .B(n_496), .C(n_495), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_556), .B(n_471), .Y(n_587) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_523), .B(n_473), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_517), .B(n_473), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_533), .B(n_498), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_562), .B(n_498), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_569), .B(n_500), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_517), .B(n_506), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_562), .B(n_500), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_544), .B(n_506), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_544), .B(n_507), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_551), .B(n_507), .Y(n_599) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_531), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_546), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g602 ( .A1(n_535), .A2(n_557), .B(n_520), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_563), .B(n_518), .C(n_566), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_527), .B(n_566), .Y(n_604) );
INVxp33_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_541), .Y(n_606) );
INVx2_ASAP7_75t_SL g607 ( .A(n_527), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_559), .B(n_558), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_552), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_565), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_547), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_527), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_547), .B(n_569), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
INVxp67_ASAP7_75t_SL g615 ( .A(n_600), .Y(n_615) );
OAI31xp33_ASAP7_75t_SL g616 ( .A1(n_603), .A2(n_542), .A3(n_545), .B(n_519), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_584), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_606), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_577), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_580), .B(n_555), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_602), .A2(n_523), .B1(n_543), .B2(n_521), .Y(n_621) );
AOI21xp33_ASAP7_75t_SL g622 ( .A1(n_603), .A2(n_579), .B(n_576), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g623 ( .A1(n_588), .A2(n_563), .B(n_560), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_578), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_580), .B(n_555), .Y(n_625) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_576), .A2(n_523), .B1(n_526), .B2(n_538), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_576), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_578), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_613), .B(n_516), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_572), .A2(n_524), .B1(n_568), .B2(n_539), .C(n_550), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_606), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_609), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_609), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_581), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_581), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_611), .B(n_537), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_579), .A2(n_561), .B1(n_532), .B2(n_567), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_613), .B(n_516), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_573), .B(n_525), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_611), .B(n_549), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_622), .A2(n_605), .B1(n_608), .B2(n_574), .C(n_570), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_616), .A2(n_570), .B(n_604), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_619), .B(n_571), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_636), .Y(n_644) );
O2A1O1Ixp5_ASAP7_75t_L g645 ( .A1(n_615), .A2(n_596), .B(n_598), .C(n_597), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_623), .B(n_588), .Y(n_646) );
OAI31xp33_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_610), .A3(n_596), .B(n_590), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_624), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_626), .A2(n_604), .B1(n_596), .B2(n_607), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_637), .A2(n_610), .B(n_596), .C(n_607), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_628), .Y(n_651) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_621), .A2(n_612), .B1(n_587), .B2(n_599), .C(n_589), .Y(n_652) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_627), .A2(n_612), .B(n_585), .C(n_593), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_620), .B(n_571), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_627), .B(n_601), .C(n_586), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_625), .B(n_575), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g657 ( .A1(n_645), .A2(n_604), .B(n_636), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_646), .B(n_640), .Y(n_658) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_647), .A2(n_640), .B(n_635), .C(n_634), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_649), .B(n_639), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_642), .A2(n_573), .B(n_575), .C(n_593), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_649), .B(n_585), .C(n_593), .D(n_594), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g663 ( .A1(n_641), .A2(n_633), .B(n_631), .C(n_632), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_650), .A2(n_631), .B(n_633), .Y(n_664) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_652), .A2(n_614), .B1(n_632), .B2(n_601), .C1(n_586), .C2(n_582), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_661), .A2(n_653), .B(n_655), .C(n_644), .Y(n_666) );
OR3x1_ASAP7_75t_L g667 ( .A(n_662), .B(n_656), .C(n_648), .Y(n_667) );
AOI21x1_ASAP7_75t_L g668 ( .A1(n_658), .A2(n_651), .B(n_643), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_659), .B(n_614), .C(n_617), .Y(n_669) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_657), .B(n_654), .C(n_593), .D(n_583), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_667), .A2(n_660), .B1(n_664), .B2(n_663), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_669), .Y(n_672) );
NOR2x1p5_ASAP7_75t_L g673 ( .A(n_670), .B(n_665), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_666), .B1(n_668), .B2(n_638), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_672), .B(n_617), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_675), .Y(n_676) );
OAI22xp5_ASAP7_75t_SL g677 ( .A1(n_674), .A2(n_671), .B1(n_618), .B2(n_582), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_676), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_678), .A2(n_677), .B(n_618), .Y(n_679) );
AOI22x1_ASAP7_75t_L g680 ( .A1(n_679), .A2(n_638), .B1(n_629), .B2(n_639), .Y(n_680) );
OAI21x1_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_629), .B(n_583), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_681), .A2(n_595), .B1(n_592), .B2(n_591), .Y(n_682) );
endmodule