module real_jpeg_24280_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_4),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_16),
.B1(n_34),
.B2(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_4),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_4),
.B(n_14),
.C(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_4),
.B(n_20),
.C(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_4),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_4),
.B(n_88),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_67),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_65),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_52),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_11),
.B(n_52),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_27),
.B(n_38),
.C(n_49),
.Y(n_11)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_12),
.A2(n_51),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_51),
.B1(n_71),
.B2(n_72),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_12),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_18),
.Y(n_12)
);

INVx5_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_14),
.B(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx3_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_23),
.B(n_84),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_37),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_34),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_38),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_48),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_48),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_39),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_39),
.B(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_51),
.C(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_92),
.B(n_98),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_80),
.B(n_91),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_70),
.B(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);


endmodule