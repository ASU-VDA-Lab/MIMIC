module fake_jpeg_14318_n_30 (n_3, n_2, n_1, n_0, n_4, n_5, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_5),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_16),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_9),
.B1(n_10),
.B2(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_20),
.B(n_15),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.C(n_17),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_26),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_18),
.C(n_13),
.Y(n_26)
);

AOI322xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_10),
.A3(n_19),
.B1(n_4),
.B2(n_5),
.C1(n_1),
.C2(n_2),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_10),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_10),
.Y(n_30)
);


endmodule