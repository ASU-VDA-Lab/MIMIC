module fake_jpeg_17246_n_149 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_2),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_65),
.Y(n_81)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_60),
.B1(n_53),
.B2(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_58),
.B1(n_56),
.B2(n_44),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_1),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_60),
.B1(n_58),
.B2(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_102),
.B1(n_81),
.B2(n_4),
.Y(n_105)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_100),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_48),
.B1(n_55),
.B2(n_52),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_98),
.B(n_8),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_55),
.B1(n_45),
.B2(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_23),
.B1(n_41),
.B2(n_40),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_107),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_10),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_7),
.B(n_8),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_112),
.B(n_98),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_103),
.B1(n_109),
.B2(n_104),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_93),
.C(n_89),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_94),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_120),
.B1(n_119),
.B2(n_121),
.Y(n_130)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_132),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_88),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_86),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_107),
.B1(n_104),
.B2(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_128),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.C(n_136),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_131),
.C(n_85),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_12),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_15),
.A3(n_17),
.B1(n_19),
.B2(n_21),
.C1(n_24),
.C2(n_25),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_28),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_29),
.B(n_30),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_31),
.C(n_32),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_33),
.C(n_35),
.Y(n_149)
);


endmodule