module fake_netlist_6_1299_n_992 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_992);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_992;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_742;
wire n_532;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_663;
wire n_361;
wire n_508;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_101),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_80),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_63),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_100),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_20),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_56),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_92),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_189),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_155),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_73),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_16),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_139),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_91),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_4),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_25),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_48),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_40),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_109),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_13),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_54),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_136),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_140),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_112),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_74),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_37),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_99),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_113),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_13),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_149),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_69),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_12),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_176),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_130),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_161),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_111),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_177),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_95),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_191),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_5),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_77),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_158),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_55),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_135),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_173),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_82),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_107),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_31),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_123),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_227),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_210),
.B(n_204),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_250),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_36),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

BUFx8_ASAP7_75t_SL g287 ( 
.A(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_194),
.B(n_38),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_209),
.B(n_0),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_0),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_215),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_1),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_241),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_2),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_2),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_194),
.B(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_214),
.B(n_4),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_225),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_193),
.B(n_5),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_214),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_239),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_7),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_7),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_8),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_199),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_8),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_216),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_237),
.B(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_200),
.B(n_9),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_230),
.B(n_10),
.Y(n_321)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_230),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_220),
.B(n_10),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_201),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_203),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_207),
.B(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_247),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_192),
.B1(n_195),
.B2(n_228),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_319),
.A2(n_192),
.B1(n_195),
.B2(n_248),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_281),
.A2(n_258),
.B1(n_264),
.B2(n_271),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_257),
.B1(n_222),
.B2(n_273),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_291),
.Y(n_335)
);

OR2x6_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_276),
.Y(n_336)
);

AO22x2_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_224),
.B1(n_226),
.B2(n_233),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_12),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_290),
.A2(n_235),
.B1(n_236),
.B2(n_242),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_307),
.B1(n_311),
.B2(n_306),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_196),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_329),
.A2(n_246),
.B1(n_253),
.B2(n_266),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_197),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_267),
.Y(n_345)
);

AO22x1_ASAP7_75t_L g346 ( 
.A1(n_293),
.A2(n_275),
.B1(n_269),
.B2(n_268),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_265),
.B1(n_263),
.B2(n_262),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_287),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_292),
.B(n_198),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_296),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_293),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_261),
.B1(n_260),
.B2(n_256),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_289),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_294),
.A2(n_255),
.B1(n_254),
.B2(n_252),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_290),
.A2(n_251),
.B1(n_249),
.B2(n_244),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_279),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_202),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_329),
.A2(n_243),
.B1(n_240),
.B2(n_234),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_305),
.A2(n_231),
.B1(n_229),
.B2(n_221),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_205),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_290),
.B(n_206),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_287),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_301),
.A2(n_318),
.B1(n_317),
.B2(n_322),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_289),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_285),
.A2(n_298),
.B1(n_304),
.B2(n_312),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_208),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_301),
.B(n_211),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_301),
.A2(n_317),
.B1(n_318),
.B2(n_322),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_213),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_317),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_317),
.B(n_217),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_L g375 ( 
.A1(n_317),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_318),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_318),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_279),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_302),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_322),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_292),
.B(n_19),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_39),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_285),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g385 ( 
.A1(n_295),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_356),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_292),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_322),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_358),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_288),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_344),
.A2(n_303),
.B(n_300),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_333),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_330),
.B(n_302),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_347),
.B(n_320),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_331),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_328),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_348),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_370),
.A2(n_280),
.B(n_278),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_338),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_349),
.B(n_298),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_353),
.B(n_310),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_360),
.B(n_295),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_353),
.B(n_304),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_334),
.B(n_284),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_337),
.Y(n_421)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_383),
.B(n_300),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

XNOR2x2_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_309),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_41),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_355),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_370),
.A2(n_303),
.B(n_284),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_368),
.B(n_43),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

BUFx6f_ASAP7_75t_SL g433 ( 
.A(n_336),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_374),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_324),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_351),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_346),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_373),
.B(n_277),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_385),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_381),
.B(n_309),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_362),
.B(n_323),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_357),
.B(n_324),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_340),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_336),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_336),
.B(n_323),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

AND2x6_ASAP7_75t_SL g455 ( 
.A(n_345),
.B(n_315),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_345),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_345),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_334),
.B(n_277),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_371),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_420),
.B(n_310),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_327),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_422),
.B(n_357),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_310),
.Y(n_464)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_458),
.B(n_310),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_418),
.B(n_327),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_327),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_310),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_395),
.B(n_324),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_399),
.A2(n_375),
.B1(n_326),
.B2(n_324),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_427),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_324),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_399),
.B(n_326),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_417),
.B(n_326),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_458),
.B(n_277),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_410),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_326),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_410),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_459),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_401),
.B(n_326),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_452),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_401),
.B(n_279),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_284),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_449),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_436),
.B(n_375),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_436),
.B(n_278),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_389),
.B(n_279),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_284),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_421),
.B(n_284),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_429),
.A2(n_284),
.B(n_283),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_387),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_388),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_402),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_441),
.B(n_278),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_413),
.B(n_286),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_386),
.B(n_428),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_447),
.B(n_286),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_423),
.B(n_44),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_450),
.B(n_24),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_449),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_447),
.B(n_286),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_389),
.B(n_286),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_391),
.B(n_286),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_416),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_391),
.B(n_278),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_278),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_386),
.B(n_25),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_443),
.A2(n_283),
.B(n_282),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_442),
.B(n_280),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_444),
.B(n_280),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_419),
.B(n_26),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_400),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_414),
.B(n_280),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_403),
.B(n_280),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_456),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_456),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_404),
.B(n_45),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_411),
.B(n_282),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_426),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_466),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_517),
.Y(n_546)
);

NAND2x1_ASAP7_75t_SL g547 ( 
.A(n_534),
.B(n_433),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_499),
.B(n_411),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_496),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_476),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_469),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_511),
.B(n_437),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_496),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_519),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_484),
.B(n_437),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_519),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_486),
.B(n_397),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_455),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_499),
.B(n_431),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_512),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_451),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_535),
.B(n_27),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_495),
.B(n_451),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_478),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_495),
.B(n_27),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_490),
.B(n_28),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_463),
.B(n_28),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_478),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_507),
.B(n_282),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_478),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_527),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_517),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_282),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_479),
.B(n_46),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_512),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_479),
.B(n_47),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_522),
.B(n_282),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_482),
.B(n_283),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_528),
.B(n_29),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_514),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_465),
.B(n_283),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_515),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_520),
.B(n_29),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_514),
.B(n_49),
.Y(n_589)
);

NAND2x1_ASAP7_75t_L g590 ( 
.A(n_460),
.B(n_52),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_53),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_460),
.B(n_520),
.Y(n_592)
);

CKINVDCx11_ASAP7_75t_R g593 ( 
.A(n_544),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_505),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_465),
.B(n_283),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_461),
.B(n_30),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_505),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_461),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_487),
.B(n_501),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_487),
.B(n_57),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_462),
.B(n_31),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_527),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_488),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_543),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_501),
.B(n_58),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_563),
.Y(n_611)
);

INVxp67_ASAP7_75t_SL g612 ( 
.A(n_584),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_592),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_552),
.B(n_474),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_554),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

BUFx4f_ASAP7_75t_L g617 ( 
.A(n_584),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_610),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_584),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

INVx3_ASAP7_75t_SL g621 ( 
.A(n_592),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_607),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_546),
.Y(n_623)
);

INVx3_ASAP7_75t_SL g624 ( 
.A(n_592),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_610),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_568),
.A2(n_482),
.B1(n_518),
.B2(n_477),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_584),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_593),
.Y(n_630)
);

INVx5_ASAP7_75t_SL g631 ( 
.A(n_591),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_548),
.B(n_488),
.Y(n_632)
);

BUFx12f_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

BUFx4f_ASAP7_75t_SL g634 ( 
.A(n_564),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_551),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_559),
.B(n_474),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_555),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_501),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_585),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_606),
.B(n_524),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_608),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_575),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_585),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_585),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_585),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_565),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_568),
.B(n_462),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_591),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_551),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_598),
.B(n_491),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_607),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_574),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_591),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

BUFx5_ASAP7_75t_L g658 ( 
.A(n_589),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_589),
.Y(n_659)
);

BUFx12f_ASAP7_75t_L g660 ( 
.A(n_593),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_598),
.B(n_491),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_598),
.B(n_467),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_574),
.Y(n_663)
);

BUFx12f_ASAP7_75t_L g664 ( 
.A(n_558),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_567),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

BUFx4f_ASAP7_75t_SL g667 ( 
.A(n_629),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_630),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_637),
.A2(n_566),
.B1(n_563),
.B2(n_583),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_626),
.A2(n_599),
.B1(n_589),
.B2(n_566),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_643),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_614),
.A2(n_583),
.B1(n_570),
.B2(n_596),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_615),
.Y(n_673)
);

BUFx6f_ASAP7_75t_SL g674 ( 
.A(n_642),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_611),
.A2(n_582),
.B1(n_570),
.B2(n_588),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_638),
.A2(n_557),
.B1(n_558),
.B2(n_572),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_660),
.Y(n_677)
);

AO22x1_ASAP7_75t_L g678 ( 
.A1(n_621),
.A2(n_476),
.B1(n_558),
.B2(n_569),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

BUFx4f_ASAP7_75t_L g682 ( 
.A(n_660),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_620),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_633),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_616),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_632),
.A2(n_558),
.B1(n_599),
.B2(n_536),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_558),
.B1(n_604),
.B2(n_599),
.Y(n_687)
);

INVx6_ASAP7_75t_L g688 ( 
.A(n_633),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_616),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_648),
.B(n_467),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_634),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_625),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_642),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_659),
.A2(n_493),
.B1(n_516),
.B2(n_602),
.Y(n_694)
);

BUFx10_ASAP7_75t_L g695 ( 
.A(n_619),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_639),
.B(n_468),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_611),
.A2(n_541),
.B1(n_476),
.B2(n_609),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_649),
.A2(n_472),
.B(n_577),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_625),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_611),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_L g701 ( 
.A1(n_639),
.A2(n_473),
.B1(n_600),
.B2(n_515),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_618),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_618),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_L g704 ( 
.A1(n_641),
.A2(n_502),
.B(n_498),
.Y(n_704)
);

INVx6_ASAP7_75t_L g705 ( 
.A(n_620),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_664),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_635),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_659),
.A2(n_662),
.B1(n_653),
.B2(n_650),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_620),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_635),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_471),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_636),
.Y(n_712)
);

INVx6_ASAP7_75t_L g713 ( 
.A(n_623),
.Y(n_713)
);

OAI21xp33_ASAP7_75t_L g714 ( 
.A1(n_662),
.A2(n_547),
.B(n_542),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_623),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_621),
.A2(n_601),
.B1(n_539),
.B2(n_540),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_666),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_668),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_669),
.A2(n_611),
.B1(n_656),
.B2(n_613),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_671),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_705),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_690),
.B(n_613),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_712),
.Y(n_724)
);

INVx5_ASAP7_75t_SL g725 ( 
.A(n_683),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_680),
.Y(n_726)
);

OAI21xp33_ASAP7_75t_L g727 ( 
.A1(n_672),
.A2(n_470),
.B(n_483),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_675),
.A2(n_656),
.B1(n_627),
.B2(n_653),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_693),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_697),
.A2(n_650),
.B1(n_653),
.B2(n_621),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_673),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_677),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_700),
.A2(n_676),
.B1(n_687),
.B2(n_670),
.Y(n_735)
);

OAI21xp5_ASAP7_75t_L g736 ( 
.A1(n_698),
.A2(n_661),
.B(n_652),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_714),
.A2(n_627),
.B1(n_650),
.B2(n_661),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_SL g738 ( 
.A1(n_706),
.A2(n_664),
.B1(n_624),
.B2(n_601),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_704),
.A2(n_652),
.B1(n_624),
.B2(n_601),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_689),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_707),
.Y(n_741)
);

BUFx6f_ASAP7_75t_SL g742 ( 
.A(n_683),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

AOI222xp33_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_468),
.B1(n_530),
.B2(n_472),
.C1(n_631),
.C2(n_578),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_686),
.A2(n_624),
.B1(n_631),
.B2(n_617),
.Y(n_745)
);

INVx8_ASAP7_75t_L g746 ( 
.A(n_674),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_695),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_715),
.B(n_623),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_716),
.A2(n_631),
.B1(n_658),
.B2(n_577),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_SL g750 ( 
.A1(n_682),
.A2(n_631),
.B1(n_658),
.B2(n_579),
.Y(n_750)
);

NOR2x1_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_644),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_701),
.B(n_658),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_711),
.A2(n_601),
.B1(n_631),
.B2(n_483),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_682),
.A2(n_562),
.B1(n_545),
.B2(n_538),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_702),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_710),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_692),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_699),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_679),
.Y(n_759)
);

AOI222xp33_ASAP7_75t_L g760 ( 
.A1(n_667),
.A2(n_468),
.B1(n_579),
.B2(n_471),
.C1(n_489),
.C2(n_504),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_SL g761 ( 
.A1(n_688),
.A2(n_658),
.B1(n_609),
.B2(n_523),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_674),
.A2(n_658),
.B1(n_609),
.B2(n_494),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_688),
.A2(n_658),
.B1(n_494),
.B2(n_523),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_705),
.A2(n_617),
.B1(n_644),
.B2(n_539),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_713),
.A2(n_617),
.B1(n_644),
.B2(n_493),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_SL g766 ( 
.A1(n_713),
.A2(n_658),
.B1(n_628),
.B2(n_645),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_703),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_684),
.A2(n_590),
.B1(n_612),
.B2(n_646),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_683),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_709),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_709),
.A2(n_493),
.B1(n_516),
.B2(n_574),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_678),
.B(n_658),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_679),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_709),
.Y(n_774)
);

OAI222xp33_ASAP7_75t_L g775 ( 
.A1(n_694),
.A2(n_665),
.B1(n_521),
.B2(n_513),
.C1(n_581),
.C2(n_594),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_669),
.B(n_516),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_705),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_728),
.A2(n_646),
.B1(n_628),
.B2(n_645),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_722),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_735),
.A2(n_776),
.B1(n_738),
.B2(n_727),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_734),
.B(n_636),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_719),
.A2(n_658),
.B1(n_536),
.B2(n_480),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_773),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_740),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_723),
.B(n_665),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_745),
.A2(n_485),
.B1(n_481),
.B2(n_619),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_717),
.Y(n_787)
);

OAI211xp5_ASAP7_75t_L g788 ( 
.A1(n_760),
.A2(n_510),
.B(n_525),
.C(n_497),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_761),
.A2(n_628),
.B1(n_645),
.B2(n_605),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_744),
.A2(n_475),
.B1(n_480),
.B2(n_496),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_743),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_743),
.A2(n_640),
.B1(n_619),
.B2(n_647),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_R g793 ( 
.A(n_772),
.B(n_752),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_647),
.B1(n_640),
.B2(n_619),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_731),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_741),
.B(n_651),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_749),
.A2(n_640),
.B1(n_619),
.B2(n_647),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_736),
.A2(n_654),
.B(n_622),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_730),
.A2(n_628),
.B1(n_645),
.B2(n_619),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_720),
.B(n_651),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_SL g801 ( 
.A1(n_771),
.A2(n_607),
.B(n_655),
.Y(n_801)
);

AOI222xp33_ASAP7_75t_L g802 ( 
.A1(n_737),
.A2(n_497),
.B1(n_594),
.B2(n_597),
.C1(n_581),
.C2(n_500),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_749),
.A2(n_647),
.B1(n_640),
.B2(n_597),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_761),
.A2(n_739),
.B1(n_762),
.B2(n_753),
.Y(n_804)
);

OAI222xp33_ASAP7_75t_L g805 ( 
.A1(n_750),
.A2(n_586),
.B1(n_595),
.B2(n_571),
.C1(n_573),
.C2(n_561),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_774),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_SL g807 ( 
.A1(n_746),
.A2(n_628),
.B1(n_645),
.B2(n_640),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_754),
.A2(n_647),
.B1(n_640),
.B2(n_553),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_754),
.A2(n_647),
.B1(n_549),
.B2(n_553),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_750),
.A2(n_549),
.B1(n_553),
.B2(n_603),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_768),
.A2(n_492),
.B1(n_527),
.B2(n_464),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_746),
.A2(n_729),
.B1(n_777),
.B2(n_721),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_763),
.A2(n_628),
.B1(n_645),
.B2(n_574),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_748),
.A2(n_549),
.B1(n_603),
.B2(n_573),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_751),
.A2(n_603),
.B1(n_571),
.B2(n_464),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_774),
.A2(n_464),
.B1(n_622),
.B2(n_654),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_766),
.A2(n_605),
.B1(n_622),
.B2(n_654),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_769),
.A2(n_464),
.B1(n_654),
.B2(n_560),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_770),
.A2(n_464),
.B1(n_560),
.B2(n_503),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_742),
.A2(n_464),
.B1(n_503),
.B2(n_605),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_742),
.A2(n_605),
.B1(n_657),
.B2(n_655),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_755),
.A2(n_605),
.B1(n_657),
.B2(n_655),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_756),
.A2(n_663),
.B1(n_657),
.B2(n_655),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_757),
.A2(n_663),
.B1(n_657),
.B2(n_655),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_758),
.A2(n_663),
.B1(n_657),
.B2(n_655),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_767),
.A2(n_663),
.B1(n_657),
.B2(n_580),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_777),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_784),
.B(n_759),
.Y(n_828)
);

OAI221xp5_ASAP7_75t_L g829 ( 
.A1(n_780),
.A2(n_788),
.B1(n_782),
.B2(n_804),
.C(n_790),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_799),
.A2(n_765),
.B1(n_764),
.B2(n_766),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_784),
.B(n_759),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_787),
.B(n_795),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_778),
.A2(n_718),
.B1(n_724),
.B2(n_726),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_793),
.B(n_747),
.C(n_732),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_SL g835 ( 
.A1(n_812),
.A2(n_797),
.B(n_811),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_806),
.B(n_725),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_779),
.A2(n_775),
.B1(n_747),
.B2(n_531),
.C(n_533),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_794),
.B(n_733),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_793),
.B(n_733),
.C(n_526),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_785),
.B(n_725),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_803),
.A2(n_725),
.B1(n_733),
.B2(n_663),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_826),
.B(n_733),
.C(n_663),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_786),
.B(n_576),
.C(n_533),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_791),
.B(n_32),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_791),
.B(n_32),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_783),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_L g847 ( 
.A(n_823),
.B(n_532),
.C(n_775),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_796),
.B(n_33),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_SL g849 ( 
.A(n_800),
.B(n_537),
.C(n_35),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_798),
.B(n_508),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_781),
.B(n_34),
.Y(n_851)
);

AOI211xp5_ASAP7_75t_L g852 ( 
.A1(n_789),
.A2(n_34),
.B(n_35),
.C(n_59),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_781),
.B(n_60),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_796),
.B(n_61),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_783),
.B(n_62),
.Y(n_855)
);

AND2x2_ASAP7_75t_SL g856 ( 
.A(n_808),
.B(n_64),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_824),
.B(n_65),
.C(n_66),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_809),
.A2(n_508),
.B1(n_68),
.B2(n_71),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_783),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_SL g860 ( 
.A1(n_807),
.A2(n_508),
.B(n_72),
.Y(n_860)
);

NAND4xp25_ASAP7_75t_L g861 ( 
.A(n_792),
.B(n_67),
.C(n_75),
.D(n_76),
.Y(n_861)
);

OA21x2_ASAP7_75t_L g862 ( 
.A1(n_805),
.A2(n_78),
.B(n_79),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_813),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_834),
.B(n_827),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_839),
.B(n_801),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_832),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_840),
.B(n_827),
.Y(n_867)
);

OAI211xp5_ASAP7_75t_SL g868 ( 
.A1(n_849),
.A2(n_814),
.B(n_825),
.C(n_810),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_828),
.B(n_817),
.Y(n_869)
);

NAND4xp75_ASAP7_75t_L g870 ( 
.A(n_838),
.B(n_827),
.C(n_821),
.D(n_801),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_846),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_846),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_832),
.B(n_831),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_836),
.Y(n_874)
);

XOR2x2_ASAP7_75t_L g875 ( 
.A(n_829),
.B(n_86),
.Y(n_875)
);

AOI211xp5_ASAP7_75t_L g876 ( 
.A1(n_835),
.A2(n_827),
.B(n_88),
.C(n_89),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_852),
.B(n_802),
.C(n_822),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_844),
.B(n_815),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_843),
.B(n_820),
.C(n_816),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_859),
.B(n_818),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_861),
.B(n_819),
.C(n_90),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_859),
.B(n_846),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_845),
.B(n_87),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_844),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_851),
.B(n_848),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_848),
.B(n_837),
.Y(n_886)
);

AOI211xp5_ASAP7_75t_L g887 ( 
.A1(n_860),
.A2(n_857),
.B(n_842),
.C(n_841),
.Y(n_887)
);

NAND4xp75_ASAP7_75t_SL g888 ( 
.A(n_864),
.B(n_862),
.C(n_870),
.D(n_876),
.Y(n_888)
);

XNOR2xp5_ASAP7_75t_L g889 ( 
.A(n_875),
.B(n_854),
.Y(n_889)
);

OAI22xp33_ASAP7_75t_L g890 ( 
.A1(n_877),
.A2(n_862),
.B1(n_847),
.B2(n_838),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_873),
.B(n_854),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_874),
.Y(n_892)
);

XOR2xp5_ASAP7_75t_L g893 ( 
.A(n_885),
.B(n_833),
.Y(n_893)
);

XOR2x2_ASAP7_75t_L g894 ( 
.A(n_886),
.B(n_856),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_L g895 ( 
.A(n_887),
.B(n_853),
.C(n_850),
.Y(n_895)
);

NAND4xp75_ASAP7_75t_L g896 ( 
.A(n_865),
.B(n_856),
.C(n_862),
.D(n_855),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_884),
.B(n_830),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_866),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_872),
.B(n_855),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_882),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_873),
.B(n_850),
.Y(n_901)
);

NAND4xp75_ASAP7_75t_L g902 ( 
.A(n_886),
.B(n_863),
.C(n_858),
.D(n_96),
.Y(n_902)
);

INVx1_ASAP7_75t_SL g903 ( 
.A(n_883),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_872),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_897),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_904),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_900),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_899),
.B(n_867),
.Y(n_908)
);

XOR2x2_ASAP7_75t_L g909 ( 
.A(n_894),
.B(n_881),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_901),
.Y(n_910)
);

XOR2x2_ASAP7_75t_L g911 ( 
.A(n_894),
.B(n_879),
.Y(n_911)
);

XNOR2x1_ASAP7_75t_L g912 ( 
.A(n_889),
.B(n_878),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_904),
.B(n_871),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_907),
.Y(n_914)
);

OA22x2_ASAP7_75t_L g915 ( 
.A1(n_905),
.A2(n_897),
.B1(n_893),
.B2(n_892),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_910),
.B(n_891),
.Y(n_916)
);

OA22x2_ASAP7_75t_L g917 ( 
.A1(n_911),
.A2(n_903),
.B1(n_904),
.B2(n_899),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_907),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_906),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_911),
.A2(n_909),
.B1(n_890),
.B2(n_896),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_906),
.Y(n_921)
);

OAI22x1_ASAP7_75t_L g922 ( 
.A1(n_913),
.A2(n_895),
.B1(n_898),
.B2(n_888),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_922),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_914),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_920),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_919),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_921),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_924),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_926),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_925),
.Y(n_930)
);

AO22x2_ASAP7_75t_L g931 ( 
.A1(n_929),
.A2(n_923),
.B1(n_927),
.B2(n_912),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_930),
.A2(n_923),
.B1(n_917),
.B2(n_915),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_928),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_930),
.A2(n_912),
.B1(n_890),
.B2(n_916),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_931),
.B(n_918),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_932),
.A2(n_909),
.B1(n_914),
.B2(n_902),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_934),
.A2(n_913),
.B1(n_868),
.B2(n_908),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_933),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_934),
.B(n_913),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_931),
.A2(n_869),
.B1(n_880),
.B2(n_882),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_933),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_938),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_936),
.A2(n_939),
.B1(n_935),
.B2(n_937),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_941),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_940),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_936),
.A2(n_880),
.B1(n_94),
.B2(n_97),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_938),
.Y(n_947)
);

INVxp67_ASAP7_75t_SL g948 ( 
.A(n_939),
.Y(n_948)
);

OAI211xp5_ASAP7_75t_L g949 ( 
.A1(n_943),
.A2(n_93),
.B(n_98),
.C(n_102),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_942),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_948),
.A2(n_103),
.B(n_104),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_944),
.Y(n_952)
);

AND2x4_ASAP7_75t_SL g953 ( 
.A(n_947),
.B(n_945),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_946),
.A2(n_106),
.B1(n_108),
.B2(n_114),
.Y(n_954)
);

NAND4xp25_ASAP7_75t_L g955 ( 
.A(n_943),
.B(n_115),
.C(n_116),
.D(n_117),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_953),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_949),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_957)
);

OR3x2_ASAP7_75t_L g958 ( 
.A(n_955),
.B(n_122),
.C(n_124),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_950),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_952),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_953),
.Y(n_963)
);

OAI211xp5_ASAP7_75t_SL g964 ( 
.A1(n_950),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_956),
.A2(n_128),
.B1(n_131),
.B2(n_138),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_SL g966 ( 
.A1(n_963),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_962),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_960),
.Y(n_968)
);

OAI22x1_ASAP7_75t_L g969 ( 
.A1(n_959),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_961),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_958),
.A2(n_153),
.B1(n_154),
.B2(n_159),
.Y(n_971)
);

NAND4xp25_ASAP7_75t_L g972 ( 
.A(n_957),
.B(n_160),
.C(n_162),
.D(n_163),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_964),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_957),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_968),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_969),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_974),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_970),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_973),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_971),
.Y(n_980)
);

OAI22xp33_ASAP7_75t_L g981 ( 
.A1(n_975),
.A2(n_972),
.B1(n_965),
.B2(n_966),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_977),
.A2(n_967),
.B1(n_165),
.B2(n_166),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_976),
.A2(n_979),
.B1(n_980),
.B2(n_975),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_983),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_981),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_984),
.A2(n_985),
.B1(n_978),
.B2(n_982),
.Y(n_986)
);

OA22x2_ASAP7_75t_L g987 ( 
.A1(n_984),
.A2(n_164),
.B1(n_167),
.B2(n_170),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_984),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_986),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_987),
.Y(n_990)
);

AOI221xp5_ASAP7_75t_L g991 ( 
.A1(n_989),
.A2(n_988),
.B1(n_178),
.B2(n_179),
.C(n_181),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_990),
.B1(n_182),
.B2(n_183),
.Y(n_992)
);


endmodule