module fake_jpeg_31868_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_27),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_17),
.B1(n_20),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_29),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_61),
.Y(n_82)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_71),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_52),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_73),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_24),
.B(n_37),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_35),
.C(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_53),
.B(n_21),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_0),
.B(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_34),
.B1(n_43),
.B2(n_3),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_57),
.B1(n_47),
.B2(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_11),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_91),
.B(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_69),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_76),
.B1(n_68),
.B2(n_71),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_86),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_79),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_81),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_93),
.C(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_102),
.C(n_94),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_88),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_63),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_119),
.C(n_112),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_104),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_78),
.B1(n_77),
.B2(n_57),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_107),
.C(n_109),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_73),
.A3(n_67),
.B1(n_65),
.B2(n_2),
.Y(n_120)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_2),
.B(n_3),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_122),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_118),
.A3(n_106),
.B1(n_113),
.B2(n_74),
.C1(n_11),
.C2(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_4),
.C(n_49),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_4),
.B(n_49),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_123),
.C(n_126),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_127),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.C(n_130),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_4),
.Y(n_138)
);


endmodule