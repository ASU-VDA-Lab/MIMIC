module fake_ariane_2696_n_1761 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1761);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1761;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_3),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_57),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_48),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_52),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_106),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

BUFx2_ASAP7_75t_SL g181 ( 
.A(n_68),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_80),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_66),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_36),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_39),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_45),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_59),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_41),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_44),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_103),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_13),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_131),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_29),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_133),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_56),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_97),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_25),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_93),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_49),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_64),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_118),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_32),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_165),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_22),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_122),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_37),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_111),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_36),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_163),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_30),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_83),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_28),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_34),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_84),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_30),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_25),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_86),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_32),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_119),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_29),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_5),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_125),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_78),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_50),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_143),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_27),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_94),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_116),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_148),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_45),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_38),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_100),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_19),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_41),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_69),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_102),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_62),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_98),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_46),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_91),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_149),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_130),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_7),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_5),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_55),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_42),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_105),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_135),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_123),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_7),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_136),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_81),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_104),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_2),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_20),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_150),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_61),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_67),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_49),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_35),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_79),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_89),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_132),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_141),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_157),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_120),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_137),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_23),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_0),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_121),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_115),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_127),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_42),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_73),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_14),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_139),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_23),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_65),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_31),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_34),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_124),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_72),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_46),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_142),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_51),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_176),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_195),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_251),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_209),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_300),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_167),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_213),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_187),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_183),
.B(n_328),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_275),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_325),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_275),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_232),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_325),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_233),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_309),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_270),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_260),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_285),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_209),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_312),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_193),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_R g363 ( 
.A(n_201),
.B(n_58),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_275),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_209),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

BUFx6f_ASAP7_75t_SL g369 ( 
.A(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_199),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_169),
.B(n_0),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_260),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_215),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_306),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_168),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_168),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_235),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_174),
.B(n_1),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_221),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_178),
.B(n_185),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_265),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_306),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_171),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_279),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_172),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_177),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_190),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_172),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_173),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_224),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_173),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_187),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_200),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_243),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_260),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_175),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_175),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_296),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_264),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_216),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_303),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_264),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_180),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_264),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_205),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_205),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_186),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_248),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_249),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_344),
.B(n_315),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_202),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_341),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_230),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_230),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_346),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_238),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_342),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_382),
.B(n_290),
.C(n_238),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_350),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_356),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_358),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_339),
.B(n_256),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_379),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_359),
.B(n_276),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_290),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_347),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_291),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_361),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_186),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_343),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_395),
.B(n_291),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_278),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_334),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_385),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_394),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_288),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_387),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_331),
.B(n_320),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_386),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_401),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_335),
.B(n_301),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_390),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_353),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

NAND3xp33_ASAP7_75t_L g466 ( 
.A(n_371),
.B(n_322),
.C(n_320),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_336),
.B(n_338),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_404),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_407),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_391),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_391),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_409),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_393),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_373),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_360),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_362),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_366),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_370),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_374),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_466),
.A2(n_352),
.B1(n_369),
.B2(n_398),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_447),
.B(n_357),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_355),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_413),
.B(n_333),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_447),
.B(n_397),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_420),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_479),
.B(n_393),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_479),
.B(n_399),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_333),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_479),
.B(n_399),
.Y(n_500)
);

BUFx10_ASAP7_75t_L g501 ( 
.A(n_460),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_479),
.B(n_337),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_402),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_337),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_400),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_478),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_448),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVx8_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_481),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_480),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_474),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_188),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_480),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_433),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_421),
.B(n_400),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_425),
.B(n_332),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_475),
.B(n_239),
.C(n_330),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_439),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_484),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_484),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_417),
.B(n_411),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_431),
.B(n_436),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_345),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

BUFx4_ASAP7_75t_L g529 ( 
.A(n_454),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_444),
.B(n_345),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_417),
.B(n_381),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_486),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_440),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_422),
.B(n_392),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_432),
.B(n_340),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_416),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_444),
.B(n_406),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_481),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_445),
.B(n_406),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_445),
.B(n_455),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_455),
.B(n_340),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_432),
.B(n_348),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_457),
.B(n_481),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_477),
.B(n_348),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_457),
.B(n_482),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_459),
.B(n_482),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_482),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_459),
.B(n_364),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_420),
.Y(n_553)
);

AND3x2_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_405),
.C(n_372),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_422),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_482),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_423),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_364),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_458),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_428),
.Y(n_561)
);

INVx6_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_466),
.A2(n_369),
.B1(n_388),
.B2(n_322),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_426),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_425),
.B(n_396),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_485),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_419),
.B(n_188),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_376),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_376),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_419),
.B(n_225),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_419),
.A2(n_435),
.B1(n_437),
.B2(n_441),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_453),
.B(n_384),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_429),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_435),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_435),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_420),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_435),
.B(n_365),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_470),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_384),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_470),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_446),
.B(n_369),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_473),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_451),
.B(n_368),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_430),
.B(n_241),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_473),
.B(n_179),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_476),
.B(n_210),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_453),
.B(n_194),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_463),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_438),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_456),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_437),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_437),
.B(n_271),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_437),
.B(n_295),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_472),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_451),
.B(n_305),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_441),
.B(n_323),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_441),
.B(n_202),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g607 ( 
.A(n_427),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_441),
.B(n_259),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_469),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_440),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_469),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_440),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_469),
.A2(n_286),
.B1(n_299),
.B2(n_324),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_427),
.B(n_442),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_427),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_442),
.B(n_326),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_442),
.B(n_180),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_418),
.B(n_274),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_440),
.Y(n_620)
);

BUFx6f_ASAP7_75t_SL g621 ( 
.A(n_461),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_442),
.B(n_182),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_443),
.A2(n_310),
.B1(n_308),
.B2(n_282),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_443),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_443),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_443),
.B(n_182),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_468),
.A2(n_253),
.B1(n_254),
.B2(n_268),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_418),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_418),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_424),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_461),
.B(n_259),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_461),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_424),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_424),
.Y(n_635)
);

INVx8_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_495),
.A2(n_198),
.B(n_196),
.C(n_194),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_588),
.B(n_601),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_526),
.A2(n_468),
.B(n_450),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_568),
.A2(n_280),
.B1(n_198),
.B2(n_246),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_493),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_528),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_545),
.B(n_184),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_531),
.B(n_196),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_582),
.A2(n_273),
.B1(n_192),
.B2(n_327),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_508),
.B(n_184),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_568),
.A2(n_273),
.B1(n_225),
.B2(n_287),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_488),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_536),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_543),
.A2(n_468),
.B(n_450),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_287),
.B1(n_181),
.B2(n_280),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_504),
.B(n_492),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_528),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_587),
.B(n_189),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_519),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_507),
.B(n_585),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_189),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_491),
.A2(n_246),
.B1(n_282),
.B2(n_293),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_SL g662 ( 
.A(n_512),
.B(n_489),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_509),
.B(n_187),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_569),
.B(n_191),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_629),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_503),
.B(n_525),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_570),
.B(n_203),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_566),
.A2(n_311),
.B1(n_293),
.B2(n_240),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_510),
.B(n_191),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_510),
.B(n_192),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_565),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_552),
.B(n_204),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_499),
.B(n_237),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_506),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_525),
.B(n_311),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_586),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_502),
.B(n_237),
.Y(n_677)
);

NAND2x1_ASAP7_75t_L g678 ( 
.A(n_540),
.B(n_450),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_SL g679 ( 
.A1(n_516),
.A2(n_219),
.B1(n_227),
.B2(n_226),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_552),
.A2(n_245),
.B1(n_281),
.B2(n_327),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_555),
.B(n_245),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_555),
.B(n_281),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_586),
.B(n_283),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_497),
.A2(n_500),
.B1(n_498),
.B2(n_527),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_548),
.A2(n_214),
.B1(n_206),
.B2(n_229),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_490),
.B(n_231),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_566),
.B(n_283),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_525),
.B(n_574),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_511),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_566),
.B(n_284),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_530),
.B(n_517),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_576),
.B(n_284),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_517),
.B(n_244),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_540),
.B(n_289),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_519),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_598),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_540),
.B(n_289),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_537),
.B(n_250),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_576),
.B(n_292),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_505),
.A2(n_292),
.B1(n_294),
.B2(n_298),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_556),
.B(n_294),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_558),
.B(n_298),
.Y(n_702)
);

AND2x6_ASAP7_75t_SL g703 ( 
.A(n_593),
.B(n_257),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_302),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_560),
.Y(n_705)
);

O2A1O1Ixp5_ASAP7_75t_L g706 ( 
.A1(n_550),
.A2(n_304),
.B(n_307),
.C(n_302),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_556),
.B(n_304),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_537),
.B(n_261),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_514),
.B(n_307),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_541),
.B(n_263),
.Y(n_710)
);

NOR2xp67_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_207),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_560),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_509),
.B(n_187),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_522),
.B(n_266),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_541),
.B(n_269),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_610),
.B(n_187),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_619),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_505),
.A2(n_258),
.B1(n_212),
.B2(n_217),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_SL g719 ( 
.A(n_520),
.B(n_595),
.C(n_516),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_SL g721 ( 
.A(n_595),
.B(n_313),
.C(n_314),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_523),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_497),
.B(n_318),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_524),
.B(n_208),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_509),
.B(n_363),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_501),
.B(n_2),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_501),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_532),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_539),
.B(n_589),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_610),
.B(n_329),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_501),
.B(n_591),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_498),
.B(n_329),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_500),
.B(n_255),
.C(n_220),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_590),
.B(n_252),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_550),
.B(n_531),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_531),
.B(n_262),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_557),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_592),
.Y(n_738)
);

CKINVDCx11_ASAP7_75t_R g739 ( 
.A(n_557),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_596),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_629),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_580),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_580),
.B(n_6),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_603),
.Y(n_744)
);

INVx5_ASAP7_75t_L g745 ( 
.A(n_513),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_534),
.B(n_247),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_518),
.A2(n_218),
.B1(n_222),
.B2(n_223),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_534),
.B(n_272),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_580),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_572),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_534),
.B(n_6),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_544),
.B(n_8),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_547),
.B(n_329),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_581),
.B(n_277),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_609),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_594),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_584),
.B(n_267),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_594),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_571),
.A2(n_329),
.B1(n_316),
.B2(n_321),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_602),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_549),
.B(n_329),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_597),
.B(n_319),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_602),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_597),
.B(n_317),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_628),
.Y(n_765)
);

BUFx6f_ASAP7_75t_SL g766 ( 
.A(n_557),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_242),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_600),
.B(n_236),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_605),
.B(n_234),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_551),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_561),
.B(n_228),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_607),
.A2(n_461),
.B(n_76),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_544),
.A2(n_461),
.B1(n_10),
.B2(n_11),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_604),
.B(n_9),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_9),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_559),
.B(n_10),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_563),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_567),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_612),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_573),
.B(n_518),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_562),
.B(n_577),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_518),
.B(n_11),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_562),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_518),
.B(n_14),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_562),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_571),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_561),
.B(n_16),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_606),
.B(n_18),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_624),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_561),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_615),
.A2(n_85),
.B(n_158),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_606),
.B(n_24),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_496),
.B(n_24),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_496),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_575),
.B(n_26),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_571),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_608),
.B(n_564),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_577),
.B(n_33),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_628),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_496),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_538),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_529),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_729),
.A2(n_618),
.B(n_626),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_689),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_684),
.A2(n_616),
.B(n_625),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_691),
.A2(n_616),
.B(n_625),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_691),
.A2(n_538),
.B(n_553),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_643),
.A2(n_647),
.B1(n_660),
.B2(n_659),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_667),
.B(n_571),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_641),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_669),
.A2(n_538),
.B(n_553),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_665),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_650),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_674),
.B(n_575),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_669),
.A2(n_694),
.B(n_670),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_667),
.B(n_571),
.Y(n_817)
);

AOI21x1_ASAP7_75t_L g818 ( 
.A1(n_753),
.A2(n_632),
.B(n_634),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_636),
.B(n_513),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_771),
.B(n_575),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_656),
.B(n_571),
.Y(n_821)
);

OAI21x1_ASAP7_75t_L g822 ( 
.A1(n_639),
.A2(n_632),
.B(n_553),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_670),
.A2(n_578),
.B(n_583),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_722),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_728),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_735),
.B(n_487),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_642),
.B(n_608),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_752),
.A2(n_723),
.B(n_698),
.C(n_708),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_753),
.A2(n_635),
.B(n_631),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_752),
.A2(n_622),
.B(n_583),
.C(n_578),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_665),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_647),
.A2(n_578),
.B1(n_583),
.B2(n_577),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_664),
.B(n_617),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_653),
.A2(n_613),
.B1(n_614),
.B2(n_633),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_671),
.B(n_579),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_648),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_645),
.A2(n_627),
.B(n_623),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_694),
.A2(n_613),
.B(n_630),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_697),
.A2(n_613),
.B(n_620),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_732),
.A2(n_513),
.B(n_621),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_697),
.A2(n_620),
.B(n_611),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_701),
.A2(n_620),
.B(n_611),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_701),
.A2(n_620),
.B(n_611),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_646),
.B(n_723),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_651),
.A2(n_513),
.B(n_621),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_707),
.A2(n_611),
.B(n_542),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_707),
.A2(n_542),
.B(n_533),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_678),
.A2(n_542),
.B(n_533),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_738),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_665),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_693),
.B(n_513),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_SL g852 ( 
.A1(n_794),
.A2(n_513),
.B(n_621),
.C(n_47),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_747),
.B(n_542),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_665),
.Y(n_854)
);

OAI321xp33_ASAP7_75t_L g855 ( 
.A1(n_787),
.A2(n_554),
.A3(n_515),
.B1(n_533),
.B2(n_50),
.C(n_38),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_693),
.B(n_533),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_704),
.A2(n_515),
.B(n_101),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_698),
.B(n_515),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_695),
.A2(n_515),
.B(n_96),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_653),
.A2(n_95),
.B(n_164),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_695),
.A2(n_90),
.B(n_146),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_SL g863 ( 
.A1(n_794),
.A2(n_40),
.B(n_47),
.C(n_52),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_708),
.A2(n_579),
.B(n_521),
.C(n_40),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_696),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_638),
.B(n_521),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_649),
.B(n_54),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_710),
.B(n_54),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_673),
.A2(n_60),
.B(n_70),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_710),
.A2(n_75),
.B1(n_77),
.B2(n_82),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_654),
.B(n_87),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_740),
.Y(n_872)
);

AO22x1_ASAP7_75t_L g873 ( 
.A1(n_803),
.A2(n_108),
.B1(n_117),
.B2(n_126),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_720),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_744),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_715),
.B(n_128),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_666),
.B(n_688),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_677),
.A2(n_129),
.B(n_140),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_755),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_702),
.A2(n_144),
.B(n_720),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_715),
.B(n_687),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_750),
.A2(n_756),
.B(n_802),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_747),
.B(n_731),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_750),
.A2(n_756),
.B(n_801),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_690),
.B(n_672),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_686),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_742),
.B(n_749),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_672),
.B(n_652),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_795),
.A2(n_777),
.B(n_770),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_778),
.A2(n_763),
.B(n_683),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_741),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_675),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_644),
.B(n_679),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_644),
.B(n_668),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_741),
.Y(n_895)
);

AOI21x1_ASAP7_75t_L g896 ( 
.A1(n_761),
.A2(n_716),
.B(n_730),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_779),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_800),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_668),
.B(n_661),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_717),
.B(n_790),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_652),
.B(n_780),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_737),
.B(n_791),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_798),
.B(n_743),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_751),
.B(n_655),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_761),
.A2(n_776),
.B(n_760),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_787),
.A2(n_797),
.B1(n_676),
.B2(n_700),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_797),
.A2(n_713),
.B1(n_663),
.B2(n_636),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_734),
.B(n_781),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_781),
.B(n_784),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_786),
.B(n_769),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_767),
.B(n_768),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_657),
.A2(n_705),
.B(n_658),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_685),
.A2(n_637),
.B(n_640),
.C(n_785),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_727),
.B(n_685),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_712),
.A2(n_758),
.B(n_732),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_799),
.A2(n_783),
.B1(n_725),
.B2(n_662),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_754),
.A2(n_757),
.B(n_724),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_799),
.A2(n_699),
.B1(n_692),
.B2(n_680),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_726),
.B(n_773),
.C(n_788),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_706),
.A2(n_733),
.B(n_774),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_775),
.A2(n_789),
.B(n_793),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_762),
.A2(n_764),
.B(n_709),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_736),
.A2(n_748),
.B1(n_746),
.B2(n_663),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_796),
.B(n_637),
.C(n_681),
.Y(n_924)
);

NOR2xp67_ASAP7_75t_L g925 ( 
.A(n_711),
.B(n_719),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_682),
.B(n_714),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_716),
.A2(n_730),
.B(n_765),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_636),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_772),
.A2(n_741),
.B(n_782),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_759),
.A2(n_718),
.B(n_792),
.C(n_745),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_782),
.A2(n_713),
.B(n_745),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_782),
.A2(n_713),
.B(n_745),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_759),
.B(n_782),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_766),
.A2(n_721),
.B1(n_745),
.B2(n_739),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_703),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_766),
.A2(n_659),
.B(n_707),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_659),
.A2(n_669),
.B(n_670),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_659),
.A2(n_669),
.B(n_670),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_674),
.B(n_512),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_684),
.A2(n_752),
.B(n_659),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_691),
.B(n_582),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_639),
.A2(n_651),
.B(n_550),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_L g944 ( 
.A1(n_672),
.A2(n_698),
.B(n_693),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_L g945 ( 
.A(n_650),
.B(n_512),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_639),
.A2(n_651),
.B(n_550),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_691),
.B(n_582),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_639),
.A2(n_651),
.B(n_550),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_691),
.B(n_582),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_691),
.B(n_582),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_689),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_671),
.B(n_452),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_639),
.A2(n_651),
.B(n_550),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_654),
.B(n_666),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_659),
.A2(n_669),
.B(n_670),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_691),
.B(n_582),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_691),
.B(n_582),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_SL g958 ( 
.A1(n_650),
.A2(n_595),
.B1(n_516),
.B2(n_383),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_691),
.B(n_582),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_689),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_641),
.Y(n_961)
);

NAND2x1_ASAP7_75t_L g962 ( 
.A(n_653),
.B(n_641),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_665),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_685),
.A2(n_660),
.B(n_661),
.C(n_643),
.Y(n_964)
);

INVx3_ASAP7_75t_SL g965 ( 
.A(n_650),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_689),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_674),
.B(n_512),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_691),
.B(n_582),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_671),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_638),
.Y(n_973)
);

AO21x1_ASAP7_75t_L g974 ( 
.A1(n_684),
.A2(n_752),
.B(n_659),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_689),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_691),
.B(n_582),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_689),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_691),
.B(n_582),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_729),
.A2(n_684),
.B(n_550),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_654),
.B(n_666),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_689),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_689),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_SL g987 ( 
.A1(n_899),
.A2(n_894),
.B1(n_893),
.B2(n_888),
.Y(n_987)
);

INVxp67_ASAP7_75t_SL g988 ( 
.A(n_907),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_950),
.B(n_956),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_957),
.A2(n_977),
.B1(n_971),
.B2(n_982),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_959),
.A2(n_828),
.B(n_809),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_954),
.B(n_984),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

INVx3_ASAP7_75t_SL g994 ( 
.A(n_965),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_944),
.A2(n_964),
.B(n_913),
.C(n_980),
.Y(n_995)
);

AO22x1_ASAP7_75t_L g996 ( 
.A1(n_952),
.A2(n_866),
.B1(n_914),
.B2(n_935),
.Y(n_996)
);

AO31x2_ASAP7_75t_L g997 ( 
.A1(n_941),
.A2(n_974),
.A3(n_905),
.B(n_890),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_885),
.B(n_881),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_911),
.A2(n_922),
.B(n_917),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_972),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_844),
.B(n_877),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_831),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_966),
.A2(n_970),
.B(n_969),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_966),
.A2(n_970),
.B(n_969),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_976),
.A2(n_979),
.B(n_978),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_973),
.B(n_886),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_811),
.Y(n_1007)
);

AOI21x1_ASAP7_75t_L g1008 ( 
.A1(n_905),
.A2(n_829),
.B(n_896),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_979),
.A2(n_983),
.B(n_980),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_983),
.A2(n_817),
.B(n_810),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_868),
.A2(n_918),
.B(n_926),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_808),
.A2(n_939),
.B(n_937),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_871),
.A2(n_837),
.B(n_903),
.C(n_876),
.Y(n_1013)
);

AND3x2_ASAP7_75t_L g1014 ( 
.A(n_835),
.B(n_902),
.C(n_892),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_890),
.A2(n_840),
.A3(n_804),
.B(n_816),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_808),
.A2(n_955),
.B(n_816),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_889),
.A2(n_830),
.B(n_804),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_855),
.A2(n_883),
.B(n_906),
.C(n_921),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_826),
.B(n_908),
.Y(n_1019)
);

AO31x2_ASAP7_75t_L g1020 ( 
.A1(n_930),
.A2(n_880),
.A3(n_882),
.B(n_884),
.Y(n_1020)
);

AOI21x1_ASAP7_75t_L g1021 ( 
.A1(n_818),
.A2(n_806),
.B(n_929),
.Y(n_1021)
);

BUFx4_ASAP7_75t_SL g1022 ( 
.A(n_814),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_856),
.A2(n_858),
.B(n_851),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_948),
.A2(n_953),
.B(n_822),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_806),
.A2(n_882),
.B(n_884),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_836),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_889),
.A2(n_807),
.B(n_823),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_900),
.B(n_945),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_807),
.A2(n_821),
.B(n_833),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_870),
.A2(n_901),
.B(n_923),
.C(n_916),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_874),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_961),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_812),
.A2(n_823),
.B(n_910),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_880),
.A2(n_927),
.B(n_841),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_824),
.B(n_825),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_849),
.B(n_872),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_875),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_819),
.A2(n_842),
.B(n_847),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_928),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_820),
.B(n_815),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_843),
.A2(n_846),
.B(n_839),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_879),
.B(n_986),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_SL g1043 ( 
.A1(n_933),
.A2(n_904),
.B(n_909),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_L g1044 ( 
.A1(n_920),
.A2(n_853),
.B(n_878),
.C(n_869),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_812),
.A2(n_834),
.B(n_838),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_936),
.B(n_813),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_869),
.A2(n_878),
.B(n_857),
.C(n_859),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_915),
.A2(n_912),
.B(n_845),
.Y(n_1048)
);

OR2x6_ASAP7_75t_L g1049 ( 
.A(n_958),
.B(n_925),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_831),
.B(n_895),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_938),
.B(n_985),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_951),
.B(n_981),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_960),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_967),
.B(n_975),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_827),
.A2(n_912),
.B(n_897),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_887),
.B(n_867),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_848),
.A2(n_931),
.B(n_932),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_924),
.B(n_919),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_863),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_940),
.A2(n_968),
.B1(n_832),
.B2(n_864),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_862),
.A2(n_962),
.B(n_860),
.C(n_850),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_935),
.B(n_934),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_SL g1063 ( 
.A(n_813),
.B(n_963),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_813),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_850),
.A2(n_891),
.B(n_895),
.C(n_854),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_852),
.A2(n_891),
.B(n_854),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_854),
.A2(n_861),
.B(n_963),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_861),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_861),
.B(n_963),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_873),
.A2(n_946),
.B(n_943),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_905),
.A2(n_829),
.B(n_896),
.Y(n_1071)
);

NAND2x1_ASAP7_75t_L g1072 ( 
.A(n_928),
.B(n_831),
.Y(n_1072)
);

NOR3xp33_ASAP7_75t_L g1073 ( 
.A(n_944),
.B(n_828),
.C(n_491),
.Y(n_1073)
);

AOI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_888),
.A2(n_868),
.B(n_944),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_888),
.A2(n_868),
.B(n_944),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_942),
.B(n_947),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_941),
.A2(n_974),
.B(n_946),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1080)
);

AOI21x1_ASAP7_75t_L g1081 ( 
.A1(n_905),
.A2(n_829),
.B(n_896),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_944),
.B(n_942),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_942),
.B(n_947),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1084)
);

AO221x2_ASAP7_75t_L g1085 ( 
.A1(n_942),
.A2(n_685),
.B1(n_947),
.B2(n_950),
.C(n_949),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_SL g1086 ( 
.A(n_965),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_943),
.A2(n_948),
.B(n_946),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_965),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_943),
.A2(n_948),
.B(n_946),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_813),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_944),
.B(n_942),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_814),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_805),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_905),
.A2(n_829),
.B(n_896),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_973),
.B(n_601),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_898),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_972),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_965),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_898),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_943),
.A2(n_948),
.B(n_946),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_942),
.B(n_947),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_898),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_828),
.B(n_944),
.Y(n_1104)
);

OA22x2_ASAP7_75t_L g1105 ( 
.A1(n_899),
.A2(n_894),
.B1(n_958),
.B2(n_893),
.Y(n_1105)
);

AOI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_888),
.A2(n_868),
.B(n_944),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_865),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_943),
.A2(n_948),
.B(n_946),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_942),
.A2(n_949),
.B(n_947),
.Y(n_1109)
);

INVx3_ASAP7_75t_L g1110 ( 
.A(n_928),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_942),
.B(n_947),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_943),
.A2(n_948),
.B(n_946),
.Y(n_1112)
);

NAND2x1_ASAP7_75t_L g1113 ( 
.A(n_928),
.B(n_831),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_954),
.B(n_666),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_947),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1105),
.A2(n_1085),
.B1(n_987),
.B2(n_1058),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_989),
.B(n_1077),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1054),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_1090),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_990),
.B(n_1001),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_991),
.A2(n_1009),
.B(n_1005),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_1095),
.B(n_1092),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_1073),
.B(n_1104),
.C(n_995),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1082),
.A2(n_1091),
.B(n_1011),
.C(n_1058),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_L g1127 ( 
.A(n_1088),
.B(n_1064),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_1107),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_993),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1000),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1026),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1022),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1090),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1083),
.B(n_1102),
.Y(n_1134)
);

AND2x6_ASAP7_75t_L g1135 ( 
.A(n_1059),
.B(n_1064),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_992),
.B(n_1097),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1099),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_SL g1138 ( 
.A(n_1073),
.B(n_1060),
.C(n_1056),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1022),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1001),
.B(n_1075),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1086),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1090),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1105),
.A2(n_1085),
.B1(n_988),
.B2(n_1019),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_988),
.A2(n_1115),
.B1(n_1111),
.B2(n_1080),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1013),
.A2(n_1018),
.B(n_1030),
.C(n_1076),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1012),
.A2(n_1016),
.B(n_1070),
.Y(n_1146)
);

CKINVDCx8_ASAP7_75t_R g1147 ( 
.A(n_1049),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1114),
.B(n_1039),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1109),
.B(n_1079),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1084),
.B(n_1098),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1018),
.A2(n_1030),
.B(n_1074),
.C(n_1106),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1086),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1085),
.A2(n_996),
.B1(n_987),
.B2(n_998),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1006),
.B(n_993),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_1099),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1110),
.B(n_1037),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1049),
.B(n_1028),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1053),
.B(n_1093),
.Y(n_1158)
);

AND2x6_ASAP7_75t_L g1159 ( 
.A(n_1068),
.B(n_1040),
.Y(n_1159)
);

INVxp67_ASAP7_75t_SL g1160 ( 
.A(n_1035),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_1036),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_994),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_SL g1163 ( 
.A1(n_1046),
.A2(n_1017),
.B(n_1033),
.C(n_1069),
.Y(n_1163)
);

BUFx2_ASAP7_75t_R g1164 ( 
.A(n_994),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1042),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1068),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1110),
.B(n_1063),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1051),
.B(n_1052),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1002),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1078),
.A2(n_999),
.B1(n_1045),
.B2(n_1055),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1014),
.B(n_1050),
.Y(n_1171)
);

CKINVDCx6p67_ASAP7_75t_R g1172 ( 
.A(n_1046),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1014),
.B(n_1067),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1078),
.A2(n_1027),
.B1(n_1002),
.B2(n_1029),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1050),
.B(n_1072),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1010),
.A2(n_1047),
.B(n_1112),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1078),
.A2(n_1065),
.B1(n_1113),
.B2(n_1096),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1065),
.B(n_1023),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1044),
.A2(n_1047),
.B(n_1061),
.C(n_1108),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1007),
.Y(n_1180)
);

BUFx4_ASAP7_75t_SL g1181 ( 
.A(n_1043),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1031),
.A2(n_1096),
.B1(n_1100),
.B2(n_1032),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1061),
.A2(n_1101),
.B(n_1089),
.C(n_1087),
.Y(n_1184)
);

NAND2x1_ASAP7_75t_L g1185 ( 
.A(n_1066),
.B(n_1103),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1041),
.A2(n_1038),
.B(n_1024),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_997),
.B(n_1015),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1057),
.B(n_1015),
.Y(n_1188)
);

INVx5_ASAP7_75t_L g1189 ( 
.A(n_1043),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1015),
.B(n_1025),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_997),
.B(n_1020),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1008),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1048),
.A2(n_1034),
.B(n_1021),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_1071),
.B(n_1081),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1020),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1020),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_997),
.B(n_1020),
.Y(n_1197)
);

AND2x6_ASAP7_75t_L g1198 ( 
.A(n_997),
.B(n_1094),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1114),
.B(n_666),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1114),
.B(n_666),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1082),
.A2(n_947),
.B1(n_949),
.B2(n_942),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_992),
.B(n_1000),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1022),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1054),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1054),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1054),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1086),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1114),
.B(n_666),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_SL g1211 ( 
.A1(n_989),
.A2(n_828),
.B(n_947),
.C(n_942),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1082),
.A2(n_1091),
.B1(n_987),
.B2(n_914),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1054),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1054),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1114),
.B(n_1039),
.Y(n_1216)
);

NAND2x1_ASAP7_75t_L g1217 ( 
.A(n_1066),
.B(n_831),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_SL g1218 ( 
.A(n_1018),
.B(n_907),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1107),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1082),
.B(n_1091),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_993),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1086),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1090),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1114),
.B(n_1039),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1090),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1107),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1086),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1107),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1082),
.B(n_536),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1054),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1082),
.A2(n_947),
.B1(n_949),
.B2(n_942),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1085),
.A2(n_899),
.B1(n_1091),
.B2(n_1082),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1086),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1090),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1090),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1114),
.B(n_666),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1082),
.A2(n_944),
.B(n_828),
.C(n_1091),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1082),
.A2(n_944),
.B(n_828),
.C(n_1091),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1003),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_989),
.B(n_1077),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_L g1244 ( 
.A(n_1073),
.B(n_636),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_989),
.B(n_1077),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1218),
.A2(n_1234),
.B1(n_1153),
.B2(n_1209),
.Y(n_1246)
);

CKINVDCx16_ASAP7_75t_R g1247 ( 
.A(n_1141),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1139),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1187),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1213),
.A2(n_1116),
.B1(n_1218),
.B2(n_1234),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1187),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1221),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1191),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1197),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1203),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1153),
.B(n_1125),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1183),
.Y(n_1257)
);

BUFx2_ASAP7_75t_SL g1258 ( 
.A(n_1135),
.Y(n_1258)
);

BUFx2_ASAP7_75t_R g1259 ( 
.A(n_1147),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1213),
.A2(n_1230),
.B1(n_1209),
.B2(n_1126),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_1121),
.B(n_1242),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1206),
.A2(n_1238),
.B(n_1212),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1263)
);

BUFx4_ASAP7_75t_R g1264 ( 
.A(n_1228),
.Y(n_1264)
);

CKINVDCx11_ASAP7_75t_R g1265 ( 
.A(n_1137),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1126),
.A2(n_1220),
.B1(n_1232),
.B2(n_1201),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1150),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1150),
.A2(n_1170),
.B(n_1233),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1224),
.A2(n_1170),
.B(n_1174),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1128),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1129),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1190),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1235),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1130),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1190),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1152),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1195),
.Y(n_1277)
);

AOI222xp33_ASAP7_75t_L g1278 ( 
.A1(n_1220),
.A2(n_1120),
.B1(n_1232),
.B2(n_1201),
.C1(n_1138),
.C2(n_1245),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1123),
.A2(n_1144),
.B1(n_1161),
.B2(n_1160),
.Y(n_1279)
);

BUFx6f_ASAP7_75t_L g1280 ( 
.A(n_1135),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1135),
.A2(n_1157),
.B1(n_1171),
.B2(n_1144),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1132),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1143),
.B(n_1158),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1196),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1154),
.Y(n_1285)
);

AO21x2_ASAP7_75t_L g1286 ( 
.A1(n_1194),
.A2(n_1179),
.B(n_1145),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1188),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_SL g1288 ( 
.A(n_1164),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1184),
.A2(n_1123),
.B(n_1151),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1142),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1166),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1208),
.Y(n_1292)
);

AOI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1185),
.A2(n_1149),
.B(n_1177),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1178),
.A2(n_1188),
.B(n_1149),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1117),
.A2(n_1134),
.B1(n_1243),
.B2(n_1140),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1161),
.A2(n_1124),
.B1(n_1131),
.B2(n_1200),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1130),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1219),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1146),
.A2(n_1177),
.B(n_1217),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1136),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1227),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1202),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1124),
.A2(n_1165),
.B1(n_1168),
.B2(n_1231),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1118),
.B(n_1205),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1192),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1199),
.A2(n_1210),
.B1(n_1239),
.B2(n_1180),
.Y(n_1306)
);

BUFx2_ASAP7_75t_SL g1307 ( 
.A(n_1159),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1192),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1198),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1204),
.A2(n_1207),
.B1(n_1214),
.B2(n_1215),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1198),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1119),
.A2(n_1223),
.B(n_1236),
.Y(n_1312)
);

OAI21xp33_ASAP7_75t_L g1313 ( 
.A1(n_1244),
.A2(n_1211),
.B(n_1155),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1172),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1119),
.A2(n_1237),
.B(n_1236),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1189),
.Y(n_1316)
);

INVx3_ASAP7_75t_SL g1317 ( 
.A(n_1208),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1189),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1226),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1156),
.B(n_1223),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1133),
.A2(n_1182),
.B(n_1181),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1229),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1148),
.A2(n_1225),
.B1(n_1216),
.B2(n_1122),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1127),
.A2(n_1159),
.B(n_1175),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_SL g1325 ( 
.A1(n_1216),
.A2(n_1225),
.B1(n_1159),
.B2(n_1169),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1167),
.B(n_1175),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1167),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1169),
.A2(n_1162),
.B1(n_1175),
.B2(n_1222),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1222),
.Y(n_1329)
);

BUFx10_ASAP7_75t_L g1330 ( 
.A(n_1139),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1135),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1176),
.A2(n_1193),
.B(n_1186),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_1105),
.B1(n_1085),
.B2(n_899),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1187),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1187),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1218),
.A2(n_1234),
.B1(n_1153),
.B2(n_1209),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_828),
.B2(n_1125),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1187),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_1173),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1230),
.A2(n_1234),
.B1(n_828),
.B2(n_1125),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1187),
.Y(n_1341)
);

CKINVDCx6p67_ASAP7_75t_R g1342 ( 
.A(n_1141),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1187),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1218),
.A2(n_1234),
.B1(n_1153),
.B2(n_1220),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1213),
.A2(n_1105),
.B1(n_1218),
.B2(n_1085),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1213),
.A2(n_1105),
.B1(n_1085),
.B2(n_899),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1234),
.B(n_1153),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1324),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1294),
.B(n_1347),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1294),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1294),
.B(n_1347),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1280),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1344),
.A2(n_1256),
.B1(n_1337),
.B2(n_1340),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1272),
.B(n_1275),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1274),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1294),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1267),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1253),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1268),
.Y(n_1359)
);

OR2x6_ASAP7_75t_L g1360 ( 
.A(n_1258),
.B(n_1280),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1299),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1287),
.B(n_1263),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1253),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1252),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1271),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1254),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1254),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1268),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1246),
.A2(n_1336),
.B(n_1293),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1249),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1251),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1334),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1261),
.A2(n_1269),
.B(n_1262),
.Y(n_1373)
);

OAI21xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1256),
.A2(n_1278),
.B(n_1260),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1285),
.B(n_1335),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1338),
.B(n_1341),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1338),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1298),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1341),
.B(n_1343),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1343),
.B(n_1262),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1266),
.B(n_1260),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1289),
.B(n_1269),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1332),
.A2(n_1316),
.B(n_1318),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1299),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1286),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1301),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1257),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1316),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1286),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1277),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1255),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1284),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1289),
.B(n_1283),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1301),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1322),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1284),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1305),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1305),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1321),
.A2(n_1315),
.B(n_1312),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1286),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1333),
.A2(n_1346),
.B(n_1308),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1308),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1331),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1304),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1289),
.B(n_1283),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1289),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1265),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1258),
.B(n_1307),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1309),
.B(n_1311),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1247),
.B(n_1264),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1304),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1382),
.B(n_1281),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1409),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1382),
.B(n_1281),
.Y(n_1415)
);

AND2x2_ASAP7_75t_SL g1416 ( 
.A(n_1350),
.B(n_1250),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1349),
.B(n_1339),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1409),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1376),
.B(n_1279),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1351),
.B(n_1380),
.Y(n_1420)
);

INVx4_ASAP7_75t_R g1421 ( 
.A(n_1355),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1376),
.B(n_1379),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1361),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1394),
.B(n_1345),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1394),
.B(n_1320),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1406),
.B(n_1320),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1379),
.B(n_1344),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1406),
.B(n_1407),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1412),
.B(n_1302),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1357),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1387),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1350),
.Y(n_1432)
);

NAND2x1_ASAP7_75t_L g1433 ( 
.A(n_1409),
.B(n_1327),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1356),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1356),
.B(n_1315),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1362),
.B(n_1312),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1358),
.B(n_1310),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1387),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1358),
.B(n_1313),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1390),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1390),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1384),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1373),
.B(n_1290),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1374),
.B(n_1381),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1363),
.B(n_1300),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1393),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1400),
.B(n_1326),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1386),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1397),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_L g1450 ( 
.A(n_1444),
.B(n_1374),
.C(n_1353),
.Y(n_1450)
);

AOI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1444),
.A2(n_1392),
.B1(n_1405),
.B2(n_1363),
.C(n_1366),
.Y(n_1451)
);

NAND4xp25_ASAP7_75t_L g1452 ( 
.A(n_1448),
.B(n_1329),
.C(n_1291),
.D(n_1411),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1420),
.B(n_1375),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1422),
.B(n_1364),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1422),
.B(n_1364),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1448),
.B(n_1314),
.C(n_1383),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1420),
.B(n_1375),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1420),
.B(n_1395),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

OAI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1413),
.A2(n_1399),
.B(n_1398),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1419),
.B(n_1365),
.Y(n_1462)
);

OAI211xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1446),
.A2(n_1378),
.B(n_1292),
.C(n_1396),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1425),
.B(n_1355),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.B(n_1385),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1413),
.B(n_1388),
.Y(n_1466)
);

OA211x2_ASAP7_75t_L g1467 ( 
.A1(n_1433),
.A2(n_1408),
.B(n_1328),
.C(n_1323),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1439),
.B(n_1399),
.C(n_1398),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1416),
.A2(n_1424),
.B1(n_1419),
.B2(n_1415),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1416),
.A2(n_1369),
.B1(n_1402),
.B2(n_1303),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1424),
.A2(n_1314),
.B(n_1329),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1424),
.A2(n_1401),
.B(n_1389),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1416),
.A2(n_1288),
.B1(n_1409),
.B2(n_1325),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1426),
.B(n_1389),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1431),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1413),
.B(n_1388),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1426),
.B(n_1389),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1413),
.B(n_1352),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1424),
.A2(n_1401),
.B(n_1389),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1429),
.B(n_1370),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1429),
.B(n_1371),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1427),
.A2(n_1367),
.B1(n_1366),
.B2(n_1401),
.C(n_1369),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1427),
.B(n_1371),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1426),
.B(n_1445),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1439),
.B(n_1443),
.C(n_1438),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1443),
.B(n_1403),
.C(n_1367),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1415),
.A2(n_1360),
.B1(n_1402),
.B2(n_1404),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1428),
.B(n_1401),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1416),
.A2(n_1360),
.B1(n_1306),
.B2(n_1296),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1354),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1438),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1417),
.A2(n_1369),
.B1(n_1402),
.B2(n_1360),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1428),
.B(n_1372),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1436),
.B(n_1354),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1436),
.B(n_1372),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1436),
.B(n_1354),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1443),
.B(n_1403),
.C(n_1377),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1460),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1475),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1492),
.B(n_1440),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1477),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1457),
.B(n_1432),
.Y(n_1503)
);

NAND2x1_ASAP7_75t_L g1504 ( 
.A(n_1498),
.B(n_1421),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1489),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_1408),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1465),
.B(n_1432),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1489),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1481),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1492),
.B(n_1440),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1465),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1468),
.B(n_1487),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1494),
.B(n_1440),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1484),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1474),
.B(n_1432),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1482),
.B(n_1440),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1478),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1478),
.B(n_1434),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1491),
.Y(n_1522)
);

AND2x4_ASAP7_75t_SL g1523 ( 
.A(n_1495),
.B(n_1414),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1491),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1497),
.B(n_1434),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1453),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1479),
.B(n_1414),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1451),
.B(n_1483),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1485),
.B(n_1441),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1453),
.B(n_1443),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1458),
.B(n_1435),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1459),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1450),
.B(n_1291),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1458),
.B(n_1435),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1454),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1455),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1459),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1461),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1456),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1464),
.B(n_1435),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1513),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1469),
.C(n_1470),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1499),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1499),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1539),
.B(n_1446),
.Y(n_1547)
);

INVx3_ASAP7_75t_L g1548 ( 
.A(n_1527),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1500),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

NAND4xp75_ASAP7_75t_L g1551 ( 
.A(n_1528),
.B(n_1467),
.C(n_1493),
.D(n_1479),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1524),
.B(n_1466),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1538),
.B(n_1466),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1538),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1528),
.A2(n_1473),
.B1(n_1488),
.B2(n_1369),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1533),
.B(n_1408),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1500),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1541),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1541),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1476),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1501),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1539),
.B(n_1446),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1519),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1476),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1519),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1471),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1533),
.B(n_1391),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1414),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1502),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1535),
.B(n_1430),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1502),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1505),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1509),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1536),
.B(n_1430),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1509),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1531),
.B(n_1414),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1516),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1501),
.B(n_1441),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1508),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_L g1580 ( 
.A(n_1506),
.B(n_1463),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1517),
.B(n_1449),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1543),
.B(n_1515),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1544),
.A2(n_1515),
.B(n_1504),
.Y(n_1583)
);

NAND4xp25_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1503),
.C(n_1532),
.D(n_1511),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1545),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1554),
.B(n_1517),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1545),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1546),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1553),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1578),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1569),
.B(n_1510),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1510),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1570),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1574),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1571),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1571),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1526),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1551),
.A2(n_1555),
.B1(n_1480),
.B2(n_1472),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1552),
.B(n_1527),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_1534),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1556),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1580),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1561),
.B(n_1547),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1560),
.B(n_1532),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1547),
.B(n_1534),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1581),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1551),
.A2(n_1504),
.B1(n_1520),
.B2(n_1527),
.Y(n_1618)
);

OAI21xp33_ASAP7_75t_L g1619 ( 
.A1(n_1562),
.A2(n_1560),
.B(n_1559),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1562),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1578),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1548),
.B(n_1527),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1605),
.A2(n_1580),
.B1(n_1490),
.B2(n_1402),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1612),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1558),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1614),
.B(n_1585),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1586),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1610),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1615),
.B(n_1548),
.Y(n_1631)
);

NOR2x1p5_ASAP7_75t_L g1632 ( 
.A(n_1584),
.B(n_1548),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1548),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1591),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1624),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1582),
.B(n_1587),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1611),
.B(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1589),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1618),
.A2(n_1527),
.B1(n_1520),
.B2(n_1525),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1590),
.Y(n_1641)
);

CKINVDCx16_ASAP7_75t_R g1642 ( 
.A(n_1618),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1582),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1583),
.A2(n_1558),
.B1(n_1559),
.B2(n_1563),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1587),
.B(n_1577),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1592),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1568),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1593),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1620),
.B(n_1577),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1604),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1601),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1594),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1595),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1602),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1619),
.B(n_1565),
.C(n_1563),
.Y(n_1655)
);

AO21x2_ASAP7_75t_L g1656 ( 
.A1(n_1603),
.A2(n_1550),
.B(n_1542),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1565),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1606),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1623),
.B(n_1576),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1634),
.B(n_1624),
.Y(n_1661)
);

AO32x1_ASAP7_75t_L g1662 ( 
.A1(n_1640),
.A2(n_1617),
.A3(n_1613),
.B1(n_1621),
.B2(n_1600),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1651),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1654),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1642),
.A2(n_1608),
.B(n_1598),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1635),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1654),
.Y(n_1667)
);

OAI31xp33_ASAP7_75t_L g1668 ( 
.A1(n_1643),
.A2(n_1616),
.A3(n_1567),
.B(n_1598),
.Y(n_1668)
);

A2O1A1Ixp33_ASAP7_75t_L g1669 ( 
.A1(n_1625),
.A2(n_1616),
.B(n_1597),
.C(n_1609),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1650),
.Y(n_1670)
);

AO22x2_ASAP7_75t_L g1671 ( 
.A1(n_1626),
.A2(n_1596),
.B1(n_1597),
.B2(n_1542),
.Y(n_1671)
);

AO21x1_ASAP7_75t_L g1672 ( 
.A1(n_1637),
.A2(n_1609),
.B(n_1550),
.Y(n_1672)
);

NOR4xp25_ASAP7_75t_SL g1673 ( 
.A(n_1642),
.B(n_1526),
.C(n_1423),
.D(n_1442),
.Y(n_1673)
);

OAI32xp33_ASAP7_75t_L g1674 ( 
.A1(n_1644),
.A2(n_1579),
.A3(n_1572),
.B1(n_1550),
.B2(n_1542),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1572),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1628),
.B(n_1572),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1629),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1579),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1655),
.A2(n_1579),
.B(n_1576),
.Y(n_1679)
);

NAND2x1p5_ASAP7_75t_L g1680 ( 
.A(n_1635),
.B(n_1270),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1635),
.B(n_1525),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1632),
.A2(n_1348),
.B1(n_1447),
.B2(n_1410),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1629),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1636),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1671),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1684),
.B(n_1631),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1670),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1671),
.A2(n_1632),
.B1(n_1655),
.B2(n_1656),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1677),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1661),
.B(n_1638),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1673),
.B(n_1248),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1669),
.A2(n_1631),
.B1(n_1638),
.B2(n_1633),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1661),
.B(n_1633),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1676),
.B(n_1645),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1683),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1666),
.B(n_1647),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1685),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1682),
.A2(n_1647),
.B1(n_1659),
.B2(n_1627),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1674),
.A2(n_1660),
.B1(n_1639),
.B2(n_1641),
.C1(n_1658),
.C2(n_1646),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1639),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1659),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1686),
.Y(n_1704)
);

OAI222xp33_ASAP7_75t_L g1705 ( 
.A1(n_1665),
.A2(n_1645),
.B1(n_1627),
.B2(n_1658),
.C1(n_1648),
.C2(n_1660),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1672),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1664),
.B1(n_1667),
.B2(n_1668),
.C(n_1678),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1690),
.A2(n_1662),
.B(n_1675),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_SL g1709 ( 
.A(n_1701),
.B(n_1687),
.C(n_1702),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1687),
.A2(n_1656),
.B1(n_1681),
.B2(n_1663),
.Y(n_1710)
);

AOI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1705),
.A2(n_1679),
.B1(n_1662),
.B2(n_1656),
.C(n_1646),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1696),
.A2(n_1662),
.B1(n_1641),
.B2(n_1653),
.C(n_1648),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1693),
.A2(n_1657),
.B(n_1653),
.Y(n_1713)
);

OAI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1693),
.A2(n_1689),
.B1(n_1696),
.B2(n_1694),
.C(n_1688),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_SL g1715 ( 
.A(n_1703),
.B(n_1652),
.C(n_1276),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1692),
.A2(n_1652),
.B(n_1649),
.Y(n_1716)
);

OAI211xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1691),
.A2(n_1511),
.B(n_1520),
.C(n_1537),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1691),
.A2(n_1273),
.B(n_1270),
.C(n_1342),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1710),
.B(n_1273),
.Y(n_1719)
);

NOR4xp25_ASAP7_75t_L g1720 ( 
.A(n_1709),
.B(n_1699),
.C(n_1704),
.D(n_1697),
.Y(n_1720)
);

OAI211xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1711),
.A2(n_1699),
.B(n_1700),
.C(n_1695),
.Y(n_1721)
);

NOR3x1_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_1695),
.C(n_1692),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1715),
.B(n_1698),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1698),
.C(n_1703),
.Y(n_1724)
);

OA22x2_ASAP7_75t_L g1725 ( 
.A1(n_1718),
.A2(n_1503),
.B1(n_1525),
.B2(n_1518),
.Y(n_1725)
);

AOI211xp5_ASAP7_75t_L g1726 ( 
.A1(n_1708),
.A2(n_1317),
.B(n_1255),
.C(n_1342),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1713),
.B(n_1534),
.Y(n_1727)
);

AOI211x1_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1503),
.B(n_1507),
.C(n_1518),
.Y(n_1728)
);

NOR2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1707),
.B(n_1330),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1724),
.B(n_1717),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1720),
.B(n_1247),
.C(n_1290),
.Y(n_1731)
);

OAI211xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1726),
.A2(n_1511),
.B(n_1330),
.C(n_1537),
.Y(n_1732)
);

NAND3xp33_ASAP7_75t_SL g1733 ( 
.A(n_1719),
.B(n_1330),
.C(n_1259),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1721),
.B(n_1525),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1722),
.B(n_1518),
.C(n_1507),
.D(n_1521),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1730),
.A2(n_1723),
.B1(n_1729),
.B2(n_1727),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1731),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1735),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1734),
.Y(n_1739)
);

AOI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1733),
.A2(n_1725),
.B1(n_1728),
.B2(n_1282),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1732),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1739),
.B(n_1282),
.Y(n_1742)
);

NAND4xp75_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1282),
.C(n_1530),
.D(n_1317),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1737),
.B(n_1530),
.Y(n_1744)
);

OR5x1_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1317),
.C(n_1421),
.D(n_1530),
.E(n_1525),
.Y(n_1745)
);

NAND2x1p5_ASAP7_75t_L g1746 ( 
.A(n_1741),
.B(n_1421),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1745),
.Y(n_1747)
);

NOR3xp33_ASAP7_75t_L g1748 ( 
.A(n_1742),
.B(n_1740),
.C(n_1437),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1744),
.B(n_1743),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1747),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1749),
.B2(n_1746),
.Y(n_1751)
);

OAI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1751),
.A2(n_1522),
.B1(n_1514),
.B2(n_1512),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1751),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1753),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1752),
.A2(n_1522),
.B1(n_1514),
.B2(n_1512),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1754),
.A2(n_1529),
.B(n_1516),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1755),
.Y(n_1757)
);

AOI21xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1757),
.A2(n_1756),
.B(n_1529),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1758),
.A2(n_1540),
.B1(n_1368),
.B2(n_1359),
.Y(n_1759)
);

OAI221xp5_ASAP7_75t_R g1760 ( 
.A1(n_1759),
.A2(n_1418),
.B1(n_1540),
.B2(n_1507),
.C(n_1521),
.Y(n_1760)
);

AOI211xp5_ASAP7_75t_L g1761 ( 
.A1(n_1760),
.A2(n_1540),
.B(n_1521),
.C(n_1319),
.Y(n_1761)
);


endmodule