module fake_jpeg_25957_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g72 ( 
.A(n_66),
.B(n_68),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_62),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_80),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_42),
.B1(n_61),
.B2(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_83),
.B1(n_58),
.B2(n_82),
.Y(n_98)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_47),
.B1(n_43),
.B2(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_96),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_57),
.B1(n_56),
.B2(n_58),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_100),
.B1(n_77),
.B2(n_44),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_101),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_79),
.B(n_55),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_57),
.B1(n_44),
.B2(n_53),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_93),
.B1(n_89),
.B2(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_106),
.B1(n_93),
.B2(n_90),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_55),
.B1(n_48),
.B2(n_3),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_50),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_99),
.C(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_1),
.Y(n_116)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_113),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_9),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_28),
.Y(n_133)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_88),
.B1(n_24),
.B2(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_22),
.B1(n_41),
.B2(n_37),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_127),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_107),
.C(n_51),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_29),
.C(n_12),
.Y(n_137)
);

NAND2x1_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_1),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_130),
.B(n_133),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_128),
.B1(n_11),
.B2(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_7),
.CON(n_130),
.SN(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_8),
.B(n_9),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_124),
.Y(n_139)
);

XOR2x1_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_139),
.Y(n_146)
);

OAI22x1_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_134),
.B1(n_130),
.B2(n_131),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_31),
.B(n_14),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_34),
.B1(n_20),
.B2(n_21),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_146),
.C(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_35),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_136),
.C(n_141),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_144),
.B(n_138),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_121),
.Y(n_157)
);


endmodule