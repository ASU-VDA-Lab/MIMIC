module fake_netlist_6_1999_n_5271 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_5271);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_5271;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_677;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_5239;
wire n_1971;
wire n_1781;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_2625;
wire n_1400;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_687;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_1932;
wire n_925;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_2767;
wire n_963;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_648;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_663;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_664;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4996;
wire n_4990;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_662;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_695;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_3288;
wire n_2918;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_3552;
wire n_941;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_633;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_3017;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_666;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_3294;
wire n_2457;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_4004;
wire n_2206;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_637;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_3133;
wire n_1959;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_4386;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_2803;
wire n_856;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_936;
wire n_885;
wire n_2970;
wire n_2342;
wire n_2167;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_671;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_676;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_635;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_665;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_632;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_681;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_638;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_689;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_690;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_678;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_656;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_3580;
wire n_2842;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_684;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3540;
wire n_3577;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_4533;
wire n_2218;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_651;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_2289;
wire n_1390;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_2328;
wire n_1439;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_2376;
wire n_1405;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_654;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_652;
wire n_4604;
wire n_3305;
wire n_1906;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_655;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_680;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_679;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_649;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_645;
wire n_3910;
wire n_3812;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_674;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_673;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_657;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_3103;
wire n_2354;
wire n_1475;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_642;
wire n_1159;
wire n_3481;
wire n_995;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2720;
wire n_2204;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_667;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_672;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_636;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2944;
wire n_2348;
wire n_3831;
wire n_869;
wire n_1154;
wire n_646;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_1476;
wire n_841;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_661;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2969;
wire n_2787;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_669;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_647;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_608),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_305),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_536),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_333),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_404),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_432),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_55),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_395),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_566),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_527),
.Y(n_641)
);

CKINVDCx16_ASAP7_75t_R g642 ( 
.A(n_424),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_269),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_174),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_270),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_423),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_337),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_422),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_395),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_582),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_410),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_299),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_511),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_480),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_125),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_163),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_433),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_275),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_359),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_281),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_470),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_205),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_131),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_591),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_555),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_50),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_210),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_558),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_255),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_260),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_517),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_324),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_131),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_286),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_505),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_448),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_436),
.Y(n_678)
);

CKINVDCx14_ASAP7_75t_R g679 ( 
.A(n_82),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_385),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_409),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_285),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_461),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_81),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_165),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_381),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_32),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_429),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_100),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_25),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_473),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_584),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_61),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_46),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_137),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_458),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_119),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_587),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_327),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_304),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_490),
.Y(n_701)
);

BUFx2_ASAP7_75t_SL g702 ( 
.A(n_437),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_578),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_615),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_99),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_178),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_246),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_15),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_385),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_626),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_332),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_242),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_24),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_631),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_74),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_123),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_223),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_130),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_427),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_493),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_499),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_66),
.Y(n_722)
);

CKINVDCx16_ASAP7_75t_R g723 ( 
.A(n_503),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_129),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_287),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_90),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_502),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_488),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_194),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_386),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_106),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_114),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_292),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_476),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_382),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_187),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_110),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_172),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_286),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_249),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_583),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_224),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_325),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_353),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_210),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_283),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_623),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_148),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_314),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_317),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_405),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_168),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_567),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_360),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_58),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_415),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_127),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_255),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_598),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_230),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_263),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_241),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_369),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_2),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_256),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_425),
.Y(n_766)
);

BUFx10_ASAP7_75t_L g767 ( 
.A(n_306),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_542),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_54),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_29),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_330),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_481),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_391),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_171),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_494),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_384),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_526),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_375),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_520),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_78),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_452),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_388),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_97),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_121),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_604),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_22),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_48),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_130),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_149),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_98),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_496),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_313),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_467),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_364),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_218),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_196),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_215),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_35),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_108),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_372),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_357),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_125),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_325),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_28),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_152),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_20),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_33),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_320),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_202),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_309),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_576),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_371),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_519),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_355),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_334),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_533),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_457),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_553),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_462),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_245),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_169),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_465),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_15),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_181),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_611),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_321),
.Y(n_826)
);

BUFx10_ASAP7_75t_L g827 ( 
.A(n_363),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_358),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_209),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_30),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_42),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_384),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_224),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_381),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_504),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_127),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_351),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_419),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_186),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_630),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_53),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_0),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_112),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_284),
.Y(n_844)
);

BUFx5_ASAP7_75t_L g845 ( 
.A(n_418),
.Y(n_845)
);

BUFx10_ASAP7_75t_L g846 ( 
.A(n_344),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_162),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_144),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_492),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_407),
.Y(n_850)
);

CKINVDCx14_ASAP7_75t_R g851 ( 
.A(n_170),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_551),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_299),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_359),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_162),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_205),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_194),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_148),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_112),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_388),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_108),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_257),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_219),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_53),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_48),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_78),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_197),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_609),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_329),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_145),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_350),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_579),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_217),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_329),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_28),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_77),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_279),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_58),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_244),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_40),
.Y(n_880)
);

BUFx10_ASAP7_75t_L g881 ( 
.A(n_606),
.Y(n_881)
);

CKINVDCx14_ASAP7_75t_R g882 ( 
.A(n_110),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_173),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_239),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_524),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_310),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_613),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_314),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_192),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_459),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_486),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_522),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_155),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_192),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_295),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_122),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_400),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_500),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_556),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_589),
.Y(n_900)
);

BUFx5_ASAP7_75t_L g901 ( 
.A(n_137),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_302),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_68),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_100),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_94),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_464),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_240),
.Y(n_907)
);

CKINVDCx14_ASAP7_75t_R g908 ( 
.A(n_273),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_568),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_81),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_506),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_92),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_335),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_170),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_625),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_408),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_102),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_549),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_317),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_569),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_54),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_344),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_89),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_320),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_563),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_232),
.Y(n_926)
);

BUFx8_ASAP7_75t_SL g927 ( 
.A(n_483),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_107),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_368),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_270),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_91),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_9),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_354),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_61),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_440),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_466),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_541),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_588),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_89),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_1),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_72),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_426),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_24),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_540),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_509),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_207),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_275),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_279),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_571),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_18),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_82),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_472),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_93),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_32),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_269),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_333),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_83),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_228),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_246),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_223),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_447),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_248),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_198),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_624),
.Y(n_964)
);

CKINVDCx14_ASAP7_75t_R g965 ( 
.A(n_165),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_471),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_191),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_147),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_627),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_321),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_60),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_227),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_605),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_332),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_114),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_38),
.Y(n_976)
);

BUFx2_ASAP7_75t_SL g977 ( 
.A(n_368),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_200),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_298),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_63),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_64),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_382),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_217),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_38),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_30),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_365),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_361),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_34),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_195),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_49),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_363),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_99),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_590),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_6),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_510),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_273),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_287),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_442),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_101),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_106),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_113),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_12),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_96),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_200),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_18),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_123),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_603),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_62),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_134),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_167),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_102),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_122),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_20),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_441),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_319),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_113),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_280),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_104),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_539),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_573),
.Y(n_1020)
);

BUFx10_ASAP7_75t_L g1021 ( 
.A(n_80),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_43),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_63),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_565),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_180),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_450),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_547),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_398),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_172),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_242),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_59),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_431),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_47),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_55),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_610),
.Y(n_1035)
);

BUFx10_ASAP7_75t_L g1036 ( 
.A(n_283),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_319),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_202),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_64),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_50),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_544),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_141),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_324),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_399),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_182),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_252),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_575),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_301),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_143),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_134),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_8),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_322),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_365),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_72),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_453),
.Y(n_1055)
);

BUFx5_ASAP7_75t_L g1056 ( 
.A(n_618),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_374),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_445),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_180),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_248),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_378),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_187),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_150),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_396),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_586),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_186),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_139),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_237),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_175),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_208),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_400),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_430),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_340),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_243),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_44),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_516),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_617),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_361),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_525),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_59),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_628),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_87),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_159),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_290),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_434),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_399),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_16),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_135),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_451),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_296),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_278),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_338),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_237),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_455),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_284),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_175),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_5),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_228),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_73),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_901),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_766),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_679),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_901),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1060),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_766),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_901),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_901),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_901),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_901),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_901),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_639),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_712),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_901),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_901),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_634),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_634),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_636),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_649),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_636),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1069),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1060),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_743),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_666),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_666),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_688),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_688),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_696),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_696),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_706),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_771),
.Y(n_1130)
);

INVxp33_ASAP7_75t_SL g1131 ( 
.A(n_958),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_714),
.Y(n_1132)
);

INVxp33_ASAP7_75t_SL g1133 ( 
.A(n_977),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_851),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_714),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_727),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_738),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_727),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_747),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_747),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_882),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_750),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_756),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_712),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_977),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_756),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_908),
.B(n_0),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_772),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_772),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_717),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_777),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1069),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_745),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_777),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_785),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_785),
.Y(n_1156)
);

INVxp33_ASAP7_75t_SL g1157 ( 
.A(n_633),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_710),
.Y(n_1158)
);

INVxp67_ASAP7_75t_L g1159 ( 
.A(n_638),
.Y(n_1159)
);

INVxp33_ASAP7_75t_SL g1160 ( 
.A(n_635),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_791),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_791),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1069),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_965),
.Y(n_1164)
);

CKINVDCx14_ASAP7_75t_R g1165 ( 
.A(n_881),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_811),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_811),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_717),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_790),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_818),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_818),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_835),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_835),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_840),
.Y(n_1174)
);

CKINVDCx16_ASAP7_75t_R g1175 ( 
.A(n_939),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_826),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_840),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_939),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_850),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_850),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_852),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_852),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_950),
.Y(n_1183)
);

INVxp33_ASAP7_75t_L g1184 ( 
.A(n_638),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_872),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_790),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_790),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_950),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_872),
.Y(n_1189)
);

INVxp67_ASAP7_75t_SL g1190 ( 
.A(n_650),
.Y(n_1190)
);

INVxp33_ASAP7_75t_SL g1191 ( 
.A(n_643),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_828),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_906),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_650),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_906),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_937),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_937),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_966),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_966),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_644),
.Y(n_1200)
);

CKINVDCx14_ASAP7_75t_R g1201 ( 
.A(n_881),
.Y(n_1201)
);

INVxp33_ASAP7_75t_SL g1202 ( 
.A(n_652),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1026),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1026),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_790),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_659),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_655),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1035),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1035),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1055),
.Y(n_1210)
);

CKINVDCx16_ASAP7_75t_R g1211 ( 
.A(n_642),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1055),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1058),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_790),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_874),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1073),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1058),
.Y(n_1217)
);

INVxp67_ASAP7_75t_SL g1218 ( 
.A(n_655),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_661),
.Y(n_1219)
);

INVxp33_ASAP7_75t_L g1220 ( 
.A(n_645),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1076),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1076),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1089),
.Y(n_1223)
);

INVxp33_ASAP7_75t_SL g1224 ( 
.A(n_664),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1089),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_710),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1073),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_814),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_814),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_721),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_721),
.Y(n_1231)
);

INVxp33_ASAP7_75t_L g1232 ( 
.A(n_645),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_855),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_855),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_857),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1073),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_857),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_858),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_858),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_873),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_873),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_929),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_929),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1085),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_888),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1018),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_953),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1018),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1085),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_955),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_667),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_647),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1029),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1029),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1063),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1063),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1092),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_960),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1096),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_996),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1073),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1073),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_881),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_647),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_656),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_656),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1009),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_663),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_670),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_845),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_663),
.Y(n_1273)
);

INVxp67_ASAP7_75t_L g1274 ( 
.A(n_668),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1025),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_668),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_675),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_671),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_675),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_687),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_687),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_673),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_674),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_822),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_693),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_693),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_700),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_700),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_705),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_705),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_720),
.B(n_1),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_822),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_715),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_822),
.B(n_403),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_682),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_715),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_725),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_710),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_684),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_725),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_845),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_726),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_726),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_736),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_736),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_744),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_744),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_658),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1028),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_710),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_881),
.Y(n_1311)
);

INVxp33_ASAP7_75t_SL g1312 ( 
.A(n_685),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_760),
.Y(n_1313)
);

INVxp33_ASAP7_75t_SL g1314 ( 
.A(n_686),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_891),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_760),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_765),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_690),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_703),
.Y(n_1319)
);

INVxp33_ASAP7_75t_SL g1320 ( 
.A(n_694),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1042),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_765),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_695),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_769),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_769),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_845),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_845),
.Y(n_1327)
);

BUFx2_ASAP7_75t_SL g1328 ( 
.A(n_637),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_780),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_780),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_797),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_797),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_708),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_720),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_642),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_809),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_891),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_723),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1067),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_809),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_831),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_831),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_709),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_837),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_837),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_723),
.Y(n_1346)
);

INVxp33_ASAP7_75t_L g1347 ( 
.A(n_844),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_844),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_848),
.Y(n_1349)
);

INVxp33_ASAP7_75t_SL g1350 ( 
.A(n_713),
.Y(n_1350)
);

INVxp33_ASAP7_75t_SL g1351 ( 
.A(n_716),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_718),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_848),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_859),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_859),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_722),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_864),
.Y(n_1357)
);

INVxp33_ASAP7_75t_L g1358 ( 
.A(n_864),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_720),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_720),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_865),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_865),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_870),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_710),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_870),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_871),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_703),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_724),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_651),
.B(n_2),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_871),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_876),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_876),
.Y(n_1372)
);

INVxp33_ASAP7_75t_SL g1373 ( 
.A(n_729),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_879),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_879),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_883),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_730),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_734),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_883),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_891),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_896),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_731),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_896),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_914),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_733),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_735),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_845),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_914),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_917),
.Y(n_1389)
);

INVx4_ASAP7_75t_R g1390 ( 
.A(n_651),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_917),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_931),
.Y(n_1392)
);

CKINVDCx14_ASAP7_75t_R g1393 ( 
.A(n_891),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_931),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_932),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_932),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_951),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_737),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_951),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_956),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_956),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_957),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_734),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_957),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_962),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_962),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_971),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_971),
.Y(n_1408)
);

INVxp33_ASAP7_75t_SL g1409 ( 
.A(n_739),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_892),
.Y(n_1410)
);

CKINVDCx16_ASAP7_75t_R g1411 ( 
.A(n_745),
.Y(n_1411)
);

CKINVDCx14_ASAP7_75t_R g1412 ( 
.A(n_632),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_972),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_972),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_892),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_978),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_745),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_978),
.Y(n_1418)
);

INVxp33_ASAP7_75t_L g1419 ( 
.A(n_981),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_981),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_984),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_740),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_742),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_746),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_984),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_719),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_989),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_748),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_749),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_989),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_997),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_898),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_997),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_752),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_845),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_898),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_973),
.B(n_3),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1000),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1000),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_657),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_973),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1001),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_754),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1001),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_845),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1002),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1002),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1006),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_755),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1006),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1008),
.Y(n_1451)
);

CKINVDCx16_ASAP7_75t_R g1452 ( 
.A(n_745),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1008),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_757),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1011),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_758),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1011),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1016),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1016),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_1007),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1031),
.B(n_3),
.Y(n_1461)
);

BUFx10_ASAP7_75t_L g1462 ( 
.A(n_689),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1031),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1033),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_761),
.Y(n_1465)
);

BUFx2_ASAP7_75t_SL g1466 ( 
.A(n_653),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_764),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1033),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1034),
.Y(n_1469)
);

INVxp33_ASAP7_75t_L g1470 ( 
.A(n_1034),
.Y(n_1470)
);

CKINVDCx14_ASAP7_75t_R g1471 ( 
.A(n_640),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1007),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1037),
.Y(n_1473)
);

INVxp67_ASAP7_75t_SL g1474 ( 
.A(n_812),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1037),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_770),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_845),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_773),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1061),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1061),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1066),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_762),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1066),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_774),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_719),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1071),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1071),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1043),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1074),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1074),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1082),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1082),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_776),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1090),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1090),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1099),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_778),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1099),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_660),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_782),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_660),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_641),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_845),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_961),
.B(n_4),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_699),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_699),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_803),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_803),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1158),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1485),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1169),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1169),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1263),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1264),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1485),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1102),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1108),
.A2(n_1023),
.B(n_1003),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

AOI22x1_ASAP7_75t_SL g1519 ( 
.A1(n_1111),
.A2(n_784),
.B1(n_786),
.B2(n_783),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1120),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1186),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1152),
.Y(n_1522)
);

CKINVDCx14_ASAP7_75t_R g1523 ( 
.A(n_1165),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1440),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

AND2x6_ASAP7_75t_L g1526 ( 
.A(n_1294),
.B(n_719),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1158),
.Y(n_1527)
);

INVx5_ASAP7_75t_L g1528 ( 
.A(n_1158),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1190),
.B(n_1218),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1152),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1186),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1163),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1187),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1108),
.A2(n_1023),
.B(n_1003),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1163),
.Y(n_1535)
);

AOI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1131),
.A2(n_698),
.B1(n_781),
.B2(n_753),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1462),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1168),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1158),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1187),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1158),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1112),
.A2(n_707),
.B1(n_732),
.B2(n_680),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_SL g1543 ( 
.A(n_1211),
.B(n_927),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1168),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1100),
.A2(n_1106),
.B(n_1103),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1230),
.B(n_1081),
.Y(n_1546)
);

AND2x6_ASAP7_75t_L g1547 ( 
.A(n_1294),
.B(n_719),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1205),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1226),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1178),
.Y(n_1550)
);

BUFx8_ASAP7_75t_L g1551 ( 
.A(n_1294),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1107),
.A2(n_1110),
.B(n_1109),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1102),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1226),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1134),
.Y(n_1555)
);

XNOR2xp5_ASAP7_75t_L g1556 ( 
.A(n_1111),
.B(n_801),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1226),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1284),
.B(n_719),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1205),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1226),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1328),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1226),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1298),
.Y(n_1563)
);

OAI22x1_ASAP7_75t_SL g1564 ( 
.A1(n_1118),
.A2(n_1086),
.B1(n_1087),
.B2(n_1084),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1298),
.Y(n_1565)
);

CKINVDCx6p67_ASAP7_75t_R g1566 ( 
.A(n_1335),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1298),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1214),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1298),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1178),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1113),
.A2(n_1068),
.B(n_1044),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1194),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1214),
.Y(n_1573)
);

BUFx8_ASAP7_75t_L g1574 ( 
.A(n_1153),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1216),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1188),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1216),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1292),
.B(n_1065),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1227),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1227),
.Y(n_1580)
);

INVx5_ASAP7_75t_L g1581 ( 
.A(n_1298),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1194),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1236),
.Y(n_1583)
);

BUFx12f_ASAP7_75t_L g1584 ( 
.A(n_1134),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1334),
.B(n_1065),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1310),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1150),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1310),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1249),
.B(n_689),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1310),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1188),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1207),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1310),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1236),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_L g1595 ( 
.A(n_1310),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1207),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1364),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1231),
.B(n_697),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1114),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1364),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1231),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1141),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1244),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1131),
.A2(n_1346),
.B1(n_1338),
.B2(n_1147),
.Y(n_1604)
);

INVx5_ASAP7_75t_L g1605 ( 
.A(n_1364),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1364),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1359),
.B(n_1065),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1115),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1364),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1206),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1116),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1426),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1426),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1117),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1119),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1123),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1272),
.A2(n_1068),
.B(n_1044),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1426),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1426),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1426),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1403),
.Y(n_1621)
);

INVx4_ASAP7_75t_L g1622 ( 
.A(n_1319),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1360),
.B(n_1065),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1124),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1125),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1502),
.B(n_1094),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1272),
.A2(n_702),
.B(n_1056),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1206),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1403),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1319),
.Y(n_1630)
);

BUFx12f_ASAP7_75t_L g1631 ( 
.A(n_1141),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1319),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_1466),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1164),
.Y(n_1634)
);

AND2x6_ASAP7_75t_L g1635 ( 
.A(n_1301),
.B(n_1065),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1164),
.Y(n_1636)
);

INVx5_ASAP7_75t_L g1637 ( 
.A(n_1301),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1326),
.Y(n_1638)
);

BUFx12f_ASAP7_75t_L g1639 ( 
.A(n_1271),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1326),
.A2(n_702),
.B(n_1056),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1126),
.Y(n_1641)
);

BUFx8_ASAP7_75t_SL g1642 ( 
.A(n_1118),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1502),
.B(n_646),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1327),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1271),
.Y(n_1645)
);

INVx5_ASAP7_75t_L g1646 ( 
.A(n_1327),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1278),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1387),
.Y(n_1648)
);

OAI22x1_ASAP7_75t_R g1649 ( 
.A1(n_1129),
.A2(n_800),
.B1(n_824),
.B2(n_789),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1278),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1127),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1435),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1282),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1244),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_L g1655 ( 
.A(n_1415),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1462),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1282),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1367),
.B(n_1019),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1412),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1283),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1128),
.A2(n_1135),
.B(n_1132),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1136),
.A2(n_711),
.B(n_697),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1283),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1435),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1138),
.Y(n_1665)
);

BUFx8_ASAP7_75t_SL g1666 ( 
.A(n_1129),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1445),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1228),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1139),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1477),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1415),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1432),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1308),
.B(n_1077),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1412),
.B(n_1079),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1229),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1137),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1477),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1140),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1471),
.B(n_1265),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1503),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1144),
.A2(n_1183),
.B1(n_1175),
.B2(n_1105),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1462),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1471),
.B(n_648),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1295),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1143),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1146),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1378),
.B(n_711),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1432),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1148),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1436),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1503),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1200),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1295),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1436),
.Y(n_1694)
);

BUFx6f_ASAP7_75t_L g1695 ( 
.A(n_1266),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1149),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1151),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1101),
.A2(n_825),
.B1(n_944),
.B2(n_813),
.Y(n_1698)
);

BUFx12f_ASAP7_75t_L g1699 ( 
.A(n_1318),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1499),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1121),
.A2(n_787),
.B1(n_794),
.B2(n_788),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1265),
.B(n_654),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1410),
.B(n_763),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1154),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1267),
.Y(n_1705)
);

AOI22x1_ASAP7_75t_SL g1706 ( 
.A1(n_1137),
.A2(n_796),
.B1(n_798),
.B2(n_795),
.Y(n_1706)
);

INVx4_ASAP7_75t_L g1707 ( 
.A(n_1461),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1268),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1318),
.Y(n_1709)
);

BUFx8_ASAP7_75t_SL g1710 ( 
.A(n_1176),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1270),
.Y(n_1711)
);

BUFx12f_ASAP7_75t_L g1712 ( 
.A(n_1323),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1155),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1273),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1156),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1276),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1411),
.A2(n_1014),
.B1(n_952),
.B2(n_799),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1461),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1323),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1161),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1162),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1452),
.A2(n_1482),
.B1(n_1504),
.B2(n_1157),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1166),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1167),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1170),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1171),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1157),
.B(n_662),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1172),
.A2(n_889),
.B(n_763),
.Y(n_1728)
);

INVx4_ASAP7_75t_L g1729 ( 
.A(n_1311),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1160),
.B(n_665),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1173),
.A2(n_954),
.B(n_889),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1343),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1441),
.B(n_954),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1277),
.Y(n_1734)
);

INVx5_ASAP7_75t_L g1735 ( 
.A(n_1311),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1174),
.Y(n_1736)
);

BUFx6f_ASAP7_75t_L g1737 ( 
.A(n_1279),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1501),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1343),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1177),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1233),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1160),
.B(n_669),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_L g1743 ( 
.A(n_1281),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1191),
.B(n_672),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1219),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1179),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1505),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1285),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1506),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1286),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1315),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1180),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1181),
.A2(n_1056),
.B(n_677),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1287),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1356),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1182),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1356),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1185),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1189),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1193),
.Y(n_1760)
);

INVx5_ASAP7_75t_L g1761 ( 
.A(n_1315),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1337),
.B(n_676),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1191),
.B(n_678),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1337),
.B(n_681),
.Y(n_1764)
);

BUFx3_ASAP7_75t_L g1765 ( 
.A(n_1235),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1195),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1380),
.B(n_1072),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1251),
.Y(n_1768)
);

AOI22x1_ASAP7_75t_SL g1769 ( 
.A1(n_1176),
.A2(n_804),
.B1(n_805),
.B2(n_802),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1196),
.Y(n_1770)
);

INVx5_ASAP7_75t_L g1771 ( 
.A(n_1380),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1237),
.B(n_990),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1238),
.B(n_990),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1197),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_R g1775 ( 
.A(n_1133),
.B(n_806),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1198),
.Y(n_1776)
);

INVx5_ASAP7_75t_L g1777 ( 
.A(n_1234),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1474),
.B(n_1488),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1199),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1460),
.B(n_1472),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1203),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1202),
.A2(n_808),
.B1(n_810),
.B2(n_807),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1204),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1208),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1368),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1289),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1290),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1239),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1293),
.Y(n_1789)
);

BUFx6f_ASAP7_75t_L g1790 ( 
.A(n_1297),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1240),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1507),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1291),
.B(n_1004),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1209),
.A2(n_1048),
.B(n_1004),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1210),
.B(n_834),
.Y(n_1795)
);

INVx5_ASAP7_75t_L g1796 ( 
.A(n_1153),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1508),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1300),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1212),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1302),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1213),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1299),
.Y(n_1802)
);

BUFx12f_ASAP7_75t_L g1803 ( 
.A(n_1368),
.Y(n_1803)
);

BUFx8_ASAP7_75t_SL g1804 ( 
.A(n_1192),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1165),
.B(n_683),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1417),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1217),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1377),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1221),
.A2(n_1056),
.B(n_692),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_R g1810 ( 
.A(n_1201),
.B(n_691),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1303),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1222),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1377),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1333),
.Y(n_1814)
);

INVxp67_ASAP7_75t_L g1815 ( 
.A(n_1497),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1201),
.B(n_701),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1223),
.Y(n_1817)
);

AND2x6_ASAP7_75t_L g1818 ( 
.A(n_1369),
.B(n_893),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1225),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1304),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1305),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1202),
.A2(n_820),
.B1(n_821),
.B2(n_815),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1241),
.B(n_1048),
.Y(n_1823)
);

OA21x2_ASAP7_75t_L g1824 ( 
.A1(n_1437),
.A2(n_1054),
.B(n_829),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1393),
.B(n_704),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1385),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1306),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1242),
.Y(n_1828)
);

AND2x2_ASAP7_75t_SL g1829 ( 
.A(n_1382),
.B(n_762),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1307),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1313),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1316),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1385),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1317),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1322),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1398),
.Y(n_1836)
);

BUFx8_ASAP7_75t_SL g1837 ( 
.A(n_1192),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1398),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1243),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1246),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1417),
.B(n_1054),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1324),
.Y(n_1842)
);

BUFx12f_ASAP7_75t_L g1843 ( 
.A(n_1423),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1393),
.B(n_728),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1325),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1330),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1331),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1248),
.B(n_762),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1133),
.B(n_762),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1423),
.Y(n_1850)
);

BUFx12f_ASAP7_75t_L g1851 ( 
.A(n_1428),
.Y(n_1851)
);

BUFx8_ASAP7_75t_SL g1852 ( 
.A(n_1215),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1428),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1429),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1429),
.B(n_767),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1332),
.Y(n_1856)
);

INVx6_ASAP7_75t_L g1857 ( 
.A(n_1184),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1253),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1510),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1524),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1694),
.B(n_1336),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1511),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1511),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1642),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1780),
.B(n_1434),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1780),
.B(n_1434),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1510),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1857),
.B(n_1145),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1512),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1828),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1541),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1829),
.A2(n_1215),
.B1(n_1247),
.B2(n_1245),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1839),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1840),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1510),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1510),
.Y(n_1876)
);

BUFx6f_ASAP7_75t_L g1877 ( 
.A(n_1515),
.Y(n_1877)
);

AND2x2_ASAP7_75t_SL g1878 ( 
.A(n_1829),
.B(n_1386),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1512),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1858),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1521),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1694),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1521),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1621),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1531),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1780),
.B(n_1449),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1642),
.Y(n_1887)
);

INVx3_ASAP7_75t_L g1888 ( 
.A(n_1541),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1541),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1515),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1558),
.B(n_1449),
.Y(n_1891)
);

XNOR2xp5_ASAP7_75t_L g1892 ( 
.A(n_1556),
.B(n_1245),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1531),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1572),
.B(n_1340),
.Y(n_1894)
);

BUFx8_ASAP7_75t_L g1895 ( 
.A(n_1516),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1621),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1533),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1515),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1541),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1558),
.B(n_1454),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1533),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1548),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1548),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1583),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1621),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1541),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1558),
.B(n_1454),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1578),
.B(n_1456),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1583),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1578),
.B(n_1585),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1621),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1857),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1629),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1638),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1629),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1578),
.B(n_1456),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1629),
.Y(n_1917)
);

OA21x2_ASAP7_75t_L g1918 ( 
.A1(n_1517),
.A2(n_1498),
.B(n_1342),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1629),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1638),
.Y(n_1920)
);

INVx3_ASAP7_75t_L g1921 ( 
.A(n_1549),
.Y(n_1921)
);

BUFx6f_ASAP7_75t_L g1922 ( 
.A(n_1515),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1644),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1525),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1688),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1688),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1688),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1688),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1690),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1658),
.B(n_1484),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1690),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1644),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1690),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1690),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1585),
.B(n_1484),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1655),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1655),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1525),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1525),
.Y(n_1939)
);

CKINVDCx16_ASAP7_75t_R g1940 ( 
.A(n_1676),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1655),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1549),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1857),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1655),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1655),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1679),
.B(n_1478),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1648),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_L g1948 ( 
.A(n_1857),
.B(n_1224),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1525),
.Y(n_1949)
);

AND2x2_ASAP7_75t_SL g1950 ( 
.A(n_1849),
.B(n_1824),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1572),
.Y(n_1951)
);

OA21x2_ASAP7_75t_L g1952 ( 
.A1(n_1517),
.A2(n_1480),
.B(n_1479),
.Y(n_1952)
);

BUFx8_ASAP7_75t_L g1953 ( 
.A(n_1516),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1589),
.B(n_1254),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1648),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1671),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1589),
.B(n_1255),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1671),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1549),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1671),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1585),
.B(n_1500),
.Y(n_1961)
);

INVx6_ASAP7_75t_L g1962 ( 
.A(n_1671),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1671),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1672),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1527),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1582),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1672),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1652),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1582),
.B(n_1341),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1549),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1672),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1592),
.B(n_1344),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1592),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1652),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1596),
.B(n_1345),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1664),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1658),
.B(n_1500),
.Y(n_1977)
);

INVx3_ASAP7_75t_L g1978 ( 
.A(n_1549),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1672),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1672),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1664),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1608),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1687),
.B(n_1256),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1527),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1775),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1554),
.Y(n_1986)
);

NAND2xp33_ASAP7_75t_SL g1987 ( 
.A(n_1855),
.B(n_1707),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1527),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1596),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1611),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1658),
.B(n_1224),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1607),
.B(n_1312),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1687),
.B(n_1703),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1614),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1667),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1667),
.Y(n_1996)
);

NOR2x1_ASAP7_75t_L g1997 ( 
.A(n_1805),
.B(n_1257),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1601),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1670),
.Y(n_1999)
);

CKINVDCx16_ASAP7_75t_R g2000 ( 
.A(n_1676),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1554),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1615),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1670),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1554),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1607),
.B(n_1312),
.Y(n_2005)
);

INVxp33_ASAP7_75t_SL g2006 ( 
.A(n_1536),
.Y(n_2006)
);

XOR2xp5_ASAP7_75t_L g2007 ( 
.A(n_1556),
.B(n_1247),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1601),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1680),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1616),
.Y(n_2010)
);

INVx3_ASAP7_75t_L g2011 ( 
.A(n_1554),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1687),
.B(n_1258),
.Y(n_2012)
);

BUFx6f_ASAP7_75t_L g2013 ( 
.A(n_1527),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1680),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1624),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1691),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1625),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1557),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1607),
.B(n_1314),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1703),
.B(n_1260),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_SL g2021 ( 
.A1(n_1542),
.A2(n_1262),
.B1(n_1275),
.B2(n_1259),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1703),
.B(n_1261),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_1623),
.B(n_1314),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1641),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1623),
.B(n_1320),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1623),
.B(n_1320),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1557),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1651),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1691),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1665),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1540),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1559),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1666),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1669),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1554),
.Y(n_2035)
);

OAI21x1_ASAP7_75t_L g2036 ( 
.A1(n_1545),
.A2(n_1483),
.B(n_1481),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1733),
.B(n_1184),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1733),
.B(n_1220),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1678),
.Y(n_2039)
);

BUFx6f_ASAP7_75t_L g2040 ( 
.A(n_1563),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1563),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1563),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1685),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1686),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1689),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1696),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1697),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1568),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1573),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1796),
.B(n_1350),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1704),
.Y(n_2051)
);

BUFx8_ASAP7_75t_L g2052 ( 
.A(n_1553),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1796),
.B(n_1350),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1796),
.B(n_1351),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1603),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1796),
.B(n_1351),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1603),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1713),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1715),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1775),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1720),
.Y(n_2061)
);

OR2x6_ASAP7_75t_L g2062 ( 
.A(n_1639),
.B(n_1159),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_SL g2063 ( 
.A(n_1838),
.B(n_1352),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_1654),
.B(n_1348),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1725),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1726),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1796),
.B(n_1373),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1806),
.B(n_1373),
.Y(n_2068)
);

BUFx2_ASAP7_75t_L g2069 ( 
.A(n_1654),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1563),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1575),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1806),
.B(n_1409),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1577),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1579),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1736),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1580),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_SL g2077 ( 
.A(n_1838),
.B(n_1352),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1666),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1806),
.B(n_1409),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1752),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1594),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1758),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1766),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1677),
.Y(n_2084)
);

INVx3_ASAP7_75t_L g2085 ( 
.A(n_1593),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1520),
.B(n_1793),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1565),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1806),
.B(n_741),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1776),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1799),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1793),
.B(n_1349),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1710),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1677),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1565),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_1710),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1793),
.B(n_1534),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1819),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1668),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_1733),
.B(n_1220),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1677),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_1707),
.A2(n_919),
.B1(n_1022),
.B2(n_913),
.Y(n_2101)
);

BUFx3_ASAP7_75t_L g2102 ( 
.A(n_1571),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1599),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1534),
.B(n_1353),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1617),
.B(n_1354),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1599),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1598),
.B(n_1232),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1668),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1675),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1675),
.Y(n_2110)
);

BUFx3_ASAP7_75t_L g2111 ( 
.A(n_1571),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1593),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1571),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1587),
.Y(n_2114)
);

BUFx6f_ASAP7_75t_L g2115 ( 
.A(n_1565),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1777),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1741),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_1617),
.B(n_1741),
.Y(n_2118)
);

OAI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_1707),
.A2(n_1130),
.B1(n_1122),
.B2(n_1422),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1806),
.B(n_751),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1600),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1765),
.Y(n_2122)
);

INVx5_ASAP7_75t_L g2123 ( 
.A(n_1526),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1765),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1788),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1546),
.B(n_759),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1598),
.B(n_1232),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1718),
.B(n_1252),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1600),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1606),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1788),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_1791),
.B(n_1355),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1606),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1791),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1724),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_SL g2136 ( 
.A(n_1838),
.B(n_1422),
.Y(n_2136)
);

NOR2x1_ASAP7_75t_L g2137 ( 
.A(n_1816),
.B(n_1844),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1724),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1529),
.B(n_1526),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1612),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1593),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1565),
.Y(n_2142)
);

INVxp67_ASAP7_75t_SL g2143 ( 
.A(n_1518),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_1804),
.Y(n_2144)
);

NOR3xp33_ASAP7_75t_L g2145 ( 
.A(n_1855),
.B(n_1250),
.C(n_1142),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1612),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1526),
.B(n_768),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1718),
.B(n_1104),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1613),
.Y(n_2149)
);

AND2x4_ASAP7_75t_L g2150 ( 
.A(n_1772),
.B(n_1357),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1718),
.B(n_1252),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1569),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1613),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1526),
.B(n_775),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1724),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1618),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1724),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1593),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1724),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1569),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1772),
.B(n_1296),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1770),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1569),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1618),
.Y(n_2164)
);

HB1xp67_ASAP7_75t_L g2165 ( 
.A(n_1777),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_1569),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1620),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1770),
.Y(n_2168)
);

BUFx6f_ASAP7_75t_L g2169 ( 
.A(n_1586),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1770),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_1778),
.B(n_1296),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1770),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1620),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1513),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1526),
.B(n_779),
.Y(n_2175)
);

BUFx8_ASAP7_75t_L g2176 ( 
.A(n_1553),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1586),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1514),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1673),
.B(n_1329),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_1818),
.A2(n_1443),
.B1(n_1465),
.B2(n_1424),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_1593),
.Y(n_2181)
);

INVx4_ASAP7_75t_L g2182 ( 
.A(n_1637),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1586),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1770),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1586),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1774),
.Y(n_2186)
);

AND2x6_ASAP7_75t_L g2187 ( 
.A(n_1848),
.B(n_1361),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1774),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1774),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1774),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_1825),
.B(n_1362),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1526),
.B(n_1547),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1588),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1804),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_1777),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1588),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1777),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1774),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1695),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1588),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1695),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1695),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1588),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1590),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1695),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1590),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1773),
.B(n_1363),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1705),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1692),
.B(n_1329),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1818),
.A2(n_1802),
.B1(n_1768),
.B2(n_1745),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1590),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1705),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1590),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1773),
.B(n_1365),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1705),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_1818),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1547),
.B(n_793),
.Y(n_2217)
);

BUFx6f_ASAP7_75t_L g2218 ( 
.A(n_1595),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1705),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1595),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1595),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1595),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_SL g2223 ( 
.A(n_1555),
.B(n_1584),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1609),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1708),
.Y(n_2225)
);

BUFx6f_ASAP7_75t_L g2226 ( 
.A(n_1609),
.Y(n_2226)
);

AND2x4_ASAP7_75t_L g2227 ( 
.A(n_1823),
.B(n_1366),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1609),
.Y(n_2228)
);

AND2x6_ASAP7_75t_L g2229 ( 
.A(n_1848),
.B(n_1370),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1609),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1708),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1619),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1547),
.B(n_816),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_1823),
.B(n_1347),
.Y(n_2234)
);

BUFx8_ASAP7_75t_L g2235 ( 
.A(n_1555),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1619),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1708),
.Y(n_2237)
);

OA21x2_ASAP7_75t_L g2238 ( 
.A1(n_1627),
.A2(n_1495),
.B(n_1372),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_1619),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1619),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1824),
.B(n_1347),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1818),
.A2(n_1443),
.B1(n_1465),
.B2(n_1424),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1528),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1547),
.B(n_817),
.Y(n_2244)
);

OAI22x1_ASAP7_75t_L g2245 ( 
.A1(n_2007),
.A2(n_1892),
.B1(n_2242),
.B2(n_2180),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2179),
.B(n_1818),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2104),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_2118),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2104),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2104),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2179),
.B(n_1818),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_L g2252 ( 
.A1(n_2241),
.A2(n_1824),
.B1(n_1547),
.B2(n_1728),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_1894),
.Y(n_2253)
);

INVx2_ASAP7_75t_SL g2254 ( 
.A(n_1894),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2209),
.B(n_1269),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_1950),
.B(n_1561),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2105),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2171),
.B(n_1802),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_2241),
.A2(n_1547),
.B1(n_1728),
.B2(n_1662),
.Y(n_2259)
);

INVx4_ASAP7_75t_L g2260 ( 
.A(n_2118),
.Y(n_2260)
);

AND3x1_ASAP7_75t_L g2261 ( 
.A(n_2145),
.B(n_1698),
.C(n_1717),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2107),
.B(n_1537),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2105),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2105),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_2118),
.Y(n_2265)
);

NAND2xp33_ASAP7_75t_R g2266 ( 
.A(n_2006),
.B(n_1826),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1914),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1914),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_1920),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1910),
.B(n_1551),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_2102),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1861),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1861),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1861),
.Y(n_2274)
);

NAND3xp33_ASAP7_75t_L g2275 ( 
.A(n_2171),
.B(n_2148),
.C(n_2209),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1882),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1993),
.B(n_1551),
.Y(n_2277)
);

BUFx3_ASAP7_75t_L g2278 ( 
.A(n_1912),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1982),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1990),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1920),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2096),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1994),
.Y(n_2283)
);

NAND2xp33_ASAP7_75t_L g2284 ( 
.A(n_2187),
.B(n_1056),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1923),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_SL g2286 ( 
.A(n_1950),
.B(n_1561),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2002),
.Y(n_2287)
);

NOR2x1p5_ASAP7_75t_L g2288 ( 
.A(n_1992),
.B(n_1566),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_1923),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2010),
.Y(n_2290)
);

NAND3xp33_ASAP7_75t_L g2291 ( 
.A(n_2148),
.B(n_1730),
.C(n_1727),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_1993),
.B(n_1633),
.Y(n_2292)
);

INVxp67_ASAP7_75t_SL g2293 ( 
.A(n_2102),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2096),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_SL g2295 ( 
.A(n_2062),
.Y(n_2295)
);

INVx8_ASAP7_75t_L g2296 ( 
.A(n_2187),
.Y(n_2296)
);

INVx1_ASAP7_75t_SL g2297 ( 
.A(n_2114),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_2111),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1932),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2187),
.B(n_1551),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1932),
.Y(n_2301)
);

INVx3_ASAP7_75t_L g2302 ( 
.A(n_2096),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_1987),
.A2(n_1744),
.B1(n_1763),
.B2(n_1742),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1947),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1864),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_1912),
.Y(n_2306)
);

AND3x2_ASAP7_75t_L g2307 ( 
.A(n_2216),
.B(n_1543),
.C(n_1634),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_1918),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2123),
.B(n_1633),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2187),
.B(n_1751),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2114),
.Y(n_2311)
);

INVx2_ASAP7_75t_SL g2312 ( 
.A(n_1894),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1985),
.B(n_1814),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1947),
.Y(n_2314)
);

AO21x2_ASAP7_75t_L g2315 ( 
.A1(n_2192),
.A2(n_2139),
.B(n_1937),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1955),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_1969),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1955),
.Y(n_2318)
);

BUFx3_ASAP7_75t_L g2319 ( 
.A(n_1951),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1864),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2015),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2060),
.B(n_1815),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2017),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_1865),
.B(n_1626),
.Y(n_2324)
);

NOR2x1p5_ASAP7_75t_L g2325 ( 
.A(n_2019),
.B(n_1566),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2024),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2187),
.B(n_1751),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2028),
.Y(n_2328)
);

INVx8_ASAP7_75t_L g2329 ( 
.A(n_2187),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_1918),
.Y(n_2330)
);

NAND2xp33_ASAP7_75t_L g2331 ( 
.A(n_2229),
.B(n_1056),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_2123),
.B(n_1537),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_2123),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_1887),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_1951),
.Y(n_2335)
);

NAND2xp33_ASAP7_75t_R g2336 ( 
.A(n_2006),
.B(n_1826),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2229),
.B(n_1643),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1968),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2123),
.B(n_1656),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_L g2340 ( 
.A(n_2229),
.B(n_1056),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2030),
.Y(n_2341)
);

AO21x2_ASAP7_75t_L g2342 ( 
.A1(n_1936),
.A2(n_1809),
.B(n_1753),
.Y(n_2342)
);

INVx3_ASAP7_75t_L g2343 ( 
.A(n_1918),
.Y(n_2343)
);

NAND3xp33_ASAP7_75t_L g2344 ( 
.A(n_2128),
.B(n_1822),
.C(n_1782),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2034),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_1973),
.Y(n_2346)
);

BUFx4f_ASAP7_75t_L g2347 ( 
.A(n_2062),
.Y(n_2347)
);

INVx4_ASAP7_75t_L g2348 ( 
.A(n_2123),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_1969),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2039),
.Y(n_2350)
);

NOR2x1p5_ASAP7_75t_L g2351 ( 
.A(n_2025),
.B(n_1584),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2043),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_2119),
.B(n_1544),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2044),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1968),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2111),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2045),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2046),
.Y(n_2358)
);

INVx1_ASAP7_75t_SL g2359 ( 
.A(n_2107),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_1860),
.B(n_1544),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1974),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_1887),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_2216),
.B(n_1656),
.Y(n_2363)
);

NAND2xp33_ASAP7_75t_R g2364 ( 
.A(n_2128),
.B(n_1853),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2047),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2051),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1974),
.Y(n_2367)
);

AND2x2_ASAP7_75t_SL g2368 ( 
.A(n_1878),
.B(n_1662),
.Y(n_2368)
);

INVx5_ASAP7_75t_L g2369 ( 
.A(n_2243),
.Y(n_2369)
);

INVx2_ASAP7_75t_SL g2370 ( 
.A(n_1969),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_1952),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_SL g2372 ( 
.A(n_2062),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2026),
.B(n_1682),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1976),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2058),
.Y(n_2375)
);

INVx4_ASAP7_75t_L g2376 ( 
.A(n_1973),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2229),
.B(n_1702),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_1976),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1981),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1981),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2229),
.B(n_1762),
.Y(n_2381)
);

INVx3_ASAP7_75t_L g2382 ( 
.A(n_1952),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2229),
.B(n_2151),
.Y(n_2383)
);

BUFx3_ASAP7_75t_L g2384 ( 
.A(n_1989),
.Y(n_2384)
);

INVx1_ASAP7_75t_SL g2385 ( 
.A(n_2127),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2059),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2151),
.B(n_1764),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1995),
.Y(n_2388)
);

AOI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2113),
.A2(n_1728),
.B1(n_1731),
.B2(n_1662),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2061),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2065),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_SL g2392 ( 
.A1(n_1878),
.A2(n_1523),
.B1(n_1574),
.B2(n_1309),
.Y(n_2392)
);

BUFx6f_ASAP7_75t_L g2393 ( 
.A(n_2113),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2066),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2075),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_1995),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_1866),
.B(n_1610),
.Y(n_2397)
);

INVx4_ASAP7_75t_L g2398 ( 
.A(n_1962),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1996),
.Y(n_2399)
);

OAI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_1935),
.A2(n_1604),
.B1(n_1722),
.B2(n_1683),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1996),
.Y(n_2401)
);

OR2x6_ASAP7_75t_L g2402 ( 
.A(n_2062),
.B(n_1639),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_1999),
.Y(n_2403)
);

OR2x6_ASAP7_75t_L g2404 ( 
.A(n_2021),
.B(n_1650),
.Y(n_2404)
);

OAI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2210),
.A2(n_1961),
.B1(n_1891),
.B2(n_1907),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_1987),
.A2(n_1854),
.B1(n_1853),
.B2(n_1657),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_SL g2407 ( 
.A(n_2037),
.B(n_1682),
.Y(n_2407)
);

INVx5_ASAP7_75t_L g2408 ( 
.A(n_2243),
.Y(n_2408)
);

CKINVDCx5p33_ASAP7_75t_R g2409 ( 
.A(n_2092),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_1999),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2003),
.Y(n_2411)
);

BUFx4f_ASAP7_75t_L g2412 ( 
.A(n_2037),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2080),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_2092),
.Y(n_2414)
);

BUFx10_ASAP7_75t_L g2415 ( 
.A(n_2194),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2082),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2083),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2003),
.Y(n_2418)
);

XOR2x2_ASAP7_75t_L g2419 ( 
.A(n_1892),
.B(n_1681),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_SL g2420 ( 
.A(n_2038),
.B(n_1854),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_2194),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2009),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2009),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2089),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2038),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2099),
.B(n_1767),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_1972),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2090),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_L g2429 ( 
.A(n_1886),
.B(n_1908),
.C(n_1900),
.Y(n_2429)
);

OR2x6_ASAP7_75t_L g2430 ( 
.A(n_1872),
.B(n_1650),
.Y(n_2430)
);

AND2x4_ASAP7_75t_L g2431 ( 
.A(n_2098),
.B(n_1729),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2097),
.Y(n_2432)
);

INVx3_ASAP7_75t_L g2433 ( 
.A(n_1952),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2099),
.B(n_1735),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_L g2435 ( 
.A1(n_2238),
.A2(n_1794),
.B1(n_1731),
.B2(n_1419),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_1916),
.B(n_1735),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_1989),
.Y(n_2437)
);

INVx8_ASAP7_75t_L g2438 ( 
.A(n_2086),
.Y(n_2438)
);

OAI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2063),
.A2(n_1358),
.B1(n_1470),
.B2(n_1419),
.Y(n_2439)
);

AOI21x1_ASAP7_75t_L g2440 ( 
.A1(n_1941),
.A2(n_1945),
.B(n_1944),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1870),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2127),
.B(n_1735),
.Y(n_2442)
);

INVxp67_ASAP7_75t_SL g2443 ( 
.A(n_1943),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2161),
.B(n_1523),
.Y(n_2444)
);

BUFx10_ASAP7_75t_L g2445 ( 
.A(n_1948),
.Y(n_2445)
);

OR2x6_ASAP7_75t_L g2446 ( 
.A(n_2055),
.B(n_1699),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2014),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1873),
.Y(n_2448)
);

INVx5_ASAP7_75t_L g2449 ( 
.A(n_2243),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2137),
.B(n_1735),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2126),
.B(n_2086),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2014),
.Y(n_2452)
);

INVx1_ASAP7_75t_SL g2453 ( 
.A(n_2161),
.Y(n_2453)
);

BUFx4f_ASAP7_75t_L g2454 ( 
.A(n_2086),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1874),
.Y(n_2455)
);

INVxp67_ASAP7_75t_R g2456 ( 
.A(n_2234),
.Y(n_2456)
);

INVx5_ASAP7_75t_L g2457 ( 
.A(n_2243),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1868),
.B(n_2234),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2016),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_1991),
.B(n_1735),
.Y(n_2460)
);

INVx3_ASAP7_75t_L g2461 ( 
.A(n_2121),
.Y(n_2461)
);

BUFx2_ASAP7_75t_L g2462 ( 
.A(n_2055),
.Y(n_2462)
);

CKINVDCx11_ASAP7_75t_R g2463 ( 
.A(n_2033),
.Y(n_2463)
);

OR2x2_ASAP7_75t_L g2464 ( 
.A(n_1991),
.B(n_1647),
.Y(n_2464)
);

INVx2_ASAP7_75t_SL g2465 ( 
.A(n_1972),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1880),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2016),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_1930),
.B(n_1628),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2036),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2036),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2121),
.Y(n_2471)
);

INVx4_ASAP7_75t_L g2472 ( 
.A(n_1962),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2129),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2029),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_1972),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_1948),
.B(n_1761),
.Y(n_2476)
);

AND2x6_ASAP7_75t_L g2477 ( 
.A(n_1997),
.B(n_1795),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2029),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_1930),
.B(n_1645),
.Y(n_2479)
);

INVx4_ASAP7_75t_L g2480 ( 
.A(n_1962),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_1862),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_2057),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_SL g2483 ( 
.A(n_1977),
.B(n_1761),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_1862),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_1859),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_1977),
.B(n_1653),
.Y(n_2486)
);

OR2x2_ASAP7_75t_L g2487 ( 
.A(n_1940),
.B(n_1647),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2005),
.B(n_1761),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_1868),
.B(n_1777),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1975),
.Y(n_2490)
);

OR2x6_ASAP7_75t_L g2491 ( 
.A(n_2057),
.B(n_1699),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_2000),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1863),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1975),
.Y(n_2494)
);

INVx2_ASAP7_75t_SL g2495 ( 
.A(n_1975),
.Y(n_2495)
);

BUFx6f_ASAP7_75t_SL g2496 ( 
.A(n_2064),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1863),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_1869),
.Y(n_2498)
);

AOI21x1_ASAP7_75t_L g2499 ( 
.A1(n_1956),
.A2(n_1552),
.B(n_1545),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2005),
.B(n_1660),
.Y(n_2500)
);

INVx5_ASAP7_75t_L g2501 ( 
.A(n_2243),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2023),
.B(n_1761),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_2129),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_1869),
.Y(n_2504)
);

INVx2_ASAP7_75t_SL g2505 ( 
.A(n_2064),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2064),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2132),
.Y(n_2507)
);

NAND2xp33_ASAP7_75t_L g2508 ( 
.A(n_2191),
.B(n_1056),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_1879),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2132),
.Y(n_2510)
);

BUFx3_ASAP7_75t_L g2511 ( 
.A(n_2069),
.Y(n_2511)
);

INVx1_ASAP7_75t_SL g2512 ( 
.A(n_2007),
.Y(n_2512)
);

BUFx4f_ASAP7_75t_L g2513 ( 
.A(n_2069),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2130),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2132),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2174),
.Y(n_2516)
);

OAI21xp33_ASAP7_75t_SL g2517 ( 
.A1(n_2023),
.A2(n_1640),
.B(n_1627),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2091),
.B(n_1657),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_1879),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_1881),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_1983),
.B(n_1761),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_1966),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_1881),
.Y(n_2523)
);

AOI21x1_ASAP7_75t_L g2524 ( 
.A1(n_1958),
.A2(n_1552),
.B(n_1640),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_1998),
.B(n_1663),
.Y(n_2525)
);

OAI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2077),
.A2(n_2136),
.B1(n_1358),
.B2(n_1470),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_1983),
.B(n_1771),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2174),
.Y(n_2528)
);

INVx5_ASAP7_75t_L g2529 ( 
.A(n_2182),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2178),
.Y(n_2530)
);

OR2x6_ASAP7_75t_L g2531 ( 
.A(n_2008),
.B(n_1712),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_1883),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_1883),
.Y(n_2533)
);

CKINVDCx5p33_ASAP7_75t_R g2534 ( 
.A(n_2033),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2178),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_1885),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2108),
.B(n_1684),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_1885),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2109),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2012),
.B(n_1771),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2091),
.B(n_1693),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2091),
.B(n_1693),
.Y(n_2542)
);

INVxp67_ASAP7_75t_SL g2543 ( 
.A(n_1965),
.Y(n_2543)
);

INVx5_ASAP7_75t_L g2544 ( 
.A(n_2182),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2110),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2117),
.B(n_1739),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2238),
.A2(n_1731),
.B1(n_1794),
.B2(n_1661),
.Y(n_2547)
);

NAND2xp33_ASAP7_75t_R g2548 ( 
.A(n_2012),
.B(n_1709),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_1895),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2122),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_1893),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_1895),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2020),
.B(n_1771),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_1893),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2124),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_1897),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2125),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_1897),
.Y(n_2558)
);

INVx5_ASAP7_75t_L g2559 ( 
.A(n_2182),
.Y(n_2559)
);

INVx4_ASAP7_75t_L g2560 ( 
.A(n_1962),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2131),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2134),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_2020),
.B(n_2022),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2031),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2130),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2150),
.B(n_1771),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_1901),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2022),
.B(n_1771),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_1901),
.Y(n_2569)
);

OR2x6_ASAP7_75t_L g2570 ( 
.A(n_1946),
.B(n_1712),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_1954),
.B(n_1755),
.Y(n_2571)
);

INVx5_ASAP7_75t_L g2572 ( 
.A(n_2013),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_1902),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_1902),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_1859),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_1903),
.Y(n_2576)
);

INVx5_ASAP7_75t_L g2577 ( 
.A(n_2013),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_1903),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_1954),
.B(n_1757),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_1904),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_1895),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2150),
.B(n_1709),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_1957),
.Y(n_2583)
);

INVx3_ASAP7_75t_L g2584 ( 
.A(n_2133),
.Y(n_2584)
);

INVxp33_ASAP7_75t_SL g2585 ( 
.A(n_2223),
.Y(n_2585)
);

NOR2x1p5_ASAP7_75t_L g2586 ( 
.A(n_2050),
.B(n_1602),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2031),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2032),
.Y(n_2588)
);

BUFx16f_ASAP7_75t_R g2589 ( 
.A(n_1953),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2150),
.B(n_1719),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2143),
.B(n_1674),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_1904),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_1909),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2207),
.B(n_2214),
.Y(n_2594)
);

INVx2_ASAP7_75t_SL g2595 ( 
.A(n_1957),
.Y(n_2595)
);

BUFx10_ASAP7_75t_L g2596 ( 
.A(n_2207),
.Y(n_2596)
);

AOI22xp33_ASAP7_75t_L g2597 ( 
.A1(n_2238),
.A2(n_1794),
.B1(n_2214),
.B2(n_2207),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2032),
.Y(n_2598)
);

AO22x2_ASAP7_75t_L g2599 ( 
.A1(n_2214),
.A2(n_1519),
.B1(n_1769),
.B2(n_1706),
.Y(n_2599)
);

AO22x2_ASAP7_75t_L g2600 ( 
.A1(n_2227),
.A2(n_1841),
.B1(n_1701),
.B2(n_1083),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_1884),
.B(n_1622),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2048),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_1909),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_1896),
.B(n_1622),
.Y(n_2604)
);

INVx2_ASAP7_75t_SL g2605 ( 
.A(n_2227),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2048),
.Y(n_2606)
);

BUFx10_ASAP7_75t_L g2607 ( 
.A(n_2227),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2049),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_1953),
.Y(n_2609)
);

INVxp33_ASAP7_75t_L g2610 ( 
.A(n_2116),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1953),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2103),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2049),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2071),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_L g2615 ( 
.A(n_2054),
.B(n_1833),
.C(n_1808),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2101),
.B(n_1836),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2071),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2133),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2103),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2073),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2073),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2074),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2074),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2106),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2106),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2140),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2140),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_1859),
.Y(n_2628)
);

INVx2_ASAP7_75t_SL g2629 ( 
.A(n_2165),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2199),
.B(n_1719),
.Y(n_2630)
);

BUFx10_ASAP7_75t_L g2631 ( 
.A(n_2195),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2146),
.Y(n_2632)
);

INVx3_ASAP7_75t_L g2633 ( 
.A(n_2265),
.Y(n_2633)
);

CKINVDCx20_ASAP7_75t_R g2634 ( 
.A(n_2463),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2247),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2297),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2319),
.B(n_2197),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2247),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2258),
.B(n_1732),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2319),
.B(n_1905),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2387),
.B(n_2053),
.Y(n_2641)
);

AND2x4_ASAP7_75t_L g2642 ( 
.A(n_2335),
.B(n_1911),
.Y(n_2642)
);

OAI221xp5_ASAP7_75t_L g2643 ( 
.A1(n_2275),
.A2(n_1841),
.B1(n_1813),
.B2(n_1785),
.C(n_1732),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2249),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2249),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2250),
.Y(n_2646)
);

AND2x6_ASAP7_75t_L g2647 ( 
.A(n_2271),
.B(n_1960),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2250),
.Y(n_2648)
);

BUFx3_ASAP7_75t_L g2649 ( 
.A(n_2522),
.Y(n_2649)
);

OR2x6_ASAP7_75t_L g2650 ( 
.A(n_2402),
.B(n_1803),
.Y(n_2650)
);

AOI22xp33_ASAP7_75t_L g2651 ( 
.A1(n_2368),
.A2(n_2202),
.B1(n_2205),
.B2(n_2201),
.Y(n_2651)
);

INVx6_ASAP7_75t_L g2652 ( 
.A(n_2415),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2335),
.B(n_2346),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_2258),
.B(n_1785),
.Y(n_2654)
);

AND2x6_ASAP7_75t_L g2655 ( 
.A(n_2271),
.B(n_1963),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2257),
.Y(n_2656)
);

AND2x6_ASAP7_75t_L g2657 ( 
.A(n_2271),
.B(n_2298),
.Y(n_2657)
);

OAI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_2246),
.A2(n_2056),
.B1(n_2068),
.B2(n_2067),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2263),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2264),
.Y(n_2660)
);

NAND2xp33_ASAP7_75t_L g2661 ( 
.A(n_2271),
.B(n_2298),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2282),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2265),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2282),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2462),
.Y(n_2665)
);

INVx1_ASAP7_75t_SL g2666 ( 
.A(n_2360),
.Y(n_2666)
);

AND2x2_ASAP7_75t_SL g2667 ( 
.A(n_2261),
.B(n_1813),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2294),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2272),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2294),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2273),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2302),
.Y(n_2672)
);

NAND2x1p5_ASAP7_75t_L g2673 ( 
.A(n_2278),
.B(n_2054),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2412),
.B(n_2303),
.Y(n_2674)
);

AOI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2324),
.A2(n_1913),
.B1(n_1917),
.B2(n_1915),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2274),
.Y(n_2676)
);

INVx4_ASAP7_75t_L g2677 ( 
.A(n_2265),
.Y(n_2677)
);

BUFx6f_ASAP7_75t_L g2678 ( 
.A(n_2265),
.Y(n_2678)
);

AND2x2_ASAP7_75t_SL g2679 ( 
.A(n_2347),
.B(n_1634),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2612),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2612),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2302),
.Y(n_2682)
);

INVx2_ASAP7_75t_SL g2683 ( 
.A(n_2518),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2262),
.B(n_2571),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2267),
.Y(n_2685)
);

OAI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2251),
.A2(n_2072),
.B1(n_2079),
.B2(n_1850),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2255),
.B(n_1259),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2291),
.B(n_1262),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2619),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2298),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2619),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2624),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2267),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2313),
.B(n_1275),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2346),
.B(n_1919),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2624),
.Y(n_2696)
);

AND2x6_ASAP7_75t_L g2697 ( 
.A(n_2298),
.B(n_1964),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2625),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2268),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_2522),
.Y(n_2700)
);

INVxp67_ASAP7_75t_L g2701 ( 
.A(n_2571),
.Y(n_2701)
);

BUFx6f_ASAP7_75t_L g2702 ( 
.A(n_2356),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2453),
.B(n_1538),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2324),
.B(n_1925),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2268),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2625),
.Y(n_2706)
);

OR2x2_ASAP7_75t_SL g2707 ( 
.A(n_2353),
.B(n_1550),
.Y(n_2707)
);

INVx4_ASAP7_75t_SL g2708 ( 
.A(n_2295),
.Y(n_2708)
);

AND2x4_ASAP7_75t_L g2709 ( 
.A(n_2278),
.B(n_2306),
.Y(n_2709)
);

AND2x6_ASAP7_75t_L g2710 ( 
.A(n_2356),
.B(n_1967),
.Y(n_2710)
);

INVx4_ASAP7_75t_L g2711 ( 
.A(n_2356),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2564),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2269),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2269),
.Y(n_2714)
);

AND2x4_ASAP7_75t_L g2715 ( 
.A(n_2306),
.B(n_1926),
.Y(n_2715)
);

NAND2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2454),
.B(n_1729),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2426),
.B(n_1927),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2579),
.B(n_1636),
.Y(n_2718)
);

NAND2xp33_ASAP7_75t_L g2719 ( 
.A(n_2356),
.B(n_1659),
.Y(n_2719)
);

INVx2_ASAP7_75t_SL g2720 ( 
.A(n_2541),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2463),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2587),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2313),
.B(n_1309),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2281),
.Y(n_2724)
);

NAND2x1p5_ASAP7_75t_L g2725 ( 
.A(n_2454),
.B(n_1729),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2588),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2598),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2602),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2384),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2579),
.B(n_1636),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2393),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2606),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2376),
.B(n_1928),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2393),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2281),
.Y(n_2735)
);

BUFx2_ASAP7_75t_L g2736 ( 
.A(n_2311),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2608),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2458),
.B(n_1929),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2613),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2614),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2285),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2617),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2393),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2293),
.B(n_1931),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2285),
.Y(n_2745)
);

NOR2xp33_ASAP7_75t_L g2746 ( 
.A(n_2322),
.B(n_1321),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2289),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2620),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2376),
.B(n_1933),
.Y(n_2749)
);

INVx2_ASAP7_75t_SL g2750 ( 
.A(n_2542),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2464),
.Y(n_2751)
);

INVx3_ASAP7_75t_L g2752 ( 
.A(n_2248),
.Y(n_2752)
);

INVx1_ASAP7_75t_SL g2753 ( 
.A(n_2492),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2412),
.B(n_1574),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_L g2755 ( 
.A(n_2322),
.B(n_1321),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2359),
.B(n_1934),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2320),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2289),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2385),
.B(n_2208),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2591),
.B(n_2212),
.Y(n_2760)
);

NOR2xp33_ASAP7_75t_L g2761 ( 
.A(n_2397),
.B(n_1339),
.Y(n_2761)
);

BUFx6f_ASAP7_75t_L g2762 ( 
.A(n_2393),
.Y(n_2762)
);

AOI22xp5_ASAP7_75t_L g2763 ( 
.A1(n_2368),
.A2(n_2219),
.B1(n_2225),
.B2(n_2215),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2299),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2384),
.Y(n_2765)
);

INVx4_ASAP7_75t_L g2766 ( 
.A(n_2438),
.Y(n_2766)
);

BUFx6f_ASAP7_75t_L g2767 ( 
.A(n_2438),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2299),
.Y(n_2768)
);

INVxp67_ASAP7_75t_SL g2769 ( 
.A(n_2248),
.Y(n_2769)
);

HB1xp67_ASAP7_75t_L g2770 ( 
.A(n_2437),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2301),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2397),
.B(n_1339),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2301),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_SL g2774 ( 
.A(n_2526),
.B(n_1574),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2260),
.Y(n_2775)
);

INVxp67_ASAP7_75t_SL g2776 ( 
.A(n_2260),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_2605),
.B(n_2231),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2621),
.Y(n_2778)
);

INVx1_ASAP7_75t_SL g2779 ( 
.A(n_2487),
.Y(n_2779)
);

INVxp67_ASAP7_75t_L g2780 ( 
.A(n_2525),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2622),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2405),
.B(n_2237),
.Y(n_2782)
);

AO22x2_ASAP7_75t_L g2783 ( 
.A1(n_2400),
.A2(n_2078),
.B1(n_2144),
.B2(n_2095),
.Y(n_2783)
);

INVx1_ASAP7_75t_SL g2784 ( 
.A(n_2437),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2304),
.Y(n_2785)
);

INVx4_ASAP7_75t_L g2786 ( 
.A(n_2438),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2304),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2253),
.B(n_1820),
.Y(n_2788)
);

AO22x2_ASAP7_75t_L g2789 ( 
.A1(n_2344),
.A2(n_1649),
.B1(n_1280),
.B2(n_1288),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2254),
.B(n_1820),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2314),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2314),
.Y(n_2792)
);

INVxp67_ASAP7_75t_SL g2793 ( 
.A(n_2485),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2316),
.Y(n_2794)
);

NAND2x1p5_ASAP7_75t_L g2795 ( 
.A(n_2482),
.B(n_1971),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2316),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_L g2797 ( 
.A(n_2500),
.B(n_1467),
.Y(n_2797)
);

BUFx2_ASAP7_75t_L g2798 ( 
.A(n_2482),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2318),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2623),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2312),
.B(n_1821),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2516),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2405),
.B(n_1979),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2528),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2530),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2535),
.Y(n_2806)
);

OR2x2_ASAP7_75t_SL g2807 ( 
.A(n_2615),
.B(n_1570),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2456),
.B(n_1576),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2451),
.B(n_1980),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2318),
.Y(n_2810)
);

INVx5_ASAP7_75t_L g2811 ( 
.A(n_2446),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2338),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_2334),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2500),
.B(n_2468),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2485),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2468),
.B(n_1467),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2317),
.B(n_1821),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2338),
.Y(n_2818)
);

INVx6_ASAP7_75t_L g2819 ( 
.A(n_2415),
.Y(n_2819)
);

INVx4_ASAP7_75t_L g2820 ( 
.A(n_2485),
.Y(n_2820)
);

AND2x6_ASAP7_75t_L g2821 ( 
.A(n_2383),
.B(n_2146),
.Y(n_2821)
);

OR2x6_ASAP7_75t_L g2822 ( 
.A(n_2402),
.B(n_1803),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2355),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2355),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_2409),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2361),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2479),
.B(n_1476),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2361),
.Y(n_2828)
);

AND2x4_ASAP7_75t_L g2829 ( 
.A(n_2349),
.B(n_1827),
.Y(n_2829)
);

INVx4_ASAP7_75t_L g2830 ( 
.A(n_2485),
.Y(n_2830)
);

OR2x6_ASAP7_75t_L g2831 ( 
.A(n_2402),
.B(n_1843),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2367),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2370),
.B(n_1827),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2367),
.Y(n_2834)
);

INVx3_ASAP7_75t_L g2835 ( 
.A(n_2575),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2479),
.B(n_1476),
.Y(n_2836)
);

AND2x4_ASAP7_75t_L g2837 ( 
.A(n_2427),
.B(n_1834),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2374),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2486),
.B(n_1493),
.Y(n_2839)
);

NOR2xp33_ASAP7_75t_L g2840 ( 
.A(n_2486),
.B(n_1493),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2575),
.Y(n_2841)
);

AND2x6_ASAP7_75t_L g2842 ( 
.A(n_2308),
.B(n_2149),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2575),
.Y(n_2843)
);

AND2x6_ASAP7_75t_L g2844 ( 
.A(n_2308),
.B(n_2149),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2374),
.Y(n_2845)
);

INVx3_ASAP7_75t_L g2846 ( 
.A(n_2575),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_2526),
.B(n_1659),
.Y(n_2847)
);

INVxp67_ASAP7_75t_L g2848 ( 
.A(n_2525),
.Y(n_2848)
);

BUFx3_ASAP7_75t_L g2849 ( 
.A(n_2511),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2563),
.B(n_2084),
.Y(n_2850)
);

BUFx6f_ASAP7_75t_L g2851 ( 
.A(n_2628),
.Y(n_2851)
);

A2O1A1Ixp33_ASAP7_75t_L g2852 ( 
.A1(n_2429),
.A2(n_1753),
.B(n_1809),
.C(n_2147),
.Y(n_2852)
);

BUFx2_ASAP7_75t_L g2853 ( 
.A(n_2511),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2489),
.B(n_2084),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_2420),
.B(n_1591),
.Y(n_2855)
);

AND2x4_ASAP7_75t_L g2856 ( 
.A(n_2465),
.B(n_1834),
.Y(n_2856)
);

OR2x6_ASAP7_75t_L g2857 ( 
.A(n_2446),
.B(n_1843),
.Y(n_2857)
);

CKINVDCx11_ASAP7_75t_R g2858 ( 
.A(n_2589),
.Y(n_2858)
);

BUFx3_ASAP7_75t_L g2859 ( 
.A(n_2513),
.Y(n_2859)
);

BUFx3_ASAP7_75t_L g2860 ( 
.A(n_2513),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2420),
.B(n_1851),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2378),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2425),
.B(n_1851),
.Y(n_2863)
);

AND2x2_ASAP7_75t_L g2864 ( 
.A(n_2583),
.B(n_1602),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2378),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2379),
.Y(n_2866)
);

AOI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2256),
.A2(n_2076),
.B1(n_2081),
.B2(n_2135),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2379),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2628),
.Y(n_2869)
);

BUFx6f_ASAP7_75t_L g2870 ( 
.A(n_2628),
.Y(n_2870)
);

NAND3xp33_ASAP7_75t_L g2871 ( 
.A(n_2616),
.B(n_2176),
.C(n_2052),
.Y(n_2871)
);

BUFx6f_ASAP7_75t_L g2872 ( 
.A(n_2628),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2380),
.Y(n_2873)
);

AND2x4_ASAP7_75t_L g2874 ( 
.A(n_2475),
.B(n_2495),
.Y(n_2874)
);

BUFx6f_ASAP7_75t_L g2875 ( 
.A(n_2596),
.Y(n_2875)
);

AND2x6_ASAP7_75t_L g2876 ( 
.A(n_2330),
.B(n_2153),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2380),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2445),
.B(n_1631),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2595),
.B(n_2093),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2388),
.Y(n_2880)
);

NOR2x1p5_ASAP7_75t_L g2881 ( 
.A(n_2549),
.B(n_1631),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2388),
.Y(n_2882)
);

AND2x2_ASAP7_75t_L g2883 ( 
.A(n_2444),
.B(n_1810),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_SL g2884 ( 
.A(n_2439),
.B(n_2596),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2505),
.B(n_1835),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2279),
.B(n_2093),
.Y(n_2886)
);

BUFx6f_ASAP7_75t_L g2887 ( 
.A(n_2607),
.Y(n_2887)
);

BUFx3_ASAP7_75t_L g2888 ( 
.A(n_2414),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2396),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2256),
.A2(n_2076),
.B1(n_2081),
.B2(n_2138),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2537),
.B(n_1810),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2280),
.B(n_2100),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2286),
.A2(n_2157),
.B1(n_2159),
.B2(n_2155),
.Y(n_2893)
);

OAI22xp5_ASAP7_75t_SL g2894 ( 
.A1(n_2512),
.A2(n_2245),
.B1(n_2392),
.B2(n_2585),
.Y(n_2894)
);

INVx4_ASAP7_75t_L g2895 ( 
.A(n_2607),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2396),
.Y(n_2896)
);

CKINVDCx16_ASAP7_75t_R g2897 ( 
.A(n_2548),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2399),
.Y(n_2898)
);

BUFx2_ASAP7_75t_L g2899 ( 
.A(n_2446),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2399),
.Y(n_2900)
);

INVx4_ASAP7_75t_L g2901 ( 
.A(n_2296),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2401),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2582),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2401),
.Y(n_2904)
);

OR2x6_ASAP7_75t_L g2905 ( 
.A(n_2491),
.B(n_2052),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2445),
.B(n_1837),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2403),
.Y(n_2907)
);

AND2x6_ASAP7_75t_L g2908 ( 
.A(n_2330),
.B(n_2153),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2403),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2286),
.A2(n_2168),
.B1(n_2170),
.B2(n_2162),
.Y(n_2910)
);

INVx3_ASAP7_75t_L g2911 ( 
.A(n_2440),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2410),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2631),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2410),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2537),
.B(n_1274),
.Y(n_2915)
);

AND2x6_ASAP7_75t_L g2916 ( 
.A(n_2343),
.B(n_2156),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2411),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2411),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2418),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2418),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2631),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2407),
.B(n_1837),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2422),
.Y(n_2923)
);

OR2x2_ASAP7_75t_L g2924 ( 
.A(n_2582),
.B(n_1389),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2422),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2423),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2546),
.B(n_1397),
.Y(n_2927)
);

INVx3_ASAP7_75t_L g2928 ( 
.A(n_2423),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2507),
.B(n_1835),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2447),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2447),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2452),
.Y(n_2932)
);

INVx5_ASAP7_75t_L g2933 ( 
.A(n_2491),
.Y(n_2933)
);

AND2x4_ASAP7_75t_L g2934 ( 
.A(n_2510),
.B(n_1847),
.Y(n_2934)
);

AND2x4_ASAP7_75t_L g2935 ( 
.A(n_2515),
.B(n_2490),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_2494),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2452),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2407),
.B(n_1852),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2364),
.A2(n_2175),
.B1(n_2217),
.B2(n_2154),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2506),
.B(n_1847),
.Y(n_2940)
);

INVx4_ASAP7_75t_L g2941 ( 
.A(n_2296),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_L g2942 ( 
.A1(n_2616),
.A2(n_2594),
.B1(n_2597),
.B2(n_2287),
.Y(n_2942)
);

OAI221xp5_ASAP7_75t_L g2943 ( 
.A1(n_2594),
.A2(n_1496),
.B1(n_1453),
.B2(n_1723),
.C(n_1721),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2283),
.B(n_2290),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2373),
.B(n_1852),
.Y(n_2945)
);

AND2x4_ASAP7_75t_L g2946 ( 
.A(n_2443),
.B(n_1856),
.Y(n_2946)
);

OAI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2597),
.A2(n_2244),
.B1(n_2233),
.B2(n_2088),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2459),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2459),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2467),
.Y(n_2950)
);

AO21x2_ASAP7_75t_L g2951 ( 
.A1(n_2337),
.A2(n_2184),
.B(n_2172),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2467),
.Y(n_2952)
);

OR2x6_ASAP7_75t_L g2953 ( 
.A(n_2491),
.B(n_2052),
.Y(n_2953)
);

AND2x4_ASAP7_75t_L g2954 ( 
.A(n_2539),
.B(n_1856),
.Y(n_2954)
);

INVx4_ASAP7_75t_L g2955 ( 
.A(n_2296),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2474),
.Y(n_2956)
);

INVx2_ASAP7_75t_SL g2957 ( 
.A(n_2545),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2474),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2550),
.B(n_1371),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2478),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2478),
.Y(n_2961)
);

BUFx6f_ASAP7_75t_L g2962 ( 
.A(n_2629),
.Y(n_2962)
);

INVxp67_ASAP7_75t_SL g2963 ( 
.A(n_2543),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2481),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2321),
.B(n_2100),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2481),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2439),
.B(n_2120),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2546),
.B(n_1842),
.Y(n_2968)
);

OAI21xp33_ASAP7_75t_L g2969 ( 
.A1(n_2406),
.A2(n_830),
.B(n_823),
.Y(n_2969)
);

OR2x2_ASAP7_75t_L g2970 ( 
.A(n_2590),
.B(n_1842),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2252),
.A2(n_2188),
.B1(n_2189),
.B2(n_2186),
.Y(n_2971)
);

INVx1_ASAP7_75t_SL g2972 ( 
.A(n_2590),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_2484),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2323),
.B(n_2190),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2484),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2493),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2610),
.B(n_1842),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2373),
.B(n_1564),
.Y(n_2978)
);

OAI21xp33_ASAP7_75t_L g2979 ( 
.A1(n_2610),
.A2(n_833),
.B(n_832),
.Y(n_2979)
);

INVx1_ASAP7_75t_SL g2980 ( 
.A(n_2421),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2531),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2555),
.B(n_2557),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2493),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2497),
.Y(n_2984)
);

BUFx3_ASAP7_75t_L g2985 ( 
.A(n_2531),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2561),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2497),
.Y(n_2987)
);

HB1xp67_ASAP7_75t_L g2988 ( 
.A(n_2548),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2498),
.Y(n_2989)
);

BUFx6f_ASAP7_75t_L g2990 ( 
.A(n_2431),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2326),
.B(n_2328),
.Y(n_2991)
);

AO22x2_ASAP7_75t_L g2992 ( 
.A1(n_2363),
.A2(n_1394),
.B1(n_1405),
.B2(n_1379),
.Y(n_2992)
);

INVx5_ASAP7_75t_L g2993 ( 
.A(n_2531),
.Y(n_2993)
);

INVx4_ASAP7_75t_L g2994 ( 
.A(n_2329),
.Y(n_2994)
);

INVx2_ASAP7_75t_SL g2995 ( 
.A(n_2562),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_SL g2996 ( 
.A(n_2431),
.B(n_1622),
.Y(n_2996)
);

AOI22xp5_ASAP7_75t_L g2997 ( 
.A1(n_2814),
.A2(n_2364),
.B1(n_2292),
.B2(n_2336),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2654),
.B(n_2585),
.Y(n_2998)
);

OAI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2942),
.A2(n_2252),
.B1(n_2259),
.B2(n_2389),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2684),
.B(n_2363),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2928),
.Y(n_3001)
);

AOI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2797),
.A2(n_2292),
.B1(n_2336),
.B2(n_2266),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2641),
.B(n_2343),
.Y(n_3003)
);

OR2x2_ASAP7_75t_L g3004 ( 
.A(n_2897),
.B(n_2419),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2667),
.A2(n_2341),
.B1(n_2350),
.B2(n_2345),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2638),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2704),
.B(n_2371),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2701),
.B(n_2371),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2638),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2644),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2850),
.B(n_2382),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2928),
.Y(n_3012)
);

OAI22xp33_ASAP7_75t_L g3013 ( 
.A1(n_2816),
.A2(n_2266),
.B1(n_2570),
.B2(n_2277),
.Y(n_3013)
);

O2A1O1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2643),
.A2(n_2630),
.B(n_2270),
.C(n_2483),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2717),
.B(n_2382),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2644),
.Y(n_3016)
);

OAI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2827),
.A2(n_2570),
.B1(n_2430),
.B2(n_2404),
.Y(n_3017)
);

A2O1A1Ixp33_ASAP7_75t_L g3018 ( 
.A1(n_2836),
.A2(n_2517),
.B(n_2354),
.C(n_2357),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2639),
.B(n_2433),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2839),
.B(n_2630),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2840),
.B(n_2307),
.Y(n_3021)
);

AOI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2674),
.A2(n_2477),
.B1(n_2431),
.B2(n_2460),
.Y(n_3022)
);

INVxp33_ASAP7_75t_SL g3023 ( 
.A(n_2757),
.Y(n_3023)
);

BUFx6f_ASAP7_75t_L g3024 ( 
.A(n_2815),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2967),
.A2(n_2358),
.B1(n_2365),
.B2(n_2352),
.Y(n_3025)
);

BUFx6f_ASAP7_75t_L g3026 ( 
.A(n_2815),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2645),
.Y(n_3027)
);

AOI22xp33_ASAP7_75t_L g3028 ( 
.A1(n_2884),
.A2(n_2375),
.B1(n_2386),
.B2(n_2366),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2780),
.B(n_2307),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2738),
.B(n_2433),
.Y(n_3030)
);

AOI22xp33_ASAP7_75t_L g3031 ( 
.A1(n_2935),
.A2(n_2391),
.B1(n_2394),
.B2(n_2390),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2990),
.B(n_2347),
.Y(n_3032)
);

AND2x4_ASAP7_75t_L g3033 ( 
.A(n_2653),
.B(n_2637),
.Y(n_3033)
);

NAND2x1p5_ASAP7_75t_L g3034 ( 
.A(n_2711),
.B(n_2766),
.Y(n_3034)
);

O2A1O1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2774),
.A2(n_2483),
.B(n_2460),
.C(n_2413),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2968),
.B(n_2435),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2653),
.B(n_2395),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2645),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2990),
.B(n_2416),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2990),
.B(n_2417),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_SL g3041 ( 
.A1(n_2761),
.A2(n_2600),
.B1(n_2430),
.B2(n_2404),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2635),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2915),
.B(n_2424),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2848),
.B(n_2305),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2927),
.B(n_2428),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2718),
.B(n_2432),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2646),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2730),
.B(n_2441),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2646),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2636),
.Y(n_3050)
);

BUFx6f_ASAP7_75t_SL g3051 ( 
.A(n_2888),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2772),
.B(n_2305),
.Y(n_3052)
);

INVx2_ASAP7_75t_SL g3053 ( 
.A(n_2665),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2694),
.B(n_2362),
.Y(n_3054)
);

NAND2x1p5_ASAP7_75t_L g3055 ( 
.A(n_2711),
.B(n_2398),
.Y(n_3055)
);

AO22x1_ASAP7_75t_L g3056 ( 
.A1(n_2723),
.A2(n_2235),
.B1(n_2176),
.B2(n_2362),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2649),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2891),
.B(n_2448),
.Y(n_3058)
);

NAND3xp33_ASAP7_75t_SL g3059 ( 
.A(n_2746),
.B(n_2534),
.C(n_2552),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2755),
.B(n_2455),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2760),
.B(n_2466),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2648),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2683),
.B(n_2720),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2688),
.A2(n_2477),
.B1(n_2502),
.B2(n_2488),
.Y(n_3064)
);

INVx4_ASAP7_75t_L g3065 ( 
.A(n_2767),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2944),
.B(n_2477),
.Y(n_3066)
);

HB1xp67_ASAP7_75t_L g3067 ( 
.A(n_2798),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2991),
.B(n_2477),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2750),
.B(n_2442),
.Y(n_3069)
);

OR2x6_ASAP7_75t_L g3070 ( 
.A(n_2652),
.B(n_2819),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2759),
.B(n_2477),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2648),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2988),
.B(n_2570),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2936),
.B(n_2434),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2669),
.B(n_2276),
.Y(n_3075)
);

NAND2xp33_ASAP7_75t_L g3076 ( 
.A(n_2657),
.B(n_2690),
.Y(n_3076)
);

NAND3xp33_ASAP7_75t_SL g3077 ( 
.A(n_2687),
.B(n_2534),
.C(n_2581),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2671),
.B(n_2600),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2656),
.Y(n_3079)
);

BUFx2_ASAP7_75t_L g3080 ( 
.A(n_2853),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_2666),
.B(n_2496),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2676),
.B(n_2600),
.Y(n_3082)
);

A2O1A1Ixp33_ASAP7_75t_SL g3083 ( 
.A1(n_2978),
.A2(n_2381),
.B(n_2377),
.C(n_2508),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2808),
.B(n_2288),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2756),
.B(n_2435),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2724),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2815),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2977),
.B(n_2488),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2751),
.B(n_2325),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2936),
.B(n_2310),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2656),
.B(n_2502),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2659),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2659),
.B(n_2498),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2660),
.B(n_2504),
.Y(n_3094)
);

BUFx12f_ASAP7_75t_L g3095 ( 
.A(n_2858),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_L g3096 ( 
.A1(n_2782),
.A2(n_2259),
.B1(n_2389),
.B2(n_2547),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2660),
.B(n_2504),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_2962),
.Y(n_3098)
);

INVx4_ASAP7_75t_L g3099 ( 
.A(n_2767),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2724),
.Y(n_3100)
);

AOI22xp33_ASAP7_75t_L g3101 ( 
.A1(n_2935),
.A2(n_2508),
.B1(n_2496),
.B2(n_2331),
.Y(n_3101)
);

CKINVDCx6p67_ASAP7_75t_R g3102 ( 
.A(n_2811),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2992),
.B(n_2509),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2992),
.B(n_2509),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_2936),
.B(n_2327),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_2855),
.B(n_2521),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2809),
.B(n_2771),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2789),
.A2(n_2331),
.B1(n_2340),
.B2(n_2284),
.Y(n_3108)
);

OR2x6_ASAP7_75t_L g3109 ( 
.A(n_2652),
.B(n_2430),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2703),
.B(n_2404),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2924),
.B(n_2883),
.Y(n_3111)
);

NOR2xp67_ASAP7_75t_L g3112 ( 
.A(n_2813),
.B(n_2609),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2771),
.B(n_2315),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2773),
.B(n_2315),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2779),
.B(n_2295),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_2637),
.B(n_2586),
.Y(n_3116)
);

NOR2x1p5_ASAP7_75t_L g3117 ( 
.A(n_2859),
.B(n_2611),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2773),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2962),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2785),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2785),
.Y(n_3121)
);

AOI22xp5_ASAP7_75t_L g3122 ( 
.A1(n_2903),
.A2(n_2419),
.B1(n_2540),
.B2(n_2527),
.Y(n_3122)
);

AND2x4_ASAP7_75t_L g3123 ( 
.A(n_2715),
.B(n_2351),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2791),
.B(n_2519),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2972),
.B(n_2553),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2661),
.A2(n_2329),
.B(n_2996),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2874),
.B(n_2568),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2791),
.B(n_2519),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2794),
.Y(n_3129)
);

AOI22xp5_ASAP7_75t_L g3130 ( 
.A1(n_2894),
.A2(n_2436),
.B1(n_2566),
.B2(n_2309),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2794),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2796),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_SL g3133 ( 
.A(n_2874),
.B(n_2309),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2796),
.B(n_2520),
.Y(n_3134)
);

OAI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2852),
.A2(n_2547),
.B(n_2470),
.Y(n_3135)
);

INVx4_ASAP7_75t_L g3136 ( 
.A(n_2767),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_2861),
.A2(n_2436),
.B1(n_2566),
.B2(n_2599),
.Y(n_3137)
);

AND2x6_ASAP7_75t_SL g3138 ( 
.A(n_2906),
.B(n_2176),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2810),
.Y(n_3139)
);

NAND2xp33_ASAP7_75t_L g3140 ( 
.A(n_2657),
.B(n_2329),
.Y(n_3140)
);

BUFx6f_ASAP7_75t_L g3141 ( 
.A(n_2841),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2810),
.B(n_2812),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2812),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2824),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2824),
.B(n_2520),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2712),
.B(n_2523),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2834),
.B(n_2838),
.Y(n_3147)
);

BUFx2_ASAP7_75t_L g3148 ( 
.A(n_2709),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2834),
.B(n_2523),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2838),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2898),
.Y(n_3151)
);

NOR3xp33_ASAP7_75t_L g3152 ( 
.A(n_2863),
.B(n_2300),
.C(n_2332),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2898),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2900),
.B(n_2532),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2789),
.A2(n_2340),
.B1(n_2284),
.B2(n_2476),
.Y(n_3155)
);

NAND2x1_ASAP7_75t_L g3156 ( 
.A(n_2657),
.B(n_2398),
.Y(n_3156)
);

INVx4_ASAP7_75t_L g3157 ( 
.A(n_2657),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2900),
.Y(n_3158)
);

NOR3xp33_ASAP7_75t_L g3159 ( 
.A(n_2847),
.B(n_2339),
.C(n_2332),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2736),
.B(n_2372),
.Y(n_3160)
);

NOR3xp33_ASAP7_75t_SL g3161 ( 
.A(n_2721),
.B(n_839),
.C(n_836),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_SL g3162 ( 
.A(n_2709),
.B(n_2450),
.Y(n_3162)
);

INVx4_ASAP7_75t_L g3163 ( 
.A(n_2690),
.Y(n_3163)
);

INVx3_ASAP7_75t_L g3164 ( 
.A(n_2690),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2902),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_SL g3166 ( 
.A(n_2679),
.B(n_2572),
.Y(n_3166)
);

AOI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_2686),
.A2(n_2599),
.B1(n_2476),
.B2(n_2339),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2825),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2902),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2904),
.B(n_2532),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2904),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2907),
.Y(n_3172)
);

O2A1O1Ixp33_ASAP7_75t_L g3173 ( 
.A1(n_2754),
.A2(n_1817),
.B(n_2536),
.C(n_2533),
.Y(n_3173)
);

AOI22xp33_ASAP7_75t_L g3174 ( 
.A1(n_2929),
.A2(n_2536),
.B1(n_2538),
.B2(n_2533),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2907),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2909),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2909),
.B(n_2538),
.Y(n_3177)
);

INVx2_ASAP7_75t_SL g3178 ( 
.A(n_2962),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_SL g3179 ( 
.A(n_2982),
.B(n_2572),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2753),
.B(n_2372),
.Y(n_3180)
);

O2A1O1Ixp33_ASAP7_75t_L g3181 ( 
.A1(n_2969),
.A2(n_2970),
.B(n_2943),
.C(n_2974),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2912),
.B(n_2551),
.Y(n_3182)
);

AND2x2_ASAP7_75t_L g3183 ( 
.A(n_2784),
.B(n_2599),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2912),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_2729),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_2929),
.A2(n_2580),
.B1(n_2592),
.B2(n_2578),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2917),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_SL g3188 ( 
.A(n_2982),
.B(n_2572),
.Y(n_3188)
);

AND2x4_ASAP7_75t_L g3189 ( 
.A(n_2715),
.B(n_2551),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2917),
.B(n_2554),
.Y(n_3190)
);

BUFx3_ASAP7_75t_L g3191 ( 
.A(n_2700),
.Y(n_3191)
);

INVx8_ASAP7_75t_L g3192 ( 
.A(n_2647),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2919),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2722),
.B(n_2554),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_2934),
.A2(n_2592),
.B1(n_2593),
.B2(n_2580),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_2726),
.B(n_2556),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2919),
.Y(n_3197)
);

NAND2xp33_ASAP7_75t_L g3198 ( 
.A(n_2702),
.B(n_2556),
.Y(n_3198)
);

BUFx3_ASAP7_75t_L g3199 ( 
.A(n_2849),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2923),
.Y(n_3200)
);

OAI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2803),
.A2(n_2469),
.B(n_2524),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2727),
.B(n_2728),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2934),
.A2(n_2603),
.B1(n_2567),
.B2(n_2569),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2732),
.B(n_2558),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_2737),
.B(n_2558),
.Y(n_3205)
);

AND2x2_ASAP7_75t_L g3206 ( 
.A(n_2770),
.B(n_1846),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_2864),
.B(n_1846),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2947),
.A2(n_2348),
.B(n_2333),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2854),
.A2(n_2348),
.B(n_2333),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2739),
.B(n_2567),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2740),
.B(n_2569),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_2923),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2948),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2742),
.B(n_2573),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_2819),
.Y(n_3215)
);

AOI22xp33_ASAP7_75t_L g3216 ( 
.A1(n_2940),
.A2(n_2574),
.B1(n_2576),
.B2(n_2573),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2948),
.B(n_2574),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_2946),
.B(n_2572),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2957),
.B(n_2601),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_2940),
.A2(n_2578),
.B1(n_2593),
.B2(n_2576),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2986),
.B(n_2604),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_2995),
.B(n_2235),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_2946),
.B(n_2577),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2949),
.Y(n_3224)
);

AOI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_2954),
.A2(n_2603),
.B1(n_2461),
.B2(n_2473),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2949),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2765),
.B(n_2235),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2860),
.B(n_1846),
.Y(n_3228)
);

INVx3_ASAP7_75t_L g3229 ( 
.A(n_2702),
.Y(n_3229)
);

BUFx6f_ASAP7_75t_L g3230 ( 
.A(n_2841),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2961),
.Y(n_3231)
);

OAI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_2971),
.A2(n_2499),
.B(n_2626),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_2954),
.A2(n_2461),
.B1(n_2473),
.B2(n_2471),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2961),
.Y(n_3234)
);

INVx4_ASAP7_75t_L g3235 ( 
.A(n_2702),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2788),
.A2(n_2471),
.B1(n_2514),
.B2(n_2503),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_2980),
.B(n_2878),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_2707),
.A2(n_2627),
.B1(n_2626),
.B2(n_2514),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_SL g3239 ( 
.A(n_2875),
.B(n_2577),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2964),
.Y(n_3240)
);

NOR2xp67_ASAP7_75t_L g3241 ( 
.A(n_2871),
.B(n_2627),
.Y(n_3241)
);

INVxp67_ASAP7_75t_L g3242 ( 
.A(n_2959),
.Y(n_3242)
);

BUFx2_ASAP7_75t_L g3243 ( 
.A(n_2913),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_2979),
.B(n_2503),
.Y(n_3244)
);

CKINVDCx5p33_ASAP7_75t_R g3245 ( 
.A(n_2634),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2959),
.B(n_1721),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2748),
.B(n_2565),
.Y(n_3247)
);

NOR2xp33_ASAP7_75t_L g3248 ( 
.A(n_2922),
.B(n_2565),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2964),
.Y(n_3249)
);

AOI22xp33_ASAP7_75t_L g3250 ( 
.A1(n_2788),
.A2(n_2584),
.B1(n_2632),
.B2(n_2618),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2989),
.B(n_2584),
.Y(n_3251)
);

NAND2xp33_ASAP7_75t_L g3252 ( 
.A(n_2731),
.B(n_2577),
.Y(n_3252)
);

OR2x2_ASAP7_75t_L g3253 ( 
.A(n_2879),
.B(n_1723),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2989),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2680),
.Y(n_3255)
);

NOR3xp33_ASAP7_75t_L g3256 ( 
.A(n_2938),
.B(n_1817),
.C(n_842),
.Y(n_3256)
);

OR2x2_ASAP7_75t_L g3257 ( 
.A(n_2807),
.B(n_1740),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2681),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_2658),
.B(n_2618),
.Y(n_3259)
);

CKINVDCx20_ASAP7_75t_R g3260 ( 
.A(n_2708),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_2685),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2778),
.B(n_2632),
.Y(n_3262)
);

AOI22xp5_ASAP7_75t_L g3263 ( 
.A1(n_2945),
.A2(n_2198),
.B1(n_838),
.B2(n_849),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_2790),
.A2(n_2342),
.B1(n_1056),
.B2(n_1817),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2693),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_2790),
.A2(n_2817),
.B1(n_2829),
.B2(n_2801),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2875),
.B(n_2577),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_2673),
.B(n_2560),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_2766),
.B(n_2560),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2689),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_2895),
.B(n_2472),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_2895),
.B(n_2472),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_2875),
.B(n_2480),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_L g3274 ( 
.A(n_2801),
.B(n_2480),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2781),
.B(n_2156),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_2817),
.A2(n_2342),
.B1(n_1661),
.B2(n_1746),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_2887),
.B(n_2529),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2699),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_L g3279 ( 
.A(n_2829),
.B(n_841),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2691),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2692),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2800),
.B(n_1661),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2802),
.B(n_1845),
.Y(n_3283)
);

OR2x6_ASAP7_75t_L g3284 ( 
.A(n_2905),
.B(n_1740),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2804),
.B(n_1845),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2805),
.B(n_2164),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_2887),
.B(n_2559),
.Y(n_3287)
);

AOI221xp5_ASAP7_75t_L g3288 ( 
.A1(n_2783),
.A2(n_853),
.B1(n_854),
.B2(n_847),
.C(n_843),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_2887),
.B(n_2529),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_SL g3290 ( 
.A(n_2731),
.B(n_2734),
.Y(n_3290)
);

A2O1A1Ixp33_ASAP7_75t_L g3291 ( 
.A1(n_2806),
.A2(n_2167),
.B(n_2173),
.C(n_2164),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_2696),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2698),
.B(n_2167),
.Y(n_3293)
);

NOR3xp33_ASAP7_75t_SL g3294 ( 
.A(n_2783),
.B(n_860),
.C(n_856),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2833),
.B(n_1746),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2706),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2818),
.B(n_2173),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_2705),
.Y(n_3298)
);

OR2x2_ASAP7_75t_L g3299 ( 
.A(n_2833),
.B(n_1756),
.Y(n_3299)
);

AOI21xp5_ASAP7_75t_L g3300 ( 
.A1(n_2963),
.A2(n_2544),
.B(n_2529),
.Y(n_3300)
);

INVx4_ASAP7_75t_L g3301 ( 
.A(n_2731),
.Y(n_3301)
);

NAND2xp33_ASAP7_75t_L g3302 ( 
.A(n_2734),
.B(n_2183),
.Y(n_3302)
);

AOI22xp5_ASAP7_75t_L g3303 ( 
.A1(n_2837),
.A2(n_868),
.B1(n_885),
.B2(n_819),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_2837),
.A2(n_2885),
.B1(n_2856),
.B2(n_2664),
.Y(n_3304)
);

AND2x6_ASAP7_75t_SL g3305 ( 
.A(n_2905),
.B(n_2953),
.Y(n_3305)
);

HB1xp67_ASAP7_75t_L g3306 ( 
.A(n_2856),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2862),
.Y(n_3307)
);

NOR3xp33_ASAP7_75t_L g3308 ( 
.A(n_2719),
.B(n_862),
.C(n_861),
.Y(n_3308)
);

AND2x6_ASAP7_75t_L g3309 ( 
.A(n_2734),
.B(n_2183),
.Y(n_3309)
);

AND2x4_ASAP7_75t_L g3310 ( 
.A(n_2786),
.B(n_1756),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_2885),
.B(n_1759),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_2662),
.A2(n_1760),
.B1(n_1779),
.B2(n_1759),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2777),
.B(n_1845),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2713),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2865),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2714),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2777),
.B(n_1845),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2866),
.Y(n_3318)
);

INVx2_ASAP7_75t_SL g3319 ( 
.A(n_2913),
.Y(n_3319)
);

NAND2xp33_ASAP7_75t_L g3320 ( 
.A(n_2743),
.B(n_2185),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2868),
.B(n_2185),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2873),
.B(n_2193),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2877),
.B(n_2193),
.Y(n_3323)
);

A2O1A1Ixp33_ASAP7_75t_SL g3324 ( 
.A1(n_2939),
.A2(n_2200),
.B(n_2203),
.C(n_2196),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2743),
.B(n_2529),
.Y(n_3325)
);

INVx2_ASAP7_75t_SL g3326 ( 
.A(n_2913),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2889),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3060),
.B(n_2640),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3020),
.B(n_2640),
.Y(n_3329)
);

HB1xp67_ASAP7_75t_L g3330 ( 
.A(n_3050),
.Y(n_3330)
);

OR2x2_ASAP7_75t_SL g3331 ( 
.A(n_3059),
.B(n_2921),
.Y(n_3331)
);

BUFx6f_ASAP7_75t_L g3332 ( 
.A(n_3024),
.Y(n_3332)
);

AND2x6_ASAP7_75t_SL g3333 ( 
.A(n_3237),
.B(n_2953),
.Y(n_3333)
);

INVx1_ASAP7_75t_SL g3334 ( 
.A(n_3080),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_3168),
.Y(n_3335)
);

AOI22xp5_ASAP7_75t_L g3336 ( 
.A1(n_2998),
.A2(n_2642),
.B1(n_2695),
.B2(n_2881),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_3067),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_2997),
.B(n_2921),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_SL g3339 ( 
.A(n_3002),
.B(n_2921),
.Y(n_3339)
);

INVx4_ASAP7_75t_L g3340 ( 
.A(n_3192),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_3021),
.B(n_2642),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3004),
.B(n_2695),
.Y(n_3342)
);

BUFx3_ASAP7_75t_L g3343 ( 
.A(n_3070),
.Y(n_3343)
);

AOI22x1_ASAP7_75t_L g3344 ( 
.A1(n_3208),
.A2(n_3232),
.B1(n_3118),
.B2(n_3120),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_3052),
.B(n_2811),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_3054),
.B(n_2811),
.Y(n_3346)
);

AND2x4_ASAP7_75t_SL g3347 ( 
.A(n_3070),
.B(n_2786),
.Y(n_3347)
);

OR2x6_ASAP7_75t_L g3348 ( 
.A(n_3070),
.B(n_2857),
.Y(n_3348)
);

INVx5_ASAP7_75t_L g3349 ( 
.A(n_3192),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3111),
.B(n_2933),
.Y(n_3350)
);

INVx2_ASAP7_75t_SL g3351 ( 
.A(n_3057),
.Y(n_3351)
);

AOI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3044),
.A2(n_2899),
.B1(n_2749),
.B2(n_2733),
.Y(n_3352)
);

INVx5_ASAP7_75t_L g3353 ( 
.A(n_3192),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3043),
.B(n_2733),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3053),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3079),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3092),
.Y(n_3357)
);

INVx3_ASAP7_75t_L g3358 ( 
.A(n_3157),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_3033),
.B(n_2708),
.Y(n_3359)
);

BUFx2_ASAP7_75t_L g3360 ( 
.A(n_3148),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_3023),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3045),
.B(n_2749),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3202),
.Y(n_3363)
);

INVx5_ASAP7_75t_L g3364 ( 
.A(n_3157),
.Y(n_3364)
);

INVx2_ASAP7_75t_SL g3365 ( 
.A(n_3191),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_SL g3366 ( 
.A1(n_3041),
.A2(n_2857),
.B1(n_2822),
.B2(n_2831),
.Y(n_3366)
);

CKINVDCx20_ASAP7_75t_R g3367 ( 
.A(n_3245),
.Y(n_3367)
);

AO21x2_ASAP7_75t_L g3368 ( 
.A1(n_3135),
.A2(n_2951),
.B(n_2763),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3255),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3258),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3270),
.Y(n_3371)
);

AOI22xp5_ASAP7_75t_L g3372 ( 
.A1(n_3013),
.A2(n_2650),
.B1(n_2831),
.B2(n_2822),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_3033),
.B(n_2933),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_3061),
.B(n_2886),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3280),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3086),
.Y(n_3376)
);

BUFx4f_ASAP7_75t_L g3377 ( 
.A(n_3095),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3132),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3046),
.B(n_2892),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_3269),
.Y(n_3380)
);

BUFx12f_ASAP7_75t_L g3381 ( 
.A(n_3305),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_3269),
.Y(n_3382)
);

INVx1_ASAP7_75t_SL g3383 ( 
.A(n_3199),
.Y(n_3383)
);

BUFx12f_ASAP7_75t_L g3384 ( 
.A(n_3243),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_L g3385 ( 
.A1(n_3259),
.A2(n_2775),
.B(n_2752),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3281),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3292),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_3215),
.Y(n_3388)
);

O2A1O1Ixp5_ASAP7_75t_L g3389 ( 
.A1(n_3106),
.A2(n_2911),
.B(n_2744),
.C(n_2793),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_3150),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3048),
.B(n_2965),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3296),
.Y(n_3392)
);

BUFx3_ASAP7_75t_L g3393 ( 
.A(n_3185),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_3151),
.Y(n_3394)
);

INVx2_ASAP7_75t_L g3395 ( 
.A(n_3158),
.Y(n_3395)
);

INVx5_ASAP7_75t_L g3396 ( 
.A(n_3309),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3000),
.B(n_3058),
.Y(n_3397)
);

INVx2_ASAP7_75t_SL g3398 ( 
.A(n_3319),
.Y(n_3398)
);

AOI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3122),
.A2(n_2650),
.B1(n_2985),
.B2(n_2981),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3307),
.Y(n_3400)
);

HB1xp67_ASAP7_75t_L g3401 ( 
.A(n_3306),
.Y(n_3401)
);

INVx4_ASAP7_75t_L g3402 ( 
.A(n_3065),
.Y(n_3402)
);

INVxp67_ASAP7_75t_L g3403 ( 
.A(n_3081),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3315),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3318),
.Y(n_3405)
);

INVx2_ASAP7_75t_SL g3406 ( 
.A(n_3326),
.Y(n_3406)
);

HB1xp67_ASAP7_75t_L g3407 ( 
.A(n_3242),
.Y(n_3407)
);

AND2x4_ASAP7_75t_L g3408 ( 
.A(n_3037),
.B(n_2933),
.Y(n_3408)
);

INVx5_ASAP7_75t_L g3409 ( 
.A(n_3309),
.Y(n_3409)
);

INVx2_ASAP7_75t_SL g3410 ( 
.A(n_3098),
.Y(n_3410)
);

BUFx2_ASAP7_75t_L g3411 ( 
.A(n_3037),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3327),
.Y(n_3412)
);

AOI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3110),
.A2(n_2795),
.B1(n_2993),
.B2(n_2668),
.Y(n_3413)
);

CKINVDCx5p33_ASAP7_75t_R g3414 ( 
.A(n_3051),
.Y(n_3414)
);

INVx4_ASAP7_75t_L g3415 ( 
.A(n_3065),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3165),
.Y(n_3416)
);

BUFx8_ASAP7_75t_L g3417 ( 
.A(n_3051),
.Y(n_3417)
);

INVx1_ASAP7_75t_SL g3418 ( 
.A(n_3119),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3100),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3121),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3295),
.B(n_2993),
.Y(n_3421)
);

INVx5_ASAP7_75t_L g3422 ( 
.A(n_3309),
.Y(n_3422)
);

INVx2_ASAP7_75t_SL g3423 ( 
.A(n_3178),
.Y(n_3423)
);

AOI22xp33_ASAP7_75t_L g3424 ( 
.A1(n_3029),
.A2(n_2670),
.B1(n_2682),
.B2(n_2672),
.Y(n_3424)
);

HB1xp67_ASAP7_75t_L g3425 ( 
.A(n_3189),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_3248),
.B(n_2993),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_3071),
.B(n_2633),
.Y(n_3427)
);

INVx6_ASAP7_75t_L g3428 ( 
.A(n_3117),
.Y(n_3428)
);

INVx4_ASAP7_75t_L g3429 ( 
.A(n_3099),
.Y(n_3429)
);

HB1xp67_ASAP7_75t_L g3430 ( 
.A(n_3189),
.Y(n_3430)
);

AND2x4_ASAP7_75t_L g3431 ( 
.A(n_3123),
.B(n_2677),
.Y(n_3431)
);

BUFx4f_ASAP7_75t_L g3432 ( 
.A(n_3102),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3219),
.B(n_2633),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3129),
.Y(n_3434)
);

CKINVDCx5p33_ASAP7_75t_R g3435 ( 
.A(n_3260),
.Y(n_3435)
);

NAND3xp33_ASAP7_75t_L g3436 ( 
.A(n_3288),
.B(n_2890),
.C(n_2867),
.Y(n_3436)
);

CKINVDCx20_ASAP7_75t_R g3437 ( 
.A(n_3161),
.Y(n_3437)
);

BUFx6f_ASAP7_75t_L g3438 ( 
.A(n_3024),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3131),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3206),
.Y(n_3440)
);

CKINVDCx5p33_ASAP7_75t_R g3441 ( 
.A(n_3138),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3034),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_SL g3443 ( 
.A(n_3266),
.B(n_2743),
.Y(n_3443)
);

INVx2_ASAP7_75t_SL g3444 ( 
.A(n_3123),
.Y(n_3444)
);

OR2x6_ASAP7_75t_L g3445 ( 
.A(n_3109),
.B(n_2663),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3221),
.B(n_2762),
.Y(n_3446)
);

A2O1A1Ixp33_ASAP7_75t_L g3447 ( 
.A1(n_3014),
.A2(n_2675),
.B(n_2910),
.C(n_2893),
.Y(n_3447)
);

OR2x2_ASAP7_75t_L g3448 ( 
.A(n_3299),
.B(n_3253),
.Y(n_3448)
);

INVx3_ASAP7_75t_L g3449 ( 
.A(n_3034),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3169),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3019),
.B(n_2762),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3019),
.B(n_2762),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3171),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_3073),
.B(n_2677),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3139),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3143),
.Y(n_3456)
);

INVx2_ASAP7_75t_SL g3457 ( 
.A(n_3116),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3077),
.B(n_2735),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3144),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3311),
.B(n_3107),
.Y(n_3460)
);

BUFx2_ASAP7_75t_L g3461 ( 
.A(n_3228),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_3246),
.Y(n_3462)
);

BUFx2_ASAP7_75t_L g3463 ( 
.A(n_3183),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3163),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3153),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3172),
.Y(n_3466)
);

AOI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3256),
.A2(n_2821),
.B1(n_2776),
.B2(n_2769),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3107),
.B(n_2741),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3175),
.Y(n_3469)
);

AND2x4_ASAP7_75t_L g3470 ( 
.A(n_3116),
.B(n_2663),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3304),
.B(n_2745),
.Y(n_3471)
);

NAND2x1p5_ASAP7_75t_L g3472 ( 
.A(n_3099),
.B(n_2901),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3187),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3028),
.B(n_3025),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3279),
.B(n_2747),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3088),
.B(n_2758),
.Y(n_3476)
);

BUFx2_ASAP7_75t_L g3477 ( 
.A(n_3164),
.Y(n_3477)
);

INVx5_ASAP7_75t_L g3478 ( 
.A(n_3309),
.Y(n_3478)
);

OR2x2_ASAP7_75t_SL g3479 ( 
.A(n_3257),
.B(n_2663),
.Y(n_3479)
);

BUFx2_ASAP7_75t_L g3480 ( 
.A(n_3164),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3207),
.B(n_2764),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3193),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3176),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3200),
.Y(n_3484)
);

BUFx12f_ASAP7_75t_L g3485 ( 
.A(n_3284),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3184),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3005),
.B(n_2768),
.Y(n_3487)
);

OAI22xp5_ASAP7_75t_SL g3488 ( 
.A1(n_3109),
.A2(n_866),
.B1(n_867),
.B2(n_863),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3213),
.Y(n_3489)
);

BUFx6f_ASAP7_75t_L g3490 ( 
.A(n_3024),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3224),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_3109),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3226),
.Y(n_3493)
);

INVx2_ASAP7_75t_SL g3494 ( 
.A(n_3089),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3006),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3009),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3010),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3016),
.Y(n_3498)
);

BUFx12f_ASAP7_75t_L g3499 ( 
.A(n_3284),
.Y(n_3499)
);

INVx2_ASAP7_75t_SL g3500 ( 
.A(n_3284),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3027),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3075),
.B(n_2787),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3031),
.B(n_2792),
.Y(n_3503)
);

INVx5_ASAP7_75t_L g3504 ( 
.A(n_3026),
.Y(n_3504)
);

OR2x4_ASAP7_75t_L g3505 ( 
.A(n_3222),
.B(n_2678),
.Y(n_3505)
);

CKINVDCx5p33_ASAP7_75t_R g3506 ( 
.A(n_3115),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3003),
.B(n_2799),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3003),
.B(n_2823),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3136),
.B(n_2678),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3038),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3047),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3085),
.B(n_2826),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_3163),
.Y(n_3513)
);

BUFx3_ASAP7_75t_L g3514 ( 
.A(n_3160),
.Y(n_3514)
);

AOI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_3084),
.A2(n_3166),
.B1(n_3112),
.B2(n_3137),
.Y(n_3515)
);

INVx3_ASAP7_75t_L g3516 ( 
.A(n_3235),
.Y(n_3516)
);

BUFx8_ASAP7_75t_L g3517 ( 
.A(n_3026),
.Y(n_3517)
);

BUFx6f_ASAP7_75t_L g3518 ( 
.A(n_3026),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3197),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3212),
.Y(n_3520)
);

INVx5_ASAP7_75t_L g3521 ( 
.A(n_3087),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_3017),
.B(n_2678),
.Y(n_3522)
);

INVx2_ASAP7_75t_SL g3523 ( 
.A(n_3063),
.Y(n_3523)
);

BUFx6f_ASAP7_75t_L g3524 ( 
.A(n_3087),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3231),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3180),
.A2(n_2821),
.B1(n_2725),
.B2(n_2716),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_3056),
.Y(n_3527)
);

BUFx2_ASAP7_75t_L g3528 ( 
.A(n_3229),
.Y(n_3528)
);

NOR2xp33_ASAP7_75t_R g3529 ( 
.A(n_3136),
.B(n_3076),
.Y(n_3529)
);

OR2x2_ASAP7_75t_L g3530 ( 
.A(n_3078),
.B(n_2828),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3008),
.B(n_2832),
.Y(n_3531)
);

INVxp67_ASAP7_75t_SL g3532 ( 
.A(n_2999),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3234),
.Y(n_3533)
);

INVx1_ASAP7_75t_SL g3534 ( 
.A(n_3082),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3064),
.B(n_3238),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3240),
.Y(n_3536)
);

OAI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3130),
.A2(n_2775),
.B1(n_2752),
.B2(n_2901),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3249),
.Y(n_3538)
);

AND2x2_ASAP7_75t_L g3539 ( 
.A(n_3294),
.B(n_2845),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3254),
.Y(n_3540)
);

AND2x2_ASAP7_75t_SL g3541 ( 
.A(n_3108),
.B(n_2941),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_3229),
.Y(n_3542)
);

AOI22xp5_ASAP7_75t_L g3543 ( 
.A1(n_3133),
.A2(n_2821),
.B1(n_2655),
.B2(n_2697),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3008),
.B(n_2880),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3066),
.B(n_2882),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3274),
.B(n_2914),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_L g3547 ( 
.A1(n_3068),
.A2(n_2821),
.B1(n_2651),
.B2(n_2896),
.Y(n_3547)
);

BUFx3_ASAP7_75t_L g3548 ( 
.A(n_3087),
.Y(n_3548)
);

OR2x6_ASAP7_75t_L g3549 ( 
.A(n_3032),
.B(n_2941),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3036),
.B(n_2918),
.Y(n_3550)
);

AND2x6_ASAP7_75t_L g3551 ( 
.A(n_3022),
.B(n_2841),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3238),
.B(n_2851),
.Y(n_3552)
);

INVxp67_ASAP7_75t_L g3553 ( 
.A(n_3227),
.Y(n_3553)
);

OAI21xp5_ASAP7_75t_L g3554 ( 
.A1(n_3018),
.A2(n_2926),
.B(n_2925),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3235),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3142),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3049),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3062),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3072),
.Y(n_3559)
);

OR2x6_ASAP7_75t_L g3560 ( 
.A(n_3241),
.B(n_2955),
.Y(n_3560)
);

AND2x4_ASAP7_75t_SL g3561 ( 
.A(n_3301),
.B(n_2851),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3036),
.B(n_3091),
.Y(n_3562)
);

BUFx3_ASAP7_75t_L g3563 ( 
.A(n_3141),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_3537),
.A2(n_2999),
.B(n_3096),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3397),
.B(n_3069),
.Y(n_3565)
);

OAI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_3328),
.A2(n_3167),
.B1(n_3101),
.B2(n_3155),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3460),
.B(n_3162),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_3376),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3338),
.A2(n_3083),
.B(n_3308),
.C(n_3035),
.Y(n_3569)
);

AND2x2_ASAP7_75t_L g3570 ( 
.A(n_3462),
.B(n_3042),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3374),
.A2(n_3096),
.B(n_3259),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3363),
.B(n_3379),
.Y(n_3572)
);

AOI21xp33_ASAP7_75t_L g3573 ( 
.A1(n_3474),
.A2(n_3436),
.B(n_3181),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_3504),
.Y(n_3574)
);

OAI22x1_ASAP7_75t_L g3575 ( 
.A1(n_3515),
.A2(n_3372),
.B1(n_3413),
.B2(n_3339),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3356),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_3378),
.Y(n_3577)
);

AND2x4_ASAP7_75t_L g3578 ( 
.A(n_3431),
.B(n_3310),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_3504),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_L g3580 ( 
.A1(n_3385),
.A2(n_3135),
.B(n_3535),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3391),
.B(n_3125),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3329),
.B(n_3244),
.Y(n_3582)
);

BUFx3_ASAP7_75t_L g3583 ( 
.A(n_3384),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_3330),
.Y(n_3584)
);

A2O1A1Ixp33_ASAP7_75t_L g3585 ( 
.A1(n_3447),
.A2(n_3152),
.B(n_3159),
.C(n_3263),
.Y(n_3585)
);

AOI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3539),
.A2(n_3127),
.B1(n_3040),
.B2(n_3039),
.Y(n_3586)
);

OAI21xp33_ASAP7_75t_L g3587 ( 
.A1(n_3354),
.A2(n_3362),
.B(n_3475),
.Y(n_3587)
);

O2A1O1Ixp5_ASAP7_75t_L g3588 ( 
.A1(n_3522),
.A2(n_3426),
.B(n_3458),
.C(n_3552),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3390),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3541),
.A2(n_3126),
.B(n_3140),
.Y(n_3590)
);

OAI22xp5_ASAP7_75t_SL g3591 ( 
.A1(n_3366),
.A2(n_3506),
.B1(n_3488),
.B2(n_3331),
.Y(n_3591)
);

A2O1A1Ixp33_ASAP7_75t_L g3592 ( 
.A1(n_3341),
.A2(n_3268),
.B(n_3173),
.C(n_3103),
.Y(n_3592)
);

HB1xp67_ASAP7_75t_L g3593 ( 
.A(n_3337),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3554),
.A2(n_3007),
.B(n_3015),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3440),
.B(n_3463),
.Y(n_3595)
);

O2A1O1Ixp5_ASAP7_75t_L g3596 ( 
.A1(n_3389),
.A2(n_3074),
.B(n_3105),
.C(n_3090),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3562),
.A2(n_3007),
.B(n_3015),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3448),
.B(n_3303),
.Y(n_3598)
);

O2A1O1Ixp33_ASAP7_75t_L g3599 ( 
.A1(n_3553),
.A2(n_3324),
.B(n_3104),
.C(n_3223),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3556),
.A2(n_3030),
.B(n_3198),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3534),
.B(n_3261),
.Y(n_3601)
);

OAI22xp5_ASAP7_75t_L g3602 ( 
.A1(n_3479),
.A2(n_3233),
.B1(n_3250),
.B2(n_3236),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3394),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3345),
.B(n_3310),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3357),
.Y(n_3605)
);

O2A1O1Ixp33_ASAP7_75t_L g3606 ( 
.A1(n_3403),
.A2(n_3218),
.B(n_3188),
.C(n_3179),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3342),
.B(n_3334),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3556),
.A2(n_3030),
.B(n_3300),
.Y(n_3608)
);

OAI22xp5_ASAP7_75t_L g3609 ( 
.A1(n_3352),
.A2(n_3225),
.B1(n_3272),
.B2(n_3271),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3419),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_3401),
.B(n_3265),
.Y(n_3611)
);

AOI22xp5_ASAP7_75t_L g3612 ( 
.A1(n_3350),
.A2(n_3273),
.B1(n_3317),
.B2(n_3313),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3468),
.A2(n_3252),
.B(n_3011),
.Y(n_3613)
);

OAI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3545),
.A2(n_3285),
.B(n_3283),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_L g3615 ( 
.A(n_3504),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3532),
.A2(n_3298),
.B1(n_3314),
.B2(n_3278),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_3396),
.A2(n_3011),
.B(n_3232),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3425),
.B(n_3316),
.Y(n_3618)
);

BUFx6f_ASAP7_75t_L g3619 ( 
.A(n_3521),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3396),
.A2(n_3114),
.B(n_3113),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3420),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3434),
.Y(n_3622)
);

OAI21xp33_ASAP7_75t_SL g3623 ( 
.A1(n_3543),
.A2(n_3147),
.B(n_3142),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3430),
.B(n_3001),
.Y(n_3624)
);

BUFx2_ASAP7_75t_L g3625 ( 
.A(n_3411),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3396),
.A2(n_3114),
.B(n_3113),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3461),
.B(n_3346),
.Y(n_3627)
);

O2A1O1Ixp33_ASAP7_75t_L g3628 ( 
.A1(n_3443),
.A2(n_3267),
.B(n_3239),
.C(n_1375),
.Y(n_3628)
);

NOR2xp33_ASAP7_75t_L g3629 ( 
.A(n_3454),
.B(n_3012),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3395),
.Y(n_3630)
);

NOR2xp33_ASAP7_75t_L g3631 ( 
.A(n_3514),
.B(n_3277),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_3336),
.B(n_3262),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_SL g3633 ( 
.A(n_3523),
.B(n_3262),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3409),
.A2(n_3201),
.B(n_3276),
.Y(n_3634)
);

AOI21xp5_ASAP7_75t_L g3635 ( 
.A1(n_3409),
.A2(n_3201),
.B(n_3209),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3344),
.A2(n_3297),
.B(n_3293),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3416),
.Y(n_3637)
);

NAND2x1p5_ASAP7_75t_L g3638 ( 
.A(n_3349),
.B(n_3301),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3409),
.A2(n_3156),
.B(n_3147),
.Y(n_3639)
);

HB1xp67_ASAP7_75t_L g3640 ( 
.A(n_3355),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3450),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3381),
.A2(n_3499),
.B1(n_3485),
.B2(n_3407),
.Y(n_3642)
);

BUFx6f_ASAP7_75t_L g3643 ( 
.A(n_3521),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3439),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3422),
.A2(n_3320),
.B(n_3302),
.Y(n_3645)
);

NOR2xp33_ASAP7_75t_L g3646 ( 
.A(n_3361),
.B(n_3287),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3455),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_3453),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3456),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3459),
.Y(n_3650)
);

BUFx6f_ASAP7_75t_L g3651 ( 
.A(n_3521),
.Y(n_3651)
);

O2A1O1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_3500),
.A2(n_1376),
.B(n_1381),
.C(n_1374),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3343),
.Y(n_3653)
);

BUFx6f_ASAP7_75t_L g3654 ( 
.A(n_3332),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3483),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_3422),
.A2(n_3128),
.B(n_3124),
.Y(n_3656)
);

NOR2xp67_ASAP7_75t_L g3657 ( 
.A(n_3335),
.B(n_3289),
.Y(n_3657)
);

A2O1A1Ixp33_ASAP7_75t_L g3658 ( 
.A1(n_3427),
.A2(n_3247),
.B(n_3264),
.C(n_3194),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3486),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_3332),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_SL g3661 ( 
.A(n_3399),
.B(n_3093),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3422),
.A2(n_3128),
.B(n_3124),
.Y(n_3662)
);

HB1xp67_ASAP7_75t_L g3663 ( 
.A(n_3360),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_SL g3664 ( 
.A(n_3446),
.B(n_3094),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3465),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3519),
.Y(n_3666)
);

NAND2x1p5_ASAP7_75t_L g3667 ( 
.A(n_3349),
.B(n_3141),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3502),
.B(n_3146),
.Y(n_3668)
);

A2O1A1Ixp33_ASAP7_75t_L g3669 ( 
.A1(n_3467),
.A2(n_3196),
.B(n_3205),
.C(n_3204),
.Y(n_3669)
);

NOR2xp33_ASAP7_75t_L g3670 ( 
.A(n_3383),
.B(n_3141),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_3364),
.Y(n_3671)
);

OAI22xp5_ASAP7_75t_L g3672 ( 
.A1(n_3505),
.A2(n_3174),
.B1(n_3195),
.B2(n_3186),
.Y(n_3672)
);

AO21x1_ASAP7_75t_L g3673 ( 
.A1(n_3487),
.A2(n_3290),
.B(n_3097),
.Y(n_3673)
);

O2A1O1Ixp5_ASAP7_75t_L g3674 ( 
.A1(n_3433),
.A2(n_3325),
.B(n_3546),
.C(n_3471),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3421),
.B(n_3210),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3476),
.B(n_3494),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3466),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3536),
.Y(n_3678)
);

NOR2xp67_ASAP7_75t_L g3679 ( 
.A(n_3388),
.B(n_3282),
.Y(n_3679)
);

BUFx5_ASAP7_75t_L g3680 ( 
.A(n_3551),
.Y(n_3680)
);

BUFx6f_ASAP7_75t_L g3681 ( 
.A(n_3332),
.Y(n_3681)
);

AND2x4_ASAP7_75t_L g3682 ( 
.A(n_3431),
.B(n_3470),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_SL g3683 ( 
.A(n_3481),
.B(n_3527),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_3492),
.A2(n_3216),
.B1(n_3220),
.B2(n_3203),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_L g3685 ( 
.A1(n_3478),
.A2(n_3145),
.B(n_3134),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_3367),
.B(n_3230),
.Y(n_3686)
);

O2A1O1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3369),
.A2(n_1384),
.B(n_1388),
.C(n_1383),
.Y(n_3687)
);

A2O1A1Ixp33_ASAP7_75t_L g3688 ( 
.A1(n_3526),
.A2(n_3214),
.B(n_3211),
.C(n_3312),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3478),
.A2(n_3145),
.B(n_3134),
.Y(n_3689)
);

A2O1A1Ixp33_ASAP7_75t_L g3690 ( 
.A1(n_3503),
.A2(n_3275),
.B(n_3286),
.C(n_3251),
.Y(n_3690)
);

A2O1A1Ixp33_ASAP7_75t_L g3691 ( 
.A1(n_3547),
.A2(n_3275),
.B(n_3286),
.C(n_3251),
.Y(n_3691)
);

OAI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_3445),
.A2(n_2994),
.B1(n_2955),
.B2(n_3055),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3469),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3478),
.A2(n_3154),
.B(n_3149),
.Y(n_3694)
);

BUFx6f_ASAP7_75t_L g3695 ( 
.A(n_3438),
.Y(n_3695)
);

HB1xp67_ASAP7_75t_L g3696 ( 
.A(n_3418),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3351),
.B(n_3230),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3473),
.Y(n_3698)
);

INVx4_ASAP7_75t_L g3699 ( 
.A(n_3349),
.Y(n_3699)
);

INVx4_ASAP7_75t_L g3700 ( 
.A(n_3353),
.Y(n_3700)
);

HB1xp67_ASAP7_75t_L g3701 ( 
.A(n_3393),
.Y(n_3701)
);

BUFx2_ASAP7_75t_L g3702 ( 
.A(n_3517),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3530),
.B(n_3149),
.Y(n_3703)
);

AOI22xp33_ASAP7_75t_L g3704 ( 
.A1(n_3551),
.A2(n_792),
.B1(n_827),
.B2(n_767),
.Y(n_3704)
);

A2O1A1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3370),
.A2(n_3291),
.B(n_3170),
.C(n_3177),
.Y(n_3705)
);

A2O1A1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_3371),
.A2(n_3170),
.B(n_3177),
.C(n_3154),
.Y(n_3706)
);

BUFx12f_ASAP7_75t_L g3707 ( 
.A(n_3417),
.Y(n_3707)
);

AND2x4_ASAP7_75t_L g3708 ( 
.A(n_3470),
.B(n_3230),
.Y(n_3708)
);

BUFx6f_ASAP7_75t_L g3709 ( 
.A(n_3438),
.Y(n_3709)
);

INVx1_ASAP7_75t_SL g3710 ( 
.A(n_3365),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3512),
.B(n_3182),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3408),
.B(n_3550),
.Y(n_3712)
);

BUFx3_ASAP7_75t_L g3713 ( 
.A(n_3517),
.Y(n_3713)
);

AOI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3507),
.A2(n_3190),
.B(n_3182),
.Y(n_3714)
);

NAND3xp33_ASAP7_75t_SL g3715 ( 
.A(n_3437),
.B(n_877),
.C(n_869),
.Y(n_3715)
);

O2A1O1Ixp33_ASAP7_75t_L g3716 ( 
.A1(n_3375),
.A2(n_1391),
.B(n_1395),
.C(n_1392),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3408),
.B(n_3190),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3445),
.A2(n_2994),
.B1(n_3055),
.B2(n_3217),
.Y(n_3718)
);

A2O1A1Ixp33_ASAP7_75t_L g3719 ( 
.A1(n_3386),
.A2(n_3217),
.B(n_2930),
.C(n_2937),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3540),
.B(n_3444),
.Y(n_3720)
);

INVxp67_ASAP7_75t_L g3721 ( 
.A(n_3398),
.Y(n_3721)
);

AOI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3508),
.A2(n_3297),
.B(n_3293),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3424),
.A2(n_2830),
.B1(n_2820),
.B2(n_2851),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3482),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3344),
.A2(n_3322),
.B(n_3321),
.Y(n_3725)
);

O2A1O1Ixp5_ASAP7_75t_L g3726 ( 
.A1(n_3451),
.A2(n_3321),
.B(n_3323),
.C(n_3322),
.Y(n_3726)
);

O2A1O1Ixp5_ASAP7_75t_L g3727 ( 
.A1(n_3452),
.A2(n_3323),
.B(n_2911),
.C(n_2950),
.Y(n_3727)
);

NAND3xp33_ASAP7_75t_L g3728 ( 
.A(n_3417),
.B(n_878),
.C(n_875),
.Y(n_3728)
);

NOR3xp33_ASAP7_75t_L g3729 ( 
.A(n_3457),
.B(n_1399),
.C(n_1396),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3368),
.A2(n_2830),
.B(n_2820),
.Y(n_3730)
);

A2O1A1Ixp33_ASAP7_75t_L g3731 ( 
.A1(n_3387),
.A2(n_2952),
.B(n_2958),
.C(n_2932),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_L g3732 ( 
.A(n_3435),
.B(n_3373),
.Y(n_3732)
);

AOI21xp5_ASAP7_75t_L g3733 ( 
.A1(n_3531),
.A2(n_2870),
.B(n_2869),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3392),
.B(n_2920),
.Y(n_3734)
);

AND2x4_ASAP7_75t_L g3735 ( 
.A(n_3373),
.B(n_2835),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3484),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3544),
.A2(n_2966),
.B(n_2960),
.Y(n_3737)
);

NOR2xp33_ASAP7_75t_L g3738 ( 
.A(n_3333),
.B(n_3428),
.Y(n_3738)
);

INVx3_ASAP7_75t_L g3739 ( 
.A(n_3364),
.Y(n_3739)
);

AOI21x1_ASAP7_75t_L g3740 ( 
.A1(n_3489),
.A2(n_2976),
.B(n_2975),
.Y(n_3740)
);

BUFx6f_ASAP7_75t_L g3741 ( 
.A(n_3438),
.Y(n_3741)
);

A2O1A1Ixp33_ASAP7_75t_L g3742 ( 
.A1(n_3400),
.A2(n_2984),
.B(n_2956),
.C(n_2973),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3364),
.A2(n_2870),
.B(n_2869),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3491),
.Y(n_3744)
);

BUFx2_ASAP7_75t_L g3745 ( 
.A(n_3548),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3560),
.A2(n_2870),
.B(n_2869),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3404),
.B(n_3405),
.Y(n_3747)
);

A2O1A1Ixp33_ASAP7_75t_L g3748 ( 
.A1(n_3412),
.A2(n_2983),
.B(n_2987),
.C(n_2931),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3551),
.A2(n_792),
.B1(n_827),
.B2(n_767),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3520),
.B(n_1760),
.Y(n_3750)
);

NOR2x1_ASAP7_75t_SL g3751 ( 
.A(n_3560),
.B(n_2872),
.Y(n_3751)
);

AOI21x1_ASAP7_75t_L g3752 ( 
.A1(n_3493),
.A2(n_2200),
.B(n_2196),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3428),
.B(n_3410),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3495),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3525),
.B(n_1779),
.Y(n_3755)
);

O2A1O1Ixp33_ASAP7_75t_L g3756 ( 
.A1(n_3348),
.A2(n_1400),
.B(n_1402),
.C(n_1401),
.Y(n_3756)
);

INVx2_ASAP7_75t_SL g3757 ( 
.A(n_3432),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3496),
.Y(n_3758)
);

INVx3_ASAP7_75t_L g3759 ( 
.A(n_3340),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3533),
.B(n_3538),
.Y(n_3760)
);

INVxp67_ASAP7_75t_SL g3761 ( 
.A(n_3557),
.Y(n_3761)
);

OR2x2_ASAP7_75t_L g3762 ( 
.A(n_3558),
.B(n_1522),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_L g3763 ( 
.A1(n_3549),
.A2(n_2872),
.B(n_2559),
.Y(n_3763)
);

O2A1O1Ixp33_ASAP7_75t_L g3764 ( 
.A1(n_3348),
.A2(n_1404),
.B(n_1407),
.C(n_1406),
.Y(n_3764)
);

A2O1A1Ixp33_ASAP7_75t_SL g3765 ( 
.A1(n_3358),
.A2(n_2843),
.B(n_2846),
.C(n_2835),
.Y(n_3765)
);

CKINVDCx5p33_ASAP7_75t_R g3766 ( 
.A(n_3377),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3340),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3353),
.A2(n_2872),
.B1(n_2846),
.B2(n_2843),
.Y(n_3768)
);

A2O1A1Ixp33_ASAP7_75t_SL g3769 ( 
.A1(n_3358),
.A2(n_1783),
.B(n_1784),
.C(n_1781),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3497),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3559),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_3377),
.Y(n_3772)
);

BUFx2_ASAP7_75t_L g3773 ( 
.A(n_3563),
.Y(n_3773)
);

AOI21xp5_ASAP7_75t_L g3774 ( 
.A1(n_3549),
.A2(n_2559),
.B(n_2544),
.Y(n_3774)
);

INVx1_ASAP7_75t_SL g3775 ( 
.A(n_3423),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3498),
.B(n_1781),
.Y(n_3776)
);

OAI21xp33_ASAP7_75t_L g3777 ( 
.A1(n_3501),
.A2(n_884),
.B(n_880),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3380),
.B(n_3382),
.Y(n_3778)
);

OAI22xp5_ASAP7_75t_L g3779 ( 
.A1(n_3353),
.A2(n_894),
.B1(n_895),
.B2(n_886),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3359),
.B(n_1408),
.Y(n_3780)
);

A2O1A1Ixp33_ASAP7_75t_SL g3781 ( 
.A1(n_3442),
.A2(n_1784),
.B(n_1801),
.C(n_1783),
.Y(n_3781)
);

O2A1O1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_3510),
.A2(n_1413),
.B(n_1416),
.C(n_1414),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3380),
.B(n_887),
.Y(n_3783)
);

OAI21xp5_ASAP7_75t_L g3784 ( 
.A1(n_3551),
.A2(n_2655),
.B(n_2647),
.Y(n_3784)
);

OR2x2_ASAP7_75t_L g3785 ( 
.A(n_3511),
.B(n_3477),
.Y(n_3785)
);

BUFx2_ASAP7_75t_L g3786 ( 
.A(n_3480),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3382),
.B(n_1801),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3576),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3591),
.A2(n_3441),
.B1(n_3414),
.B2(n_3359),
.Y(n_3789)
);

OAI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3704),
.A2(n_3432),
.B1(n_3347),
.B2(n_3406),
.Y(n_3790)
);

INVx3_ASAP7_75t_L g3791 ( 
.A(n_3699),
.Y(n_3791)
);

INVx1_ASAP7_75t_SL g3792 ( 
.A(n_3627),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3572),
.B(n_3528),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3568),
.Y(n_3794)
);

INVx1_ASAP7_75t_SL g3795 ( 
.A(n_3710),
.Y(n_3795)
);

INVx4_ASAP7_75t_L g3796 ( 
.A(n_3574),
.Y(n_3796)
);

BUFx2_ASAP7_75t_L g3797 ( 
.A(n_3663),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3749),
.A2(n_3542),
.B1(n_3415),
.B2(n_3429),
.Y(n_3798)
);

NOR2xp33_ASAP7_75t_L g3799 ( 
.A(n_3607),
.B(n_3490),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3595),
.B(n_3490),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3594),
.A2(n_3449),
.B(n_3442),
.Y(n_3801)
);

BUFx6f_ASAP7_75t_L g3802 ( 
.A(n_3574),
.Y(n_3802)
);

NAND2xp33_ASAP7_75t_L g3803 ( 
.A(n_3766),
.B(n_3529),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3605),
.Y(n_3804)
);

BUFx6f_ASAP7_75t_L g3805 ( 
.A(n_3574),
.Y(n_3805)
);

O2A1O1Ixp5_ASAP7_75t_SL g3806 ( 
.A1(n_3573),
.A2(n_1420),
.B(n_1421),
.C(n_1418),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3610),
.Y(n_3807)
);

INVx3_ASAP7_75t_L g3808 ( 
.A(n_3699),
.Y(n_3808)
);

BUFx6f_ASAP7_75t_L g3809 ( 
.A(n_3579),
.Y(n_3809)
);

INVx1_ASAP7_75t_SL g3810 ( 
.A(n_3775),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_3587),
.B(n_3449),
.Y(n_3811)
);

OA21x2_ASAP7_75t_L g3812 ( 
.A1(n_3580),
.A2(n_1427),
.B(n_1425),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3577),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_3683),
.B(n_3490),
.Y(n_3814)
);

AO22x1_ASAP7_75t_L g3815 ( 
.A1(n_3784),
.A2(n_3509),
.B1(n_3415),
.B2(n_3429),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3621),
.Y(n_3816)
);

AND2x4_ASAP7_75t_L g3817 ( 
.A(n_3682),
.B(n_3509),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3589),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3622),
.Y(n_3819)
);

OR2x6_ASAP7_75t_L g3820 ( 
.A(n_3707),
.B(n_3472),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_SL g3821 ( 
.A1(n_3569),
.A2(n_3513),
.B(n_3516),
.C(n_3464),
.Y(n_3821)
);

CKINVDCx5p33_ASAP7_75t_R g3822 ( 
.A(n_3772),
.Y(n_3822)
);

INVx2_ASAP7_75t_SL g3823 ( 
.A(n_3653),
.Y(n_3823)
);

INVx2_ASAP7_75t_SL g3824 ( 
.A(n_3583),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3644),
.Y(n_3825)
);

INVx3_ASAP7_75t_L g3826 ( 
.A(n_3700),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_3647),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3649),
.Y(n_3828)
);

INVx2_ASAP7_75t_L g3829 ( 
.A(n_3603),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3582),
.B(n_3518),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3575),
.A2(n_792),
.B1(n_827),
.B2(n_767),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3630),
.Y(n_3832)
);

BUFx2_ASAP7_75t_L g3833 ( 
.A(n_3786),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3570),
.B(n_3518),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_SL g3835 ( 
.A(n_3609),
.B(n_3555),
.Y(n_3835)
);

OAI22xp5_ASAP7_75t_L g3836 ( 
.A1(n_3631),
.A2(n_3402),
.B1(n_3513),
.B2(n_3464),
.Y(n_3836)
);

NOR2xp33_ASAP7_75t_L g3837 ( 
.A(n_3715),
.B(n_3518),
.Y(n_3837)
);

INVx2_ASAP7_75t_SL g3838 ( 
.A(n_3701),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3581),
.B(n_3565),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3650),
.Y(n_3840)
);

CKINVDCx5p33_ASAP7_75t_R g3841 ( 
.A(n_3713),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3584),
.Y(n_3842)
);

AOI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3661),
.A2(n_827),
.B1(n_846),
.B2(n_792),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3637),
.Y(n_3844)
);

AND2x4_ASAP7_75t_L g3845 ( 
.A(n_3682),
.B(n_3516),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3641),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3712),
.B(n_3524),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3676),
.B(n_3524),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3665),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3700),
.Y(n_3850)
);

OAI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3566),
.A2(n_3402),
.B1(n_902),
.B2(n_903),
.Y(n_3851)
);

BUFx2_ASAP7_75t_L g3852 ( 
.A(n_3593),
.Y(n_3852)
);

BUFx3_ASAP7_75t_L g3853 ( 
.A(n_3745),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3648),
.Y(n_3854)
);

AOI22xp33_ASAP7_75t_L g3855 ( 
.A1(n_3729),
.A2(n_1021),
.B1(n_1036),
.B2(n_846),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3655),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3629),
.B(n_3524),
.Y(n_3857)
);

AOI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3604),
.A2(n_904),
.B1(n_905),
.B2(n_897),
.Y(n_3858)
);

NOR2xp33_ASAP7_75t_L g3859 ( 
.A(n_3598),
.B(n_890),
.Y(n_3859)
);

OR2x6_ASAP7_75t_L g3860 ( 
.A(n_3638),
.B(n_3555),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3677),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3659),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3693),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3698),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3567),
.B(n_1530),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3675),
.B(n_3717),
.Y(n_3866)
);

AOI22xp5_ASAP7_75t_L g3867 ( 
.A1(n_3738),
.A2(n_910),
.B1(n_912),
.B2(n_907),
.Y(n_3867)
);

INVx4_ASAP7_75t_L g3868 ( 
.A(n_3579),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3724),
.Y(n_3869)
);

INVx2_ASAP7_75t_SL g3870 ( 
.A(n_3696),
.Y(n_3870)
);

INVx2_ASAP7_75t_SL g3871 ( 
.A(n_3773),
.Y(n_3871)
);

AOI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3632),
.A2(n_922),
.B1(n_923),
.B2(n_921),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3579),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3666),
.Y(n_3874)
);

AND3x1_ASAP7_75t_SL g3875 ( 
.A(n_3736),
.B(n_1431),
.C(n_1430),
.Y(n_3875)
);

BUFx12f_ASAP7_75t_L g3876 ( 
.A(n_3702),
.Y(n_3876)
);

HB1xp67_ASAP7_75t_L g3877 ( 
.A(n_3785),
.Y(n_3877)
);

BUFx6f_ASAP7_75t_L g3878 ( 
.A(n_3615),
.Y(n_3878)
);

BUFx12f_ASAP7_75t_L g3879 ( 
.A(n_3757),
.Y(n_3879)
);

NAND2x1_ASAP7_75t_L g3880 ( 
.A(n_3671),
.B(n_2647),
.Y(n_3880)
);

INVx3_ASAP7_75t_L g3881 ( 
.A(n_3615),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3703),
.B(n_1532),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3586),
.A2(n_3561),
.B1(n_926),
.B2(n_928),
.Y(n_3883)
);

INVx3_ASAP7_75t_L g3884 ( 
.A(n_3615),
.Y(n_3884)
);

OAI21x1_ASAP7_75t_SL g3885 ( 
.A1(n_3751),
.A2(n_1438),
.B(n_1433),
.Y(n_3885)
);

HB1xp67_ASAP7_75t_L g3886 ( 
.A(n_3640),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3678),
.Y(n_3887)
);

OAI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_3657),
.A2(n_930),
.B1(n_933),
.B2(n_924),
.Y(n_3888)
);

AOI21xp33_ASAP7_75t_L g3889 ( 
.A1(n_3585),
.A2(n_1442),
.B(n_1439),
.Y(n_3889)
);

BUFx3_ASAP7_75t_L g3890 ( 
.A(n_3625),
.Y(n_3890)
);

BUFx6f_ASAP7_75t_L g3891 ( 
.A(n_3619),
.Y(n_3891)
);

BUFx6f_ASAP7_75t_L g3892 ( 
.A(n_3619),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_L g3893 ( 
.A1(n_3777),
.A2(n_1021),
.B1(n_1036),
.B2(n_846),
.Y(n_3893)
);

CKINVDCx20_ASAP7_75t_R g3894 ( 
.A(n_3686),
.Y(n_3894)
);

BUFx3_ASAP7_75t_L g3895 ( 
.A(n_3670),
.Y(n_3895)
);

BUFx2_ASAP7_75t_L g3896 ( 
.A(n_3654),
.Y(n_3896)
);

INVx4_ASAP7_75t_L g3897 ( 
.A(n_3619),
.Y(n_3897)
);

AND2x6_ASAP7_75t_SL g3898 ( 
.A(n_3753),
.B(n_3732),
.Y(n_3898)
);

BUFx8_ASAP7_75t_L g3899 ( 
.A(n_3643),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3668),
.B(n_3601),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3642),
.A2(n_940),
.B1(n_941),
.B2(n_934),
.Y(n_3901)
);

HB1xp67_ASAP7_75t_L g3902 ( 
.A(n_3747),
.Y(n_3902)
);

BUFx3_ASAP7_75t_L g3903 ( 
.A(n_3697),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3744),
.Y(n_3904)
);

BUFx3_ASAP7_75t_L g3905 ( 
.A(n_3654),
.Y(n_3905)
);

CKINVDCx5p33_ASAP7_75t_R g3906 ( 
.A(n_3646),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3754),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_3679),
.Y(n_3908)
);

OAI22xp5_ASAP7_75t_L g3909 ( 
.A1(n_3721),
.A2(n_946),
.B1(n_947),
.B2(n_943),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_3620),
.A2(n_2559),
.B(n_2544),
.Y(n_3910)
);

INVx1_ASAP7_75t_SL g3911 ( 
.A(n_3611),
.Y(n_3911)
);

O2A1O1Ixp33_ASAP7_75t_L g3912 ( 
.A1(n_3592),
.A2(n_1444),
.B(n_1447),
.C(n_1446),
.Y(n_3912)
);

HB1xp67_ASAP7_75t_L g3913 ( 
.A(n_3758),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3770),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_L g3915 ( 
.A(n_3720),
.B(n_899),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3761),
.Y(n_3916)
);

OAI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_3612),
.A2(n_959),
.B1(n_963),
.B2(n_948),
.Y(n_3917)
);

AND2x4_ASAP7_75t_L g3918 ( 
.A(n_3708),
.B(n_2647),
.Y(n_3918)
);

INVx3_ASAP7_75t_SL g3919 ( 
.A(n_3780),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3602),
.A2(n_968),
.B1(n_970),
.B2(n_967),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3664),
.B(n_1535),
.Y(n_3921)
);

BUFx2_ASAP7_75t_L g3922 ( 
.A(n_3654),
.Y(n_3922)
);

AND2x4_ASAP7_75t_L g3923 ( 
.A(n_3708),
.B(n_2655),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3624),
.B(n_1448),
.Y(n_3924)
);

INVx3_ASAP7_75t_L g3925 ( 
.A(n_3643),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3618),
.B(n_1807),
.Y(n_3926)
);

AND2x4_ASAP7_75t_L g3927 ( 
.A(n_3578),
.B(n_2655),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3578),
.B(n_2697),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3771),
.Y(n_3929)
);

INVx3_ASAP7_75t_L g3930 ( 
.A(n_3643),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3760),
.Y(n_3931)
);

INVx4_ASAP7_75t_L g3932 ( 
.A(n_3651),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3762),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3633),
.B(n_1807),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3734),
.Y(n_3935)
);

O2A1O1Ixp33_ASAP7_75t_L g3936 ( 
.A1(n_3588),
.A2(n_1450),
.B(n_1455),
.C(n_1451),
.Y(n_3936)
);

BUFx6f_ASAP7_75t_L g3937 ( 
.A(n_3651),
.Y(n_3937)
);

OAI22xp5_ASAP7_75t_L g3938 ( 
.A1(n_3616),
.A2(n_975),
.B1(n_976),
.B2(n_974),
.Y(n_3938)
);

INVx1_ASAP7_75t_SL g3939 ( 
.A(n_3735),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3740),
.Y(n_3940)
);

NAND2x2_ASAP7_75t_L g3941 ( 
.A(n_3787),
.B(n_1390),
.Y(n_3941)
);

BUFx2_ASAP7_75t_L g3942 ( 
.A(n_3660),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3680),
.A2(n_1021),
.B1(n_1036),
.B2(n_846),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_3735),
.B(n_900),
.Y(n_3944)
);

INVxp67_ASAP7_75t_L g3945 ( 
.A(n_3660),
.Y(n_3945)
);

O2A1O1Ixp5_ASAP7_75t_L g3946 ( 
.A1(n_3673),
.A2(n_1458),
.B(n_1459),
.C(n_1457),
.Y(n_3946)
);

AOI22xp33_ASAP7_75t_L g3947 ( 
.A1(n_3680),
.A2(n_1036),
.B1(n_1021),
.B2(n_1463),
.Y(n_3947)
);

AND2x4_ASAP7_75t_L g3948 ( 
.A(n_3759),
.B(n_2697),
.Y(n_3948)
);

BUFx6f_ASAP7_75t_L g3949 ( 
.A(n_3651),
.Y(n_3949)
);

OR2x6_ASAP7_75t_L g3950 ( 
.A(n_3746),
.B(n_1812),
.Y(n_3950)
);

BUFx6f_ASAP7_75t_L g3951 ( 
.A(n_3660),
.Y(n_3951)
);

CKINVDCx20_ASAP7_75t_R g3952 ( 
.A(n_3681),
.Y(n_3952)
);

AOI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3680),
.A2(n_1468),
.B1(n_1469),
.B2(n_1464),
.Y(n_3953)
);

NAND2x1p5_ASAP7_75t_L g3954 ( 
.A(n_3671),
.B(n_2697),
.Y(n_3954)
);

INVx5_ASAP7_75t_L g3955 ( 
.A(n_3739),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3776),
.Y(n_3956)
);

INVx4_ASAP7_75t_L g3957 ( 
.A(n_3681),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3680),
.A2(n_1475),
.B1(n_1486),
.B2(n_1473),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3626),
.A2(n_2544),
.B(n_2710),
.Y(n_3959)
);

BUFx3_ASAP7_75t_L g3960 ( 
.A(n_3681),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_SL g3961 ( 
.A(n_3680),
.B(n_1708),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3750),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3711),
.B(n_1812),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3635),
.A2(n_2710),
.B(n_2408),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3755),
.Y(n_3965)
);

INVx4_ASAP7_75t_L g3966 ( 
.A(n_3695),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3695),
.Y(n_3967)
);

INVx4_ASAP7_75t_L g3968 ( 
.A(n_3695),
.Y(n_3968)
);

INVx2_ASAP7_75t_SL g3969 ( 
.A(n_3709),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3709),
.Y(n_3970)
);

BUFx3_ASAP7_75t_L g3971 ( 
.A(n_3709),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3727),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_3741),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3741),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3674),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3741),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3634),
.A2(n_2710),
.B(n_2408),
.Y(n_3977)
);

OR2x6_ASAP7_75t_L g3978 ( 
.A(n_3667),
.B(n_2203),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3739),
.Y(n_3979)
);

AND2x4_ASAP7_75t_L g3980 ( 
.A(n_3759),
.B(n_2710),
.Y(n_3980)
);

OR2x6_ASAP7_75t_L g3981 ( 
.A(n_3743),
.B(n_2204),
.Y(n_3981)
);

INVx3_ASAP7_75t_L g3982 ( 
.A(n_3767),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3571),
.B(n_979),
.Y(n_3983)
);

AOI22xp33_ASAP7_75t_L g3984 ( 
.A1(n_3684),
.A2(n_1489),
.B1(n_1490),
.B2(n_1487),
.Y(n_3984)
);

INVx3_ASAP7_75t_L g3985 ( 
.A(n_3767),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3597),
.B(n_980),
.Y(n_3986)
);

A2O1A1Ixp33_ASAP7_75t_L g3987 ( 
.A1(n_3564),
.A2(n_1492),
.B(n_1494),
.C(n_1491),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3714),
.B(n_982),
.Y(n_3988)
);

BUFx12f_ASAP7_75t_L g3989 ( 
.A(n_3728),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3599),
.Y(n_3990)
);

INVx2_ASAP7_75t_SL g3991 ( 
.A(n_3778),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3737),
.B(n_1700),
.Y(n_3992)
);

INVx2_ASAP7_75t_SL g3993 ( 
.A(n_3783),
.Y(n_3993)
);

BUFx2_ASAP7_75t_L g3994 ( 
.A(n_3623),
.Y(n_3994)
);

AOI221xp5_ASAP7_75t_L g3995 ( 
.A1(n_3756),
.A2(n_986),
.B1(n_987),
.B2(n_985),
.C(n_983),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3706),
.Y(n_3996)
);

A2O1A1Ixp33_ASAP7_75t_L g3997 ( 
.A1(n_3590),
.A2(n_1080),
.B(n_1053),
.C(n_991),
.Y(n_3997)
);

AOI21xp5_ASAP7_75t_L g3998 ( 
.A1(n_3617),
.A2(n_2408),
.B(n_2369),
.Y(n_3998)
);

BUFx6f_ASAP7_75t_L g3999 ( 
.A(n_3752),
.Y(n_3999)
);

A2O1A1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_3606),
.A2(n_1045),
.B(n_1059),
.C(n_999),
.Y(n_4000)
);

BUFx6f_ASAP7_75t_L g4001 ( 
.A(n_3636),
.Y(n_4001)
);

BUFx6f_ASAP7_75t_L g4002 ( 
.A(n_3765),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3672),
.A2(n_992),
.B1(n_994),
.B2(n_988),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3782),
.Y(n_4004)
);

BUFx6f_ASAP7_75t_L g4005 ( 
.A(n_3768),
.Y(n_4005)
);

INVxp67_ASAP7_75t_L g4006 ( 
.A(n_3779),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3764),
.B(n_909),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3731),
.Y(n_4008)
);

AOI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_3656),
.A2(n_2408),
.B(n_2369),
.Y(n_4009)
);

INVx5_ASAP7_75t_L g4010 ( 
.A(n_3781),
.Y(n_4010)
);

INVx3_ASAP7_75t_L g4011 ( 
.A(n_3692),
.Y(n_4011)
);

INVx3_ASAP7_75t_L g4012 ( 
.A(n_3763),
.Y(n_4012)
);

BUFx2_ASAP7_75t_L g4013 ( 
.A(n_3718),
.Y(n_4013)
);

INVxp67_ASAP7_75t_SL g4014 ( 
.A(n_3600),
.Y(n_4014)
);

INVx2_ASAP7_75t_SL g4015 ( 
.A(n_3723),
.Y(n_4015)
);

A2O1A1Ixp33_ASAP7_75t_L g4016 ( 
.A1(n_4007),
.A2(n_3628),
.B(n_3652),
.C(n_3596),
.Y(n_4016)
);

O2A1O1Ixp33_ASAP7_75t_SL g4017 ( 
.A1(n_4000),
.A2(n_3719),
.B(n_3669),
.C(n_3658),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3851),
.A2(n_1010),
.B1(n_1012),
.B2(n_1005),
.Y(n_4018)
);

AOI22xp5_ASAP7_75t_L g4019 ( 
.A1(n_4004),
.A2(n_1015),
.B1(n_1017),
.B2(n_1013),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3929),
.Y(n_4020)
);

INVxp33_ASAP7_75t_SL g4021 ( 
.A(n_3822),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_4014),
.A2(n_3685),
.B(n_3662),
.Y(n_4022)
);

AND2x4_ASAP7_75t_L g4023 ( 
.A(n_3797),
.B(n_3733),
.Y(n_4023)
);

NOR2xp33_ASAP7_75t_L g4024 ( 
.A(n_3792),
.B(n_1030),
.Y(n_4024)
);

NOR2xp33_ASAP7_75t_L g4025 ( 
.A(n_3906),
.B(n_3894),
.Y(n_4025)
);

O2A1O1Ixp33_ASAP7_75t_SL g4026 ( 
.A1(n_3908),
.A2(n_3688),
.B(n_3691),
.C(n_3742),
.Y(n_4026)
);

CKINVDCx5p33_ASAP7_75t_R g4027 ( 
.A(n_3876),
.Y(n_4027)
);

NOR2xp33_ASAP7_75t_L g4028 ( 
.A(n_3895),
.B(n_1038),
.Y(n_4028)
);

O2A1O1Ixp33_ASAP7_75t_SL g4029 ( 
.A1(n_3821),
.A2(n_3705),
.B(n_3748),
.C(n_3690),
.Y(n_4029)
);

OR2x2_ASAP7_75t_L g4030 ( 
.A(n_3877),
.B(n_3608),
.Y(n_4030)
);

INVx3_ASAP7_75t_L g4031 ( 
.A(n_3802),
.Y(n_4031)
);

AOI221xp5_ASAP7_75t_L g4032 ( 
.A1(n_3920),
.A2(n_1046),
.B1(n_1049),
.B2(n_1040),
.C(n_1039),
.Y(n_4032)
);

INVx1_ASAP7_75t_SL g4033 ( 
.A(n_3903),
.Y(n_4033)
);

AO21x2_ASAP7_75t_L g4034 ( 
.A1(n_3964),
.A2(n_3730),
.B(n_3725),
.Y(n_4034)
);

O2A1O1Ixp33_ASAP7_75t_SL g4035 ( 
.A1(n_3997),
.A2(n_3769),
.B(n_3645),
.C(n_3639),
.Y(n_4035)
);

CKINVDCx11_ASAP7_75t_R g4036 ( 
.A(n_3898),
.Y(n_4036)
);

AO31x2_ASAP7_75t_L g4037 ( 
.A1(n_3972),
.A2(n_3689),
.A3(n_3694),
.B(n_3613),
.Y(n_4037)
);

AO31x2_ASAP7_75t_L g4038 ( 
.A1(n_3940),
.A2(n_3722),
.A3(n_3774),
.B(n_2206),
.Y(n_4038)
);

AOI22xp33_ASAP7_75t_L g4039 ( 
.A1(n_4013),
.A2(n_1051),
.B1(n_1052),
.B2(n_1050),
.Y(n_4039)
);

INVx2_ASAP7_75t_SL g4040 ( 
.A(n_3853),
.Y(n_4040)
);

AOI31xp67_ASAP7_75t_L g4041 ( 
.A1(n_3961),
.A2(n_3835),
.A3(n_3811),
.B(n_3988),
.Y(n_4041)
);

CKINVDCx20_ASAP7_75t_R g4042 ( 
.A(n_3952),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3994),
.A2(n_3614),
.B(n_3726),
.Y(n_4043)
);

INVx2_ASAP7_75t_L g4044 ( 
.A(n_3788),
.Y(n_4044)
);

OAI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_4006),
.A2(n_1088),
.B1(n_1062),
.B2(n_1064),
.Y(n_4045)
);

OAI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_3983),
.A2(n_3716),
.B(n_3687),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_SL g4047 ( 
.A1(n_4003),
.A2(n_12),
.B(n_23),
.C(n_4),
.Y(n_4047)
);

HB1xp67_ASAP7_75t_L g4048 ( 
.A(n_3842),
.Y(n_4048)
);

AOI221xp5_ASAP7_75t_L g4049 ( 
.A1(n_3917),
.A2(n_1075),
.B1(n_1078),
.B2(n_1070),
.C(n_1057),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_3841),
.Y(n_4050)
);

BUFx2_ASAP7_75t_L g4051 ( 
.A(n_3852),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3801),
.A2(n_915),
.B(n_911),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3800),
.B(n_5),
.Y(n_4053)
);

O2A1O1Ixp33_ASAP7_75t_SL g4054 ( 
.A1(n_3900),
.A2(n_16),
.B(n_27),
.C(n_6),
.Y(n_4054)
);

CKINVDCx12_ASAP7_75t_R g4055 ( 
.A(n_3847),
.Y(n_4055)
);

O2A1O1Ixp33_ASAP7_75t_L g4056 ( 
.A1(n_3889),
.A2(n_1738),
.B(n_1747),
.C(n_1700),
.Y(n_4056)
);

O2A1O1Ixp33_ASAP7_75t_SL g4057 ( 
.A1(n_3839),
.A2(n_19),
.B(n_31),
.C(n_7),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3804),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3933),
.B(n_1711),
.Y(n_4059)
);

OAI21x1_ASAP7_75t_L g4060 ( 
.A1(n_3959),
.A2(n_1738),
.B(n_1700),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3913),
.Y(n_4061)
);

AOI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3837),
.A2(n_1093),
.B1(n_1095),
.B2(n_1091),
.Y(n_4062)
);

OAI211xp5_ASAP7_75t_L g4063 ( 
.A1(n_3831),
.A2(n_1098),
.B(n_1097),
.C(n_918),
.Y(n_4063)
);

AOI21xp5_ASAP7_75t_L g4064 ( 
.A1(n_3986),
.A2(n_920),
.B(n_916),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3807),
.Y(n_4065)
);

BUFx5_ASAP7_75t_L g4066 ( 
.A(n_3975),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3866),
.B(n_1738),
.Y(n_4067)
);

A2O1A1Ixp33_ASAP7_75t_L g4068 ( 
.A1(n_3859),
.A2(n_935),
.B(n_936),
.C(n_925),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3816),
.Y(n_4069)
);

O2A1O1Ixp33_ASAP7_75t_L g4070 ( 
.A1(n_3990),
.A2(n_1749),
.B(n_1792),
.C(n_1747),
.Y(n_4070)
);

BUFx12f_ASAP7_75t_L g4071 ( 
.A(n_3899),
.Y(n_4071)
);

INVx1_ASAP7_75t_SL g4072 ( 
.A(n_3795),
.Y(n_4072)
);

A2O1A1Ixp33_ASAP7_75t_L g4073 ( 
.A1(n_3843),
.A2(n_942),
.B(n_945),
.C(n_938),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3902),
.B(n_1747),
.Y(n_4074)
);

OAI21x1_ASAP7_75t_L g4075 ( 
.A1(n_3977),
.A2(n_1792),
.B(n_1749),
.Y(n_4075)
);

CKINVDCx16_ASAP7_75t_R g4076 ( 
.A(n_3834),
.Y(n_4076)
);

AOI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3910),
.A2(n_964),
.B(n_949),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3819),
.Y(n_4078)
);

OAI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_3946),
.A2(n_993),
.B(n_969),
.Y(n_4079)
);

HB1xp67_ASAP7_75t_L g4080 ( 
.A(n_3886),
.Y(n_4080)
);

A2O1A1Ixp33_ASAP7_75t_L g4081 ( 
.A1(n_3893),
.A2(n_3912),
.B(n_3996),
.C(n_3943),
.Y(n_4081)
);

NOR2xp67_ASAP7_75t_R g4082 ( 
.A(n_4011),
.B(n_1749),
.Y(n_4082)
);

O2A1O1Ixp33_ASAP7_75t_SL g4083 ( 
.A1(n_3993),
.A2(n_19),
.B(n_31),
.C(n_7),
.Y(n_4083)
);

O2A1O1Ixp33_ASAP7_75t_L g4084 ( 
.A1(n_3888),
.A2(n_1797),
.B(n_1792),
.C(n_1632),
.Y(n_4084)
);

AOI21xp5_ASAP7_75t_L g4085 ( 
.A1(n_3815),
.A2(n_998),
.B(n_995),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3825),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3911),
.B(n_1020),
.Y(n_4087)
);

O2A1O1Ixp33_ASAP7_75t_SL g4088 ( 
.A1(n_3790),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3857),
.B(n_10),
.Y(n_4089)
);

AND2x4_ASAP7_75t_L g4090 ( 
.A(n_3833),
.B(n_406),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_3827),
.Y(n_4091)
);

BUFx2_ASAP7_75t_L g4092 ( 
.A(n_3890),
.Y(n_4092)
);

AND2x4_ASAP7_75t_L g4093 ( 
.A(n_3870),
.B(n_3871),
.Y(n_4093)
);

A2O1A1Ixp33_ASAP7_75t_L g4094 ( 
.A1(n_3872),
.A2(n_1027),
.B(n_1032),
.C(n_1024),
.Y(n_4094)
);

NAND2x2_ASAP7_75t_L g4095 ( 
.A(n_3824),
.B(n_11),
.Y(n_4095)
);

BUFx6f_ASAP7_75t_L g4096 ( 
.A(n_3951),
.Y(n_4096)
);

AO31x2_ASAP7_75t_L g4097 ( 
.A1(n_3998),
.A2(n_4008),
.A3(n_4009),
.B(n_3840),
.Y(n_4097)
);

OAI22xp33_ASAP7_75t_L g4098 ( 
.A1(n_3919),
.A2(n_1047),
.B1(n_1041),
.B2(n_1711),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3828),
.Y(n_4099)
);

BUFx10_ASAP7_75t_L g4100 ( 
.A(n_3944),
.Y(n_4100)
);

CKINVDCx11_ASAP7_75t_R g4101 ( 
.A(n_3989),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3849),
.Y(n_4102)
);

AO31x2_ASAP7_75t_L g4103 ( 
.A1(n_3861),
.A2(n_2206),
.A3(n_2213),
.B(n_2204),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3810),
.B(n_1797),
.Y(n_4104)
);

OA21x2_ASAP7_75t_L g4105 ( 
.A1(n_3916),
.A2(n_1632),
.B(n_1630),
.Y(n_4105)
);

OAI21x1_ASAP7_75t_L g4106 ( 
.A1(n_4012),
.A2(n_1797),
.B(n_2213),
.Y(n_4106)
);

INVx3_ASAP7_75t_L g4107 ( 
.A(n_3802),
.Y(n_4107)
);

AOI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3815),
.A2(n_2221),
.B(n_2220),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3931),
.B(n_1630),
.Y(n_4109)
);

OA21x2_ASAP7_75t_L g4110 ( 
.A1(n_3863),
.A2(n_2221),
.B(n_2220),
.Y(n_4110)
);

OAI21xp5_ASAP7_75t_L g4111 ( 
.A1(n_3984),
.A2(n_2844),
.B(n_2842),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3864),
.Y(n_4112)
);

OR2x2_ASAP7_75t_L g4113 ( 
.A(n_3869),
.B(n_1711),
.Y(n_4113)
);

INVx2_ASAP7_75t_L g4114 ( 
.A(n_3904),
.Y(n_4114)
);

INVx1_ASAP7_75t_SL g4115 ( 
.A(n_3939),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3907),
.Y(n_4116)
);

OR2x2_ASAP7_75t_L g4117 ( 
.A(n_3914),
.B(n_1711),
.Y(n_4117)
);

A2O1A1Ixp33_ASAP7_75t_L g4118 ( 
.A1(n_3936),
.A2(n_1716),
.B(n_1734),
.C(n_1714),
.Y(n_4118)
);

AO22x2_ASAP7_75t_L g4119 ( 
.A1(n_4011),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_4119)
);

OAI21x1_ASAP7_75t_L g4120 ( 
.A1(n_4012),
.A2(n_3812),
.B(n_3806),
.Y(n_4120)
);

OA21x2_ASAP7_75t_L g4121 ( 
.A1(n_3987),
.A2(n_2228),
.B(n_2224),
.Y(n_4121)
);

AO32x2_ASAP7_75t_L g4122 ( 
.A1(n_3991),
.A2(n_17),
.A3(n_13),
.B1(n_14),
.B2(n_21),
.Y(n_4122)
);

AOI221xp5_ASAP7_75t_L g4123 ( 
.A1(n_3855),
.A2(n_1734),
.B1(n_1737),
.B2(n_1716),
.C(n_1714),
.Y(n_4123)
);

AOI22xp33_ASAP7_75t_SL g4124 ( 
.A1(n_4005),
.A2(n_1716),
.B1(n_1734),
.B2(n_1714),
.Y(n_4124)
);

OAI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3789),
.A2(n_1716),
.B1(n_1734),
.B2(n_1714),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_3799),
.B(n_3915),
.Y(n_4126)
);

INVx3_ASAP7_75t_L g4127 ( 
.A(n_3802),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3794),
.Y(n_4128)
);

O2A1O1Ixp33_ASAP7_75t_SL g4129 ( 
.A1(n_3880),
.A2(n_22),
.B(n_17),
.C(n_21),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_3830),
.B(n_23),
.Y(n_4130)
);

AO31x2_ASAP7_75t_L g4131 ( 
.A1(n_3836),
.A2(n_2228),
.A3(n_2232),
.B(n_2224),
.Y(n_4131)
);

AOI21xp5_ASAP7_75t_L g4132 ( 
.A1(n_3812),
.A2(n_2232),
.B(n_2369),
.Y(n_4132)
);

INVx3_ASAP7_75t_L g4133 ( 
.A(n_3805),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3813),
.Y(n_4134)
);

INVx3_ASAP7_75t_SL g4135 ( 
.A(n_3823),
.Y(n_4135)
);

AO31x2_ASAP7_75t_L g4136 ( 
.A1(n_3979),
.A2(n_3935),
.A3(n_3829),
.B(n_3832),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3818),
.Y(n_4137)
);

AOI22xp33_ASAP7_75t_L g4138 ( 
.A1(n_4015),
.A2(n_1743),
.B1(n_1748),
.B2(n_1737),
.Y(n_4138)
);

AO31x2_ASAP7_75t_L g4139 ( 
.A1(n_3844),
.A2(n_1562),
.A3(n_1597),
.B(n_1509),
.Y(n_4139)
);

INVx3_ASAP7_75t_L g4140 ( 
.A(n_3805),
.Y(n_4140)
);

INVx2_ASAP7_75t_SL g4141 ( 
.A(n_3951),
.Y(n_4141)
);

AND2x4_ASAP7_75t_L g4142 ( 
.A(n_3838),
.B(n_411),
.Y(n_4142)
);

AOI22xp33_ASAP7_75t_L g4143 ( 
.A1(n_3941),
.A2(n_1743),
.B1(n_1748),
.B2(n_1737),
.Y(n_4143)
);

AOI21xp5_ASAP7_75t_L g4144 ( 
.A1(n_3950),
.A2(n_2449),
.B(n_2369),
.Y(n_4144)
);

AOI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_3814),
.A2(n_1743),
.B1(n_1748),
.B2(n_1737),
.Y(n_4145)
);

NAND2x1p5_ASAP7_75t_L g4146 ( 
.A(n_3955),
.B(n_2230),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_L g4147 ( 
.A1(n_3950),
.A2(n_2457),
.B(n_2449),
.Y(n_4147)
);

AOI22xp33_ASAP7_75t_L g4148 ( 
.A1(n_4005),
.A2(n_1748),
.B1(n_1750),
.B2(n_1743),
.Y(n_4148)
);

O2A1O1Ixp5_ASAP7_75t_L g4149 ( 
.A1(n_3798),
.A2(n_2240),
.B(n_2230),
.C(n_1518),
.Y(n_4149)
);

A2O1A1Ixp33_ASAP7_75t_L g4150 ( 
.A1(n_3947),
.A2(n_1754),
.B(n_1786),
.C(n_1750),
.Y(n_4150)
);

A2O1A1Ixp33_ASAP7_75t_L g4151 ( 
.A1(n_3858),
.A2(n_1754),
.B(n_1786),
.C(n_1750),
.Y(n_4151)
);

OAI21x1_ASAP7_75t_L g4152 ( 
.A1(n_3992),
.A2(n_2240),
.B(n_2230),
.Y(n_4152)
);

AO32x2_ASAP7_75t_L g4153 ( 
.A1(n_3938),
.A2(n_27),
.A3(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_4153)
);

O2A1O1Ixp33_ASAP7_75t_SL g4154 ( 
.A1(n_3793),
.A2(n_34),
.B(n_26),
.C(n_33),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3846),
.Y(n_4155)
);

NOR2xp33_ASAP7_75t_SL g4156 ( 
.A(n_3879),
.B(n_2842),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3854),
.Y(n_4157)
);

NAND3xp33_ASAP7_75t_L g4158 ( 
.A(n_3995),
.B(n_1754),
.C(n_1750),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3856),
.Y(n_4159)
);

O2A1O1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_3901),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_4160)
);

INVxp67_ASAP7_75t_L g4161 ( 
.A(n_3848),
.Y(n_4161)
);

NOR2xp33_ASAP7_75t_SL g4162 ( 
.A(n_3796),
.B(n_2842),
.Y(n_4162)
);

AOI22xp33_ASAP7_75t_L g4163 ( 
.A1(n_4005),
.A2(n_1786),
.B1(n_1787),
.B2(n_1754),
.Y(n_4163)
);

HB1xp67_ASAP7_75t_L g4164 ( 
.A(n_3862),
.Y(n_4164)
);

BUFx10_ASAP7_75t_L g4165 ( 
.A(n_3820),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3896),
.B(n_3922),
.Y(n_4166)
);

O2A1O1Ixp33_ASAP7_75t_SL g4167 ( 
.A1(n_3945),
.A2(n_39),
.B(n_36),
.C(n_37),
.Y(n_4167)
);

HB1xp67_ASAP7_75t_L g4168 ( 
.A(n_3874),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_3942),
.B(n_39),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3956),
.B(n_40),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3963),
.A2(n_2457),
.B(n_2449),
.Y(n_4171)
);

OAI21x1_ASAP7_75t_L g4172 ( 
.A1(n_3791),
.A2(n_2240),
.B(n_1888),
.Y(n_4172)
);

AO31x2_ASAP7_75t_L g4173 ( 
.A1(n_3887),
.A2(n_1562),
.A3(n_1597),
.B(n_1509),
.Y(n_4173)
);

AOI221xp5_ASAP7_75t_L g4174 ( 
.A1(n_3909),
.A2(n_3883),
.B1(n_3867),
.B2(n_3924),
.C(n_3962),
.Y(n_4174)
);

CKINVDCx9p33_ASAP7_75t_R g4175 ( 
.A(n_3882),
.Y(n_4175)
);

OAI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3953),
.A2(n_2844),
.B(n_2842),
.Y(n_4176)
);

INVxp67_ASAP7_75t_SL g4177 ( 
.A(n_3934),
.Y(n_4177)
);

AOI22xp33_ASAP7_75t_L g4178 ( 
.A1(n_3958),
.A2(n_3965),
.B1(n_3885),
.B2(n_3928),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3921),
.Y(n_4179)
);

AO31x2_ASAP7_75t_L g4180 ( 
.A1(n_4001),
.A2(n_1562),
.A3(n_1597),
.B(n_1509),
.Y(n_4180)
);

O2A1O1Ixp33_ASAP7_75t_L g4181 ( 
.A1(n_3803),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_4181)
);

NOR2xp33_ASAP7_75t_L g4182 ( 
.A(n_3817),
.B(n_41),
.Y(n_4182)
);

A2O1A1Ixp33_ASAP7_75t_L g4183 ( 
.A1(n_3926),
.A2(n_1787),
.B(n_1789),
.C(n_1786),
.Y(n_4183)
);

INVx2_ASAP7_75t_SL g4184 ( 
.A(n_3951),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_SL g4185 ( 
.A(n_3796),
.B(n_2844),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3865),
.B(n_44),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_3927),
.A2(n_1787),
.B1(n_1790),
.B2(n_1789),
.Y(n_4187)
);

HB1xp67_ASAP7_75t_L g4188 ( 
.A(n_3955),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3982),
.B(n_45),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3967),
.Y(n_4190)
);

A2O1A1Ixp33_ASAP7_75t_L g4191 ( 
.A1(n_3927),
.A2(n_3928),
.B(n_3923),
.C(n_3918),
.Y(n_4191)
);

A2O1A1Ixp33_ASAP7_75t_L g4192 ( 
.A1(n_3918),
.A2(n_1789),
.B(n_1790),
.C(n_1787),
.Y(n_4192)
);

OAI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_3860),
.A2(n_2876),
.B(n_2844),
.Y(n_4193)
);

OR2x2_ASAP7_75t_L g4194 ( 
.A(n_3973),
.B(n_1789),
.Y(n_4194)
);

OAI21x1_ASAP7_75t_L g4195 ( 
.A1(n_3791),
.A2(n_1888),
.B(n_1871),
.Y(n_4195)
);

OAI22x1_ASAP7_75t_L g4196 ( 
.A1(n_3974),
.A2(n_3976),
.B1(n_3955),
.B2(n_3897),
.Y(n_4196)
);

BUFx10_ASAP7_75t_L g4197 ( 
.A(n_3820),
.Y(n_4197)
);

A2O1A1Ixp33_ASAP7_75t_L g4198 ( 
.A1(n_3923),
.A2(n_1798),
.B(n_1800),
.C(n_1790),
.Y(n_4198)
);

BUFx4f_ASAP7_75t_SL g4199 ( 
.A(n_3899),
.Y(n_4199)
);

AOI21xp5_ASAP7_75t_L g4200 ( 
.A1(n_3981),
.A2(n_2457),
.B(n_2449),
.Y(n_4200)
);

AO31x2_ASAP7_75t_L g4201 ( 
.A1(n_4001),
.A2(n_4010),
.A3(n_3897),
.B(n_3932),
.Y(n_4201)
);

A2O1A1Ixp33_ASAP7_75t_L g4202 ( 
.A1(n_3881),
.A2(n_3925),
.B(n_3930),
.C(n_3884),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_3982),
.B(n_45),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4001),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3985),
.B(n_46),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_3985),
.B(n_47),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3817),
.B(n_49),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3881),
.B(n_51),
.Y(n_4208)
);

OAI21xp5_ASAP7_75t_L g4209 ( 
.A1(n_3860),
.A2(n_2916),
.B(n_2908),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_3981),
.A2(n_2501),
.B(n_2457),
.Y(n_4210)
);

OAI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_3845),
.A2(n_1790),
.B1(n_1800),
.B2(n_1798),
.Y(n_4211)
);

O2A1O1Ixp33_ASAP7_75t_SL g4212 ( 
.A1(n_3969),
.A2(n_56),
.B(n_51),
.C(n_52),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_4010),
.A2(n_2908),
.A3(n_2916),
.B(n_2876),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_4010),
.A2(n_2501),
.B(n_1867),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3808),
.Y(n_4215)
);

O2A1O1Ixp33_ASAP7_75t_SL g4216 ( 
.A1(n_3884),
.A2(n_3930),
.B(n_3925),
.C(n_3826),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_3970),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_3905),
.Y(n_4218)
);

OAI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_3954),
.A2(n_3826),
.B(n_3808),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_3845),
.B(n_52),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3805),
.B(n_56),
.Y(n_4221)
);

AOI22xp33_ASAP7_75t_L g4222 ( 
.A1(n_4002),
.A2(n_3980),
.B1(n_3948),
.B2(n_3850),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_3978),
.A2(n_2501),
.B(n_1867),
.Y(n_4223)
);

NAND2x1p5_ASAP7_75t_L g4224 ( 
.A(n_3850),
.B(n_1859),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3970),
.Y(n_4225)
);

OAI21x1_ASAP7_75t_L g4226 ( 
.A1(n_3999),
.A2(n_1888),
.B(n_1871),
.Y(n_4226)
);

CKINVDCx11_ASAP7_75t_R g4227 ( 
.A(n_3809),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3809),
.B(n_57),
.Y(n_4228)
);

AOI22xp33_ASAP7_75t_L g4229 ( 
.A1(n_4002),
.A2(n_1798),
.B1(n_1811),
.B2(n_1800),
.Y(n_4229)
);

INVx2_ASAP7_75t_SL g4230 ( 
.A(n_3970),
.Y(n_4230)
);

OAI21x1_ASAP7_75t_L g4231 ( 
.A1(n_3999),
.A2(n_1889),
.B(n_1871),
.Y(n_4231)
);

OR2x2_ASAP7_75t_L g4232 ( 
.A(n_3960),
.B(n_1798),
.Y(n_4232)
);

AOI22xp33_ASAP7_75t_L g4233 ( 
.A1(n_4002),
.A2(n_1800),
.B1(n_1830),
.B2(n_1811),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3999),
.Y(n_4234)
);

O2A1O1Ixp33_ASAP7_75t_L g4235 ( 
.A1(n_3978),
.A2(n_62),
.B(n_57),
.C(n_60),
.Y(n_4235)
);

O2A1O1Ixp33_ASAP7_75t_L g4236 ( 
.A1(n_3948),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_4236)
);

O2A1O1Ixp33_ASAP7_75t_L g4237 ( 
.A1(n_3980),
.A2(n_68),
.B(n_65),
.C(n_67),
.Y(n_4237)
);

O2A1O1Ixp33_ASAP7_75t_L g4238 ( 
.A1(n_3875),
.A2(n_3971),
.B(n_71),
.C(n_69),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3809),
.Y(n_4239)
);

AO32x2_ASAP7_75t_L g4240 ( 
.A1(n_3957),
.A2(n_71),
.A3(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_4240)
);

INVx8_ASAP7_75t_L g4241 ( 
.A(n_3873),
.Y(n_4241)
);

AOI31xp67_ASAP7_75t_L g4242 ( 
.A1(n_3868),
.A2(n_2908),
.A3(n_2916),
.B(n_2876),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_3873),
.B(n_70),
.Y(n_4243)
);

INVx3_ASAP7_75t_L g4244 ( 
.A(n_3873),
.Y(n_4244)
);

OAI21xp5_ASAP7_75t_L g4245 ( 
.A1(n_3868),
.A2(n_2908),
.B(n_2876),
.Y(n_4245)
);

OAI21x1_ASAP7_75t_L g4246 ( 
.A1(n_3932),
.A2(n_1899),
.B(n_1889),
.Y(n_4246)
);

NOR2xp33_ASAP7_75t_L g4247 ( 
.A(n_3957),
.B(n_74),
.Y(n_4247)
);

AOI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_3878),
.A2(n_2501),
.B(n_1875),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_3878),
.B(n_75),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4044),
.Y(n_4250)
);

AOI22xp33_ASAP7_75t_L g4251 ( 
.A1(n_4036),
.A2(n_3891),
.B1(n_3892),
.B2(n_3878),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_L g4252 ( 
.A(n_4126),
.B(n_3966),
.Y(n_4252)
);

OAI22xp33_ASAP7_75t_SL g4253 ( 
.A1(n_4095),
.A2(n_3968),
.B1(n_3966),
.B2(n_77),
.Y(n_4253)
);

INVx3_ASAP7_75t_L g4254 ( 
.A(n_4023),
.Y(n_4254)
);

NAND2x1p5_ASAP7_75t_L g4255 ( 
.A(n_4092),
.B(n_3891),
.Y(n_4255)
);

INVx6_ASAP7_75t_L g4256 ( 
.A(n_4071),
.Y(n_4256)
);

BUFx2_ASAP7_75t_L g4257 ( 
.A(n_4051),
.Y(n_4257)
);

INVx1_ASAP7_75t_SL g4258 ( 
.A(n_4033),
.Y(n_4258)
);

NAND2xp33_ASAP7_75t_L g4259 ( 
.A(n_4081),
.B(n_3891),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4017),
.A2(n_3937),
.B(n_3892),
.Y(n_4260)
);

OAI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_4016),
.A2(n_3937),
.B1(n_3949),
.B2(n_3892),
.Y(n_4261)
);

AOI21x1_ASAP7_75t_L g4262 ( 
.A1(n_4085),
.A2(n_3968),
.B(n_3949),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4065),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_4178),
.A2(n_3949),
.B1(n_3937),
.B2(n_1830),
.Y(n_4264)
);

OR2x2_ASAP7_75t_L g4265 ( 
.A(n_4061),
.B(n_75),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4058),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4076),
.B(n_76),
.Y(n_4267)
);

AO31x2_ASAP7_75t_L g4268 ( 
.A1(n_4022),
.A2(n_80),
.A3(n_76),
.B(n_79),
.Y(n_4268)
);

INVx2_ASAP7_75t_SL g4269 ( 
.A(n_4135),
.Y(n_4269)
);

OR2x2_ASAP7_75t_L g4270 ( 
.A(n_4048),
.B(n_79),
.Y(n_4270)
);

OAI21x1_ASAP7_75t_L g4271 ( 
.A1(n_4132),
.A2(n_1899),
.B(n_1889),
.Y(n_4271)
);

AOI22xp33_ASAP7_75t_L g4272 ( 
.A1(n_4046),
.A2(n_4158),
.B1(n_4174),
.B2(n_4064),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4069),
.Y(n_4273)
);

AO21x2_ASAP7_75t_L g4274 ( 
.A1(n_4043),
.A2(n_83),
.B(n_84),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_4072),
.B(n_84),
.Y(n_4275)
);

OAI21x1_ASAP7_75t_L g4276 ( 
.A1(n_4120),
.A2(n_1906),
.B(n_1899),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4086),
.Y(n_4277)
);

OA21x2_ASAP7_75t_L g4278 ( 
.A1(n_4204),
.A2(n_85),
.B(n_86),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4078),
.Y(n_4279)
);

O2A1O1Ixp33_ASAP7_75t_SL g4280 ( 
.A1(n_4181),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_4080),
.B(n_88),
.Y(n_4281)
);

OAI21x1_ASAP7_75t_SL g4282 ( 
.A1(n_4219),
.A2(n_88),
.B(n_90),
.Y(n_4282)
);

AOI22xp5_ASAP7_75t_L g4283 ( 
.A1(n_4125),
.A2(n_1811),
.B1(n_1831),
.B2(n_1830),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4164),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4099),
.Y(n_4285)
);

AOI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4063),
.A2(n_1811),
.B1(n_1831),
.B2(n_1830),
.Y(n_4286)
);

AOI22xp33_ASAP7_75t_SL g4287 ( 
.A1(n_4119),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_4287)
);

AOI221xp5_ASAP7_75t_L g4288 ( 
.A1(n_4045),
.A2(n_1832),
.B1(n_1831),
.B2(n_1845),
.C(n_96),
.Y(n_4288)
);

NAND3x1_ASAP7_75t_L g4289 ( 
.A(n_4025),
.B(n_94),
.C(n_95),
.Y(n_4289)
);

OAI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_4222),
.A2(n_1832),
.B1(n_1831),
.B2(n_98),
.Y(n_4290)
);

INVx1_ASAP7_75t_SL g4291 ( 
.A(n_4227),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4091),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4112),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4102),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4166),
.B(n_95),
.Y(n_4295)
);

AOI22xp33_ASAP7_75t_L g4296 ( 
.A1(n_4119),
.A2(n_1832),
.B1(n_2916),
.B2(n_1518),
.Y(n_4296)
);

CKINVDCx5p33_ASAP7_75t_R g4297 ( 
.A(n_4021),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4161),
.B(n_97),
.Y(n_4298)
);

AOI22xp33_ASAP7_75t_L g4299 ( 
.A1(n_4130),
.A2(n_4030),
.B1(n_4123),
.B2(n_4028),
.Y(n_4299)
);

AND2x2_ASAP7_75t_L g4300 ( 
.A(n_4040),
.B(n_101),
.Y(n_4300)
);

CKINVDCx20_ASAP7_75t_R g4301 ( 
.A(n_4042),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4116),
.Y(n_4302)
);

AOI22xp33_ASAP7_75t_SL g4303 ( 
.A1(n_4175),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_4303)
);

OAI21x1_ASAP7_75t_L g4304 ( 
.A1(n_4075),
.A2(n_1921),
.B(n_1906),
.Y(n_4304)
);

OAI22xp5_ASAP7_75t_L g4305 ( 
.A1(n_4191),
.A2(n_1832),
.B1(n_107),
.B2(n_103),
.Y(n_4305)
);

AOI22xp33_ASAP7_75t_L g4306 ( 
.A1(n_4177),
.A2(n_1635),
.B1(n_1875),
.B2(n_1867),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4114),
.Y(n_4307)
);

O2A1O1Ixp33_ASAP7_75t_SL g4308 ( 
.A1(n_4202),
.A2(n_111),
.B(n_105),
.C(n_109),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4020),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4168),
.Y(n_4310)
);

BUFx12f_ASAP7_75t_SL g4311 ( 
.A(n_4089),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4134),
.Y(n_4312)
);

O2A1O1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_4160),
.A2(n_115),
.B(n_109),
.C(n_111),
.Y(n_4313)
);

AOI22xp33_ASAP7_75t_L g4314 ( 
.A1(n_4182),
.A2(n_1635),
.B1(n_1875),
.B2(n_1867),
.Y(n_4314)
);

OAI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4236),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_4315)
);

AOI22xp33_ASAP7_75t_L g4316 ( 
.A1(n_4039),
.A2(n_4179),
.B1(n_4101),
.B2(n_4024),
.Y(n_4316)
);

OAI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_4237),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_4317)
);

AO31x2_ASAP7_75t_L g4318 ( 
.A1(n_4196),
.A2(n_120),
.A3(n_118),
.B(n_119),
.Y(n_4318)
);

AOI22xp33_ASAP7_75t_SL g4319 ( 
.A1(n_4247),
.A2(n_124),
.B1(n_120),
.B2(n_121),
.Y(n_4319)
);

NAND2x1_ASAP7_75t_L g4320 ( 
.A(n_4215),
.B(n_1539),
.Y(n_4320)
);

INVx4_ASAP7_75t_SL g4321 ( 
.A(n_4199),
.Y(n_4321)
);

INVx6_ASAP7_75t_L g4322 ( 
.A(n_4100),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4137),
.Y(n_4323)
);

AOI22xp33_ASAP7_75t_L g4324 ( 
.A1(n_4186),
.A2(n_1635),
.B1(n_1876),
.B2(n_1875),
.Y(n_4324)
);

AND2x4_ASAP7_75t_L g4325 ( 
.A(n_4234),
.B(n_124),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4155),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4157),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4128),
.B(n_126),
.Y(n_4328)
);

OAI22xp5_ASAP7_75t_L g4329 ( 
.A1(n_4019),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_4329)
);

OAI221xp5_ASAP7_75t_L g4330 ( 
.A1(n_4018),
.A2(n_133),
.B1(n_128),
.B2(n_132),
.C(n_135),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4136),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_4159),
.B(n_132),
.Y(n_4332)
);

BUFx2_ASAP7_75t_L g4333 ( 
.A(n_4188),
.Y(n_4333)
);

AOI22xp33_ASAP7_75t_L g4334 ( 
.A1(n_4207),
.A2(n_1635),
.B1(n_1877),
.B2(n_1876),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4093),
.B(n_133),
.Y(n_4335)
);

CKINVDCx20_ASAP7_75t_R g4336 ( 
.A(n_4050),
.Y(n_4336)
);

INVx3_ASAP7_75t_L g4337 ( 
.A(n_4165),
.Y(n_4337)
);

AOI22xp33_ASAP7_75t_SL g4338 ( 
.A1(n_4052),
.A2(n_139),
.B1(n_136),
.B2(n_138),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4115),
.B(n_136),
.Y(n_4339)
);

A2O1A1Ixp33_ASAP7_75t_L g4340 ( 
.A1(n_4238),
.A2(n_141),
.B(n_138),
.C(n_140),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4136),
.Y(n_4341)
);

AOI21x1_ASAP7_75t_L g4342 ( 
.A1(n_4074),
.A2(n_140),
.B(n_142),
.Y(n_4342)
);

O2A1O1Ixp33_ASAP7_75t_L g4343 ( 
.A1(n_4088),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4136),
.Y(n_4344)
);

OR2x6_ASAP7_75t_L g4345 ( 
.A(n_4241),
.B(n_1876),
.Y(n_4345)
);

AOI21xp5_ASAP7_75t_L g4346 ( 
.A1(n_4029),
.A2(n_1921),
.B(n_1906),
.Y(n_4346)
);

AND2x4_ASAP7_75t_L g4347 ( 
.A(n_4239),
.B(n_145),
.Y(n_4347)
);

BUFx12f_ASAP7_75t_L g4348 ( 
.A(n_4027),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4190),
.Y(n_4349)
);

AOI22xp33_ASAP7_75t_L g4350 ( 
.A1(n_4067),
.A2(n_1635),
.B1(n_1877),
.B2(n_1876),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4066),
.Y(n_4351)
);

CKINVDCx11_ASAP7_75t_R g4352 ( 
.A(n_4197),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4066),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4066),
.B(n_146),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4218),
.B(n_146),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4066),
.Y(n_4356)
);

OAI21x1_ASAP7_75t_L g4357 ( 
.A1(n_4060),
.A2(n_1942),
.B(n_1921),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4103),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4170),
.B(n_147),
.Y(n_4359)
);

OAI221xp5_ASAP7_75t_L g4360 ( 
.A1(n_4062),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.C(n_152),
.Y(n_4360)
);

OAI22xp33_ASAP7_75t_L g4361 ( 
.A1(n_4145),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4113),
.B(n_153),
.Y(n_4362)
);

INVx6_ASAP7_75t_L g4363 ( 
.A(n_4096),
.Y(n_4363)
);

OAI22xp5_ASAP7_75t_L g4364 ( 
.A1(n_4235),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_4053),
.B(n_156),
.Y(n_4365)
);

OAI22xp5_ASAP7_75t_L g4366 ( 
.A1(n_4068),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4366)
);

AND2x4_ASAP7_75t_L g4367 ( 
.A(n_4217),
.B(n_157),
.Y(n_4367)
);

AOI22xp33_ASAP7_75t_SL g4368 ( 
.A1(n_4090),
.A2(n_161),
.B1(n_158),
.B2(n_160),
.Y(n_4368)
);

OAI22xp5_ASAP7_75t_L g4369 ( 
.A1(n_4073),
.A2(n_163),
.B1(n_160),
.B2(n_161),
.Y(n_4369)
);

AOI22xp33_ASAP7_75t_L g4370 ( 
.A1(n_4142),
.A2(n_1635),
.B1(n_1890),
.B2(n_1877),
.Y(n_4370)
);

A2O1A1Ixp33_ASAP7_75t_L g4371 ( 
.A1(n_4094),
.A2(n_167),
.B(n_164),
.C(n_166),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_L g4372 ( 
.A1(n_4104),
.A2(n_1890),
.B1(n_1898),
.B2(n_1877),
.Y(n_4372)
);

INVx1_ASAP7_75t_SL g4373 ( 
.A(n_4031),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4117),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4103),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_4225),
.B(n_164),
.Y(n_4376)
);

INVx2_ASAP7_75t_SL g4377 ( 
.A(n_4241),
.Y(n_4377)
);

AOI22xp33_ASAP7_75t_L g4378 ( 
.A1(n_4111),
.A2(n_1898),
.B1(n_1922),
.B2(n_1890),
.Y(n_4378)
);

OAI22xp5_ASAP7_75t_L g4379 ( 
.A1(n_4124),
.A2(n_169),
.B1(n_166),
.B2(n_168),
.Y(n_4379)
);

AOI22xp33_ASAP7_75t_SL g4380 ( 
.A1(n_4079),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4103),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4059),
.B(n_4087),
.Y(n_4382)
);

O2A1O1Ixp33_ASAP7_75t_L g4383 ( 
.A1(n_4047),
.A2(n_178),
.B(n_176),
.C(n_177),
.Y(n_4383)
);

INVx3_ASAP7_75t_L g4384 ( 
.A(n_4201),
.Y(n_4384)
);

AOI22xp33_ASAP7_75t_L g4385 ( 
.A1(n_4098),
.A2(n_1898),
.B1(n_1922),
.B2(n_1890),
.Y(n_4385)
);

AND2x4_ASAP7_75t_L g4386 ( 
.A(n_4201),
.B(n_176),
.Y(n_4386)
);

NAND2xp33_ASAP7_75t_R g4387 ( 
.A(n_4249),
.B(n_177),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_L g4388 ( 
.A1(n_4176),
.A2(n_1922),
.B1(n_1924),
.B2(n_1898),
.Y(n_4388)
);

AOI222xp33_ASAP7_75t_L g4389 ( 
.A1(n_4049),
.A2(n_182),
.B1(n_184),
.B2(n_179),
.C1(n_181),
.C2(n_183),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4055),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_SL g4391 ( 
.A(n_4109),
.B(n_1539),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4037),
.Y(n_4392)
);

OR2x2_ASAP7_75t_L g4393 ( 
.A(n_4037),
.B(n_179),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_4096),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4037),
.Y(n_4395)
);

OAI21x1_ASAP7_75t_L g4396 ( 
.A1(n_4106),
.A2(n_1959),
.B(n_1942),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4097),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_L g4398 ( 
.A1(n_4220),
.A2(n_4077),
.B1(n_4143),
.B2(n_4032),
.Y(n_4398)
);

NAND3xp33_ASAP7_75t_L g4399 ( 
.A(n_4154),
.B(n_1560),
.C(n_1539),
.Y(n_4399)
);

OAI21x1_ASAP7_75t_SL g4400 ( 
.A1(n_4189),
.A2(n_183),
.B(n_184),
.Y(n_4400)
);

AND2x4_ASAP7_75t_L g4401 ( 
.A(n_4201),
.B(n_185),
.Y(n_4401)
);

AOI22xp33_ASAP7_75t_L g4402 ( 
.A1(n_4169),
.A2(n_1924),
.B1(n_1938),
.B2(n_1922),
.Y(n_4402)
);

OR2x2_ASAP7_75t_L g4403 ( 
.A(n_4097),
.B(n_4203),
.Y(n_4403)
);

AND2x4_ASAP7_75t_L g4404 ( 
.A(n_4141),
.B(n_185),
.Y(n_4404)
);

AOI222xp33_ASAP7_75t_L g4405 ( 
.A1(n_4205),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.C1(n_191),
.C2(n_193),
.Y(n_4405)
);

AOI22xp33_ASAP7_75t_L g4406 ( 
.A1(n_4208),
.A2(n_1938),
.B1(n_1939),
.B2(n_1924),
.Y(n_4406)
);

O2A1O1Ixp33_ASAP7_75t_SL g4407 ( 
.A1(n_4221),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_4407)
);

CKINVDCx5p33_ASAP7_75t_R g4408 ( 
.A(n_4107),
.Y(n_4408)
);

AOI22xp33_ASAP7_75t_L g4409 ( 
.A1(n_4206),
.A2(n_1938),
.B1(n_1939),
.B2(n_1924),
.Y(n_4409)
);

O2A1O1Ixp33_ASAP7_75t_SL g4410 ( 
.A1(n_4228),
.A2(n_196),
.B(n_193),
.C(n_195),
.Y(n_4410)
);

AOI222xp33_ASAP7_75t_L g4411 ( 
.A1(n_4151),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.C1(n_201),
.C2(n_203),
.Y(n_4411)
);

BUFx10_ASAP7_75t_L g4412 ( 
.A(n_4184),
.Y(n_4412)
);

INVx1_ASAP7_75t_SL g4413 ( 
.A(n_4127),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4097),
.Y(n_4414)
);

AO21x2_ASAP7_75t_L g4415 ( 
.A1(n_4034),
.A2(n_199),
.B(n_201),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4038),
.Y(n_4416)
);

AND2x4_ASAP7_75t_L g4417 ( 
.A(n_4230),
.B(n_4133),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4216),
.Y(n_4418)
);

BUFx2_ASAP7_75t_L g4419 ( 
.A(n_4140),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4243),
.A2(n_4171),
.B1(n_4187),
.B2(n_4193),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4240),
.Y(n_4421)
);

AOI221xp5_ASAP7_75t_L g4422 ( 
.A1(n_4083),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.C(n_207),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4244),
.B(n_204),
.Y(n_4423)
);

BUFx12f_ASAP7_75t_L g4424 ( 
.A(n_4232),
.Y(n_4424)
);

OA21x2_ASAP7_75t_L g4425 ( 
.A1(n_4149),
.A2(n_206),
.B(n_208),
.Y(n_4425)
);

OAI22x1_ASAP7_75t_L g4426 ( 
.A1(n_4240),
.A2(n_212),
.B1(n_209),
.B2(n_211),
.Y(n_4426)
);

AOI221xp5_ASAP7_75t_L g4427 ( 
.A1(n_4054),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4240),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4152),
.B(n_213),
.Y(n_4429)
);

INVx3_ASAP7_75t_L g4430 ( 
.A(n_4194),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4026),
.B(n_214),
.Y(n_4431)
);

AOI22xp33_ASAP7_75t_L g4432 ( 
.A1(n_4209),
.A2(n_1939),
.B1(n_1949),
.B2(n_1938),
.Y(n_4432)
);

O2A1O1Ixp33_ASAP7_75t_L g4433 ( 
.A1(n_4057),
.A2(n_4167),
.B(n_4212),
.C(n_4129),
.Y(n_4433)
);

AO31x2_ASAP7_75t_L g4434 ( 
.A1(n_4214),
.A2(n_218),
.A3(n_215),
.B(n_216),
.Y(n_4434)
);

INVx3_ASAP7_75t_L g4435 ( 
.A(n_4384),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4331),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4257),
.B(n_4038),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4333),
.B(n_4038),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4344),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_4322),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4341),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4263),
.Y(n_4442)
);

BUFx2_ASAP7_75t_L g4443 ( 
.A(n_4254),
.Y(n_4443)
);

INVx2_ASAP7_75t_L g4444 ( 
.A(n_4273),
.Y(n_4444)
);

INVx3_ASAP7_75t_L g4445 ( 
.A(n_4384),
.Y(n_4445)
);

AND2x4_ASAP7_75t_L g4446 ( 
.A(n_4254),
.B(n_4353),
.Y(n_4446)
);

AOI22xp33_ASAP7_75t_L g4447 ( 
.A1(n_4389),
.A2(n_4138),
.B1(n_4163),
.B2(n_4148),
.Y(n_4447)
);

AND2x2_ASAP7_75t_L g4448 ( 
.A(n_4390),
.B(n_4131),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_4279),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4292),
.Y(n_4450)
);

NAND2x1p5_ASAP7_75t_L g4451 ( 
.A(n_4386),
.B(n_4105),
.Y(n_4451)
);

BUFx3_ASAP7_75t_L g4452 ( 
.A(n_4322),
.Y(n_4452)
);

OR2x2_ASAP7_75t_L g4453 ( 
.A(n_4284),
.B(n_4131),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4293),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4302),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4261),
.B(n_4035),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4309),
.Y(n_4457)
);

NAND2xp33_ASAP7_75t_L g4458 ( 
.A(n_4289),
.B(n_4146),
.Y(n_4458)
);

HB1xp67_ASAP7_75t_L g4459 ( 
.A(n_4309),
.Y(n_4459)
);

HB1xp67_ASAP7_75t_L g4460 ( 
.A(n_4310),
.Y(n_4460)
);

INVx3_ASAP7_75t_L g4461 ( 
.A(n_4412),
.Y(n_4461)
);

INVx2_ASAP7_75t_L g4462 ( 
.A(n_4326),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4250),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4307),
.Y(n_4464)
);

OAI21x1_ASAP7_75t_L g4465 ( 
.A1(n_4397),
.A2(n_4110),
.B(n_4105),
.Y(n_4465)
);

BUFx2_ASAP7_75t_L g4466 ( 
.A(n_4424),
.Y(n_4466)
);

OAI21x1_ASAP7_75t_L g4467 ( 
.A1(n_4392),
.A2(n_4110),
.B(n_4226),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4312),
.Y(n_4468)
);

AO21x2_ASAP7_75t_L g4469 ( 
.A1(n_4395),
.A2(n_4414),
.B(n_4358),
.Y(n_4469)
);

INVx2_ASAP7_75t_L g4470 ( 
.A(n_4266),
.Y(n_4470)
);

OA21x2_ASAP7_75t_L g4471 ( 
.A1(n_4416),
.A2(n_4231),
.B(n_4172),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4323),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4327),
.Y(n_4473)
);

OAI21xp5_ASAP7_75t_L g4474 ( 
.A1(n_4272),
.A2(n_4041),
.B(n_4150),
.Y(n_4474)
);

INVx2_ASAP7_75t_SL g4475 ( 
.A(n_4412),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4277),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4285),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_4405),
.A2(n_4153),
.B1(n_4121),
.B2(n_4211),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_4294),
.Y(n_4479)
);

AO21x2_ASAP7_75t_L g4480 ( 
.A1(n_4358),
.A2(n_4416),
.B(n_4274),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4349),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4374),
.Y(n_4482)
);

OAI21x1_ASAP7_75t_L g4483 ( 
.A1(n_4276),
.A2(n_4195),
.B(n_4246),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4430),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4430),
.Y(n_4485)
);

INVx2_ASAP7_75t_SL g4486 ( 
.A(n_4419),
.Y(n_4486)
);

OA21x2_ASAP7_75t_L g4487 ( 
.A1(n_4375),
.A2(n_4108),
.B(n_4183),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4403),
.Y(n_4488)
);

OAI21x1_ASAP7_75t_L g4489 ( 
.A1(n_4271),
.A2(n_4210),
.B(n_4200),
.Y(n_4489)
);

INVx3_ASAP7_75t_L g4490 ( 
.A(n_4386),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4393),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4421),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4351),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4428),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4356),
.Y(n_4495)
);

INVx3_ASAP7_75t_L g4496 ( 
.A(n_4401),
.Y(n_4496)
);

HB1xp67_ASAP7_75t_L g4497 ( 
.A(n_4278),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4278),
.Y(n_4498)
);

OAI22xp5_ASAP7_75t_L g4499 ( 
.A1(n_4340),
.A2(n_4192),
.B1(n_4198),
.B2(n_4229),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4381),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4418),
.Y(n_4501)
);

OR2x2_ASAP7_75t_L g4502 ( 
.A(n_4258),
.B(n_4131),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4269),
.B(n_4122),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4415),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4265),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4337),
.B(n_4122),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4268),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4268),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4268),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4270),
.Y(n_4510)
);

INVx2_ASAP7_75t_SL g4511 ( 
.A(n_4417),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_4415),
.Y(n_4512)
);

BUFx3_ASAP7_75t_L g4513 ( 
.A(n_4256),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4328),
.Y(n_4514)
);

OA21x2_ASAP7_75t_L g4515 ( 
.A1(n_4354),
.A2(n_4223),
.B(n_4118),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4337),
.B(n_4122),
.Y(n_4516)
);

BUFx2_ASAP7_75t_L g4517 ( 
.A(n_4255),
.Y(n_4517)
);

INVxp67_ASAP7_75t_L g4518 ( 
.A(n_4387),
.Y(n_4518)
);

INVx1_ASAP7_75t_SL g4519 ( 
.A(n_4352),
.Y(n_4519)
);

OR2x2_ASAP7_75t_L g4520 ( 
.A(n_4373),
.B(n_4413),
.Y(n_4520)
);

BUFx6f_ASAP7_75t_L g4521 ( 
.A(n_4401),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4274),
.Y(n_4522)
);

OA21x2_ASAP7_75t_L g4523 ( 
.A1(n_4431),
.A2(n_4147),
.B(n_4144),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4332),
.Y(n_4524)
);

HB1xp67_ASAP7_75t_L g4525 ( 
.A(n_4434),
.Y(n_4525)
);

OR2x6_ASAP7_75t_L g4526 ( 
.A(n_4260),
.B(n_4245),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4291),
.B(n_4139),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4434),
.Y(n_4528)
);

BUFx2_ASAP7_75t_R g4529 ( 
.A(n_4297),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4434),
.Y(n_4530)
);

BUFx2_ASAP7_75t_L g4531 ( 
.A(n_4417),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_4363),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4318),
.Y(n_4533)
);

AO21x2_ASAP7_75t_L g4534 ( 
.A1(n_4282),
.A2(n_4248),
.B(n_4070),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4298),
.Y(n_4535)
);

NAND3xp33_ASAP7_75t_L g4536 ( 
.A(n_4299),
.B(n_4084),
.C(n_4233),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_4318),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4318),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4429),
.Y(n_4539)
);

INVx2_ASAP7_75t_L g4540 ( 
.A(n_4320),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4281),
.Y(n_4541)
);

OA21x2_ASAP7_75t_L g4542 ( 
.A1(n_4396),
.A2(n_4153),
.B(n_4082),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4281),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4252),
.B(n_4139),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4362),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4342),
.Y(n_4546)
);

OR2x2_ASAP7_75t_L g4547 ( 
.A(n_4339),
.B(n_4139),
.Y(n_4547)
);

AO31x2_ASAP7_75t_L g4548 ( 
.A1(n_4426),
.A2(n_4153),
.A3(n_4173),
.B(n_4180),
.Y(n_4548)
);

AND2x4_ASAP7_75t_L g4549 ( 
.A(n_4325),
.B(n_4173),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4325),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4347),
.Y(n_4551)
);

CKINVDCx16_ASAP7_75t_R g4552 ( 
.A(n_4348),
.Y(n_4552)
);

CKINVDCx20_ASAP7_75t_R g4553 ( 
.A(n_4301),
.Y(n_4553)
);

INVx5_ASAP7_75t_L g4554 ( 
.A(n_4256),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4347),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4367),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_4363),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4336),
.Y(n_4558)
);

CKINVDCx5p33_ASAP7_75t_R g4559 ( 
.A(n_4394),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4425),
.Y(n_4560)
);

INVx3_ASAP7_75t_L g4561 ( 
.A(n_4367),
.Y(n_4561)
);

AND2x4_ASAP7_75t_L g4562 ( 
.A(n_4321),
.B(n_4173),
.Y(n_4562)
);

HB1xp67_ASAP7_75t_L g4563 ( 
.A(n_4425),
.Y(n_4563)
);

AO21x1_ASAP7_75t_L g4564 ( 
.A1(n_4343),
.A2(n_4224),
.B(n_4185),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4376),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4423),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4376),
.Y(n_4567)
);

OAI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4313),
.A2(n_4056),
.B(n_4156),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4295),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4304),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4357),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4400),
.Y(n_4572)
);

INVx2_ASAP7_75t_L g4573 ( 
.A(n_4404),
.Y(n_4573)
);

AOI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4564),
.A2(n_4360),
.B1(n_4380),
.B2(n_4411),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4501),
.Y(n_4575)
);

AOI221xp5_ASAP7_75t_L g4576 ( 
.A1(n_4497),
.A2(n_4280),
.B1(n_4383),
.B2(n_4329),
.C(n_4407),
.Y(n_4576)
);

AOI21xp5_ASAP7_75t_L g4577 ( 
.A1(n_4474),
.A2(n_4259),
.B(n_4433),
.Y(n_4577)
);

A2O1A1Ixp33_ASAP7_75t_L g4578 ( 
.A1(n_4458),
.A2(n_4422),
.B(n_4427),
.C(n_4303),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4459),
.Y(n_4579)
);

AND2x2_ASAP7_75t_L g4580 ( 
.A(n_4443),
.B(n_4267),
.Y(n_4580)
);

OAI22xp5_ASAP7_75t_L g4581 ( 
.A1(n_4478),
.A2(n_4287),
.B1(n_4420),
.B2(n_4251),
.Y(n_4581)
);

AOI21xp33_ASAP7_75t_L g4582 ( 
.A1(n_4456),
.A2(n_4253),
.B(n_4382),
.Y(n_4582)
);

AOI221xp5_ASAP7_75t_L g4583 ( 
.A1(n_4497),
.A2(n_4410),
.B1(n_4330),
.B2(n_4317),
.C(n_4315),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4459),
.Y(n_4584)
);

NAND2x1_ASAP7_75t_L g4585 ( 
.A(n_4490),
.B(n_4404),
.Y(n_4585)
);

OAI22xp5_ASAP7_75t_L g4586 ( 
.A1(n_4478),
.A2(n_4399),
.B1(n_4264),
.B2(n_4398),
.Y(n_4586)
);

NOR2xp33_ASAP7_75t_L g4587 ( 
.A(n_4519),
.B(n_4311),
.Y(n_4587)
);

AOI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4456),
.A2(n_4364),
.B1(n_4305),
.B2(n_4366),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4444),
.Y(n_4589)
);

BUFx2_ASAP7_75t_L g4590 ( 
.A(n_4490),
.Y(n_4590)
);

AOI22xp5_ASAP7_75t_L g4591 ( 
.A1(n_4458),
.A2(n_4319),
.B1(n_4369),
.B2(n_4288),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4490),
.Y(n_4592)
);

OAI211xp5_ASAP7_75t_SL g4593 ( 
.A1(n_4572),
.A2(n_4491),
.B(n_4518),
.C(n_4535),
.Y(n_4593)
);

INVx2_ASAP7_75t_SL g4594 ( 
.A(n_4513),
.Y(n_4594)
);

HB1xp67_ASAP7_75t_L g4595 ( 
.A(n_4460),
.Y(n_4595)
);

OAI211xp5_ASAP7_75t_L g4596 ( 
.A1(n_4525),
.A2(n_4368),
.B(n_4371),
.C(n_4338),
.Y(n_4596)
);

AO21x2_ASAP7_75t_L g4597 ( 
.A1(n_4522),
.A2(n_4359),
.B(n_4308),
.Y(n_4597)
);

AOI22xp33_ASAP7_75t_SL g4598 ( 
.A1(n_4536),
.A2(n_4275),
.B1(n_4290),
.B2(n_4379),
.Y(n_4598)
);

AOI22xp33_ASAP7_75t_L g4599 ( 
.A1(n_4572),
.A2(n_4316),
.B1(n_4361),
.B2(n_4391),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4531),
.B(n_4321),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4496),
.B(n_4408),
.Y(n_4601)
);

AOI221xp5_ASAP7_75t_L g4602 ( 
.A1(n_4498),
.A2(n_4365),
.B1(n_4300),
.B2(n_4355),
.C(n_4335),
.Y(n_4602)
);

AOI22xp33_ASAP7_75t_L g4603 ( 
.A1(n_4539),
.A2(n_4286),
.B1(n_4385),
.B2(n_4314),
.Y(n_4603)
);

OAI221xp5_ASAP7_75t_L g4604 ( 
.A1(n_4514),
.A2(n_4524),
.B1(n_4545),
.B2(n_4568),
.C(n_4525),
.Y(n_4604)
);

AOI22xp33_ASAP7_75t_L g4605 ( 
.A1(n_4539),
.A2(n_4324),
.B1(n_4409),
.B2(n_4296),
.Y(n_4605)
);

OAI22xp33_ASAP7_75t_L g4606 ( 
.A1(n_4526),
.A2(n_4283),
.B1(n_4262),
.B2(n_4377),
.Y(n_4606)
);

AOI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_4499),
.A2(n_4406),
.B(n_4378),
.Y(n_4607)
);

BUFx2_ASAP7_75t_L g4608 ( 
.A(n_4496),
.Y(n_4608)
);

AND2x4_ASAP7_75t_L g4609 ( 
.A(n_4562),
.B(n_4345),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_4460),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4496),
.Y(n_4611)
);

INVx3_ASAP7_75t_L g4612 ( 
.A(n_4521),
.Y(n_4612)
);

OAI22xp33_ASAP7_75t_L g4613 ( 
.A1(n_4526),
.A2(n_4345),
.B1(n_4162),
.B2(n_4121),
.Y(n_4613)
);

OAI22xp5_ASAP7_75t_L g4614 ( 
.A1(n_4554),
.A2(n_4402),
.B1(n_4388),
.B2(n_4432),
.Y(n_4614)
);

AOI221xp5_ASAP7_75t_L g4615 ( 
.A1(n_4522),
.A2(n_4372),
.B1(n_4346),
.B2(n_4334),
.C(n_4350),
.Y(n_4615)
);

AND2x4_ASAP7_75t_L g4616 ( 
.A(n_4562),
.B(n_4554),
.Y(n_4616)
);

OAI22xp5_ASAP7_75t_L g4617 ( 
.A1(n_4554),
.A2(n_4370),
.B1(n_4306),
.B2(n_4242),
.Y(n_4617)
);

OAI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4554),
.A2(n_4526),
.B1(n_4447),
.B2(n_4521),
.Y(n_4618)
);

OAI211xp5_ASAP7_75t_SL g4619 ( 
.A1(n_4510),
.A2(n_220),
.B(n_216),
.C(n_219),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4527),
.B(n_4180),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4503),
.B(n_4180),
.Y(n_4621)
);

AOI221xp5_ASAP7_75t_L g4622 ( 
.A1(n_4546),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.C(n_225),
.Y(n_4622)
);

AOI22xp33_ASAP7_75t_L g4623 ( 
.A1(n_4534),
.A2(n_1949),
.B1(n_1939),
.B2(n_1942),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4444),
.Y(n_4624)
);

OAI222xp33_ASAP7_75t_L g4625 ( 
.A1(n_4506),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.C1(n_226),
.C2(n_227),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4493),
.Y(n_4626)
);

INVx5_ASAP7_75t_L g4627 ( 
.A(n_4552),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4493),
.Y(n_4628)
);

AOI22xp5_ASAP7_75t_L g4629 ( 
.A1(n_4447),
.A2(n_230),
.B1(n_226),
.B2(n_229),
.Y(n_4629)
);

OAI22xp33_ASAP7_75t_L g4630 ( 
.A1(n_4521),
.A2(n_4213),
.B1(n_232),
.B2(n_229),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4449),
.Y(n_4631)
);

NAND3xp33_ASAP7_75t_L g4632 ( 
.A(n_4546),
.B(n_231),
.C(n_233),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4516),
.B(n_4213),
.Y(n_4633)
);

OA21x2_ASAP7_75t_L g4634 ( 
.A1(n_4436),
.A2(n_4213),
.B(n_231),
.Y(n_4634)
);

OAI22x1_ASAP7_75t_L g4635 ( 
.A1(n_4541),
.A2(n_4543),
.B1(n_4555),
.B2(n_4550),
.Y(n_4635)
);

OAI22xp5_ASAP7_75t_L g4636 ( 
.A1(n_4521),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4449),
.Y(n_4637)
);

AOI222xp33_ASAP7_75t_L g4638 ( 
.A1(n_4505),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.C1(n_238),
.C2(n_239),
.Y(n_4638)
);

AND2x2_ASAP7_75t_L g4639 ( 
.A(n_4511),
.B(n_236),
.Y(n_4639)
);

OAI22xp5_ASAP7_75t_L g4640 ( 
.A1(n_4550),
.A2(n_4555),
.B1(n_4561),
.B2(n_4551),
.Y(n_4640)
);

AOI222xp33_ASAP7_75t_L g4641 ( 
.A1(n_4507),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.C1(n_243),
.C2(n_244),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4511),
.B(n_4517),
.Y(n_4642)
);

AOI22xp33_ASAP7_75t_L g4643 ( 
.A1(n_4534),
.A2(n_1949),
.B1(n_1970),
.B2(n_1959),
.Y(n_4643)
);

AOI22xp33_ASAP7_75t_L g4644 ( 
.A1(n_4561),
.A2(n_1949),
.B1(n_1970),
.B2(n_1959),
.Y(n_4644)
);

OAI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4561),
.A2(n_249),
.B1(n_245),
.B2(n_247),
.Y(n_4645)
);

A2O1A1Ixp33_ASAP7_75t_L g4646 ( 
.A1(n_4538),
.A2(n_251),
.B(n_247),
.C(n_250),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_4553),
.Y(n_4647)
);

OAI22xp5_ASAP7_75t_L g4648 ( 
.A1(n_4573),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4486),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4479),
.Y(n_4650)
);

OAI21x1_ASAP7_75t_L g4651 ( 
.A1(n_4435),
.A2(n_1567),
.B(n_1560),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4450),
.Y(n_4652)
);

OAI322xp33_ASAP7_75t_L g4653 ( 
.A1(n_4530),
.A2(n_253),
.A3(n_254),
.B1(n_256),
.B2(n_257),
.C1(n_258),
.C2(n_259),
.Y(n_4653)
);

OAI221xp5_ASAP7_75t_SL g4654 ( 
.A1(n_4504),
.A2(n_253),
.B1(n_254),
.B2(n_258),
.C(n_259),
.Y(n_4654)
);

AOI22xp33_ASAP7_75t_SL g4655 ( 
.A1(n_4466),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_4655)
);

AOI22xp33_ASAP7_75t_L g4656 ( 
.A1(n_4566),
.A2(n_1978),
.B1(n_1986),
.B2(n_1970),
.Y(n_4656)
);

AOI22xp33_ASAP7_75t_L g4657 ( 
.A1(n_4566),
.A2(n_1986),
.B1(n_2001),
.B2(n_1978),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4450),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4486),
.B(n_261),
.Y(n_4659)
);

OAI22xp33_ASAP7_75t_L g4660 ( 
.A1(n_4547),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_4660)
);

OAI22xp5_ASAP7_75t_L g4661 ( 
.A1(n_4573),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_4661)
);

OAI221xp5_ASAP7_75t_L g4662 ( 
.A1(n_4508),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.C(n_268),
.Y(n_4662)
);

OR2x2_ASAP7_75t_L g4663 ( 
.A(n_4488),
.B(n_267),
.Y(n_4663)
);

OAI22xp5_ASAP7_75t_L g4664 ( 
.A1(n_4556),
.A2(n_272),
.B1(n_268),
.B2(n_271),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_4513),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4454),
.Y(n_4666)
);

AOI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_4562),
.A2(n_271),
.B(n_272),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4454),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4446),
.B(n_274),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4455),
.Y(n_4670)
);

AO31x2_ASAP7_75t_L g4671 ( 
.A1(n_4504),
.A2(n_277),
.A3(n_274),
.B(n_276),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4512),
.A2(n_276),
.B(n_277),
.Y(n_4672)
);

AOI22xp33_ASAP7_75t_L g4673 ( 
.A1(n_4565),
.A2(n_1986),
.B1(n_2001),
.B2(n_1978),
.Y(n_4673)
);

AOI22xp33_ASAP7_75t_L g4674 ( 
.A1(n_4567),
.A2(n_2004),
.B1(n_2011),
.B2(n_2001),
.Y(n_4674)
);

AOI222xp33_ASAP7_75t_L g4675 ( 
.A1(n_4509),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.C1(n_282),
.C2(n_285),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4455),
.Y(n_4676)
);

AOI22xp33_ASAP7_75t_SL g4677 ( 
.A1(n_4563),
.A2(n_289),
.B1(n_282),
.B2(n_288),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4512),
.A2(n_288),
.B(n_289),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4457),
.Y(n_4679)
);

AND2x4_ASAP7_75t_L g4680 ( 
.A(n_4461),
.B(n_290),
.Y(n_4680)
);

AOI22xp33_ASAP7_75t_L g4681 ( 
.A1(n_4569),
.A2(n_2011),
.B1(n_2035),
.B2(n_2004),
.Y(n_4681)
);

OAI22xp5_ASAP7_75t_L g4682 ( 
.A1(n_4475),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4544),
.B(n_291),
.Y(n_4683)
);

OAI21x1_ASAP7_75t_L g4684 ( 
.A1(n_4435),
.A2(n_1567),
.B(n_1560),
.Y(n_4684)
);

AOI22xp33_ASAP7_75t_L g4685 ( 
.A1(n_4440),
.A2(n_4452),
.B1(n_4448),
.B2(n_4549),
.Y(n_4685)
);

AND2x2_ASAP7_75t_L g4686 ( 
.A(n_4446),
.B(n_293),
.Y(n_4686)
);

INVxp67_ASAP7_75t_L g4687 ( 
.A(n_4482),
.Y(n_4687)
);

AOI22xp33_ASAP7_75t_L g4688 ( 
.A1(n_4440),
.A2(n_4452),
.B1(n_4549),
.B2(n_4523),
.Y(n_4688)
);

AOI22xp33_ASAP7_75t_SL g4689 ( 
.A1(n_4563),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_4689)
);

AOI22xp33_ASAP7_75t_L g4690 ( 
.A1(n_4549),
.A2(n_2004),
.B1(n_2035),
.B2(n_2011),
.Y(n_4690)
);

AOI22xp33_ASAP7_75t_L g4691 ( 
.A1(n_4523),
.A2(n_2035),
.B1(n_2112),
.B2(n_2085),
.Y(n_4691)
);

AOI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4523),
.A2(n_2085),
.B1(n_2141),
.B2(n_2112),
.Y(n_4692)
);

BUFx12f_ASAP7_75t_L g4693 ( 
.A(n_4558),
.Y(n_4693)
);

INVx3_ASAP7_75t_L g4694 ( 
.A(n_4446),
.Y(n_4694)
);

BUFx12f_ASAP7_75t_L g4695 ( 
.A(n_4558),
.Y(n_4695)
);

AOI22xp33_ASAP7_75t_L g4696 ( 
.A1(n_4533),
.A2(n_2085),
.B1(n_2141),
.B2(n_2112),
.Y(n_4696)
);

OAI21x1_ASAP7_75t_L g4697 ( 
.A1(n_4435),
.A2(n_1567),
.B(n_294),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4462),
.Y(n_4698)
);

AO21x2_ASAP7_75t_L g4699 ( 
.A1(n_4560),
.A2(n_297),
.B(n_298),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4442),
.Y(n_4700)
);

AOI22xp33_ASAP7_75t_L g4701 ( 
.A1(n_4533),
.A2(n_2158),
.B1(n_2181),
.B2(n_2141),
.Y(n_4701)
);

AOI22xp33_ASAP7_75t_L g4702 ( 
.A1(n_4537),
.A2(n_2181),
.B1(n_2158),
.B2(n_1984),
.Y(n_4702)
);

AOI22xp5_ASAP7_75t_L g4703 ( 
.A1(n_4553),
.A2(n_301),
.B1(n_297),
.B2(n_300),
.Y(n_4703)
);

OR2x6_ASAP7_75t_L g4704 ( 
.A(n_4528),
.B(n_300),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4464),
.B(n_302),
.Y(n_4705)
);

HB1xp67_ASAP7_75t_L g4706 ( 
.A(n_4595),
.Y(n_4706)
);

INVxp67_ASAP7_75t_L g4707 ( 
.A(n_4597),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4575),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4683),
.B(n_4437),
.Y(n_4709)
);

OR2x2_ASAP7_75t_L g4710 ( 
.A(n_4621),
.B(n_4492),
.Y(n_4710)
);

BUFx3_ASAP7_75t_L g4711 ( 
.A(n_4627),
.Y(n_4711)
);

INVx2_ASAP7_75t_L g4712 ( 
.A(n_4666),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4700),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4670),
.Y(n_4714)
);

OR2x2_ASAP7_75t_SL g4715 ( 
.A(n_4632),
.B(n_4529),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4616),
.B(n_4475),
.Y(n_4716)
);

INVx3_ASAP7_75t_L g4717 ( 
.A(n_4616),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4687),
.B(n_4468),
.Y(n_4718)
);

AND2x2_ASAP7_75t_L g4719 ( 
.A(n_4694),
.B(n_4461),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4626),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4694),
.B(n_4461),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4590),
.B(n_4494),
.Y(n_4722)
);

INVx1_ASAP7_75t_L g4723 ( 
.A(n_4679),
.Y(n_4723)
);

BUFx6f_ASAP7_75t_L g4724 ( 
.A(n_4627),
.Y(n_4724)
);

AND2x4_ASAP7_75t_L g4725 ( 
.A(n_4608),
.B(n_4540),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4628),
.Y(n_4726)
);

INVx4_ASAP7_75t_L g4727 ( 
.A(n_4627),
.Y(n_4727)
);

AND2x4_ASAP7_75t_L g4728 ( 
.A(n_4592),
.B(n_4540),
.Y(n_4728)
);

BUFx2_ASAP7_75t_L g4729 ( 
.A(n_4649),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4698),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4659),
.B(n_4472),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4611),
.B(n_4557),
.Y(n_4732)
);

OAI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_4577),
.A2(n_4537),
.B(n_4528),
.Y(n_4733)
);

HB1xp67_ASAP7_75t_L g4734 ( 
.A(n_4610),
.Y(n_4734)
);

AO211x2_ASAP7_75t_L g4735 ( 
.A1(n_4672),
.A2(n_4484),
.B(n_4485),
.C(n_4500),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4589),
.Y(n_4736)
);

BUFx6f_ASAP7_75t_L g4737 ( 
.A(n_4665),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4579),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4705),
.B(n_4473),
.Y(n_4739)
);

INVx2_ASAP7_75t_L g4740 ( 
.A(n_4624),
.Y(n_4740)
);

AOI22xp33_ASAP7_75t_L g4741 ( 
.A1(n_4574),
.A2(n_4515),
.B1(n_4520),
.B2(n_4557),
.Y(n_4741)
);

AND2x4_ASAP7_75t_L g4742 ( 
.A(n_4612),
.B(n_4445),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4584),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4612),
.B(n_4557),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4620),
.B(n_4685),
.Y(n_4745)
);

BUFx2_ASAP7_75t_L g4746 ( 
.A(n_4704),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4631),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4642),
.B(n_4532),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4637),
.Y(n_4749)
);

INVx2_ASAP7_75t_L g4750 ( 
.A(n_4652),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4600),
.B(n_4532),
.Y(n_4751)
);

BUFx3_ASAP7_75t_L g4752 ( 
.A(n_4693),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4658),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4668),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4688),
.B(n_4479),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4601),
.B(n_4495),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4676),
.Y(n_4757)
);

INVx1_ASAP7_75t_SL g4758 ( 
.A(n_4695),
.Y(n_4758)
);

NOR2xp33_ASAP7_75t_L g4759 ( 
.A(n_4582),
.B(n_4559),
.Y(n_4759)
);

BUFx3_ASAP7_75t_L g4760 ( 
.A(n_4665),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4650),
.Y(n_4761)
);

BUFx2_ASAP7_75t_L g4762 ( 
.A(n_4704),
.Y(n_4762)
);

AO21x2_ASAP7_75t_L g4763 ( 
.A1(n_4678),
.A2(n_4560),
.B(n_4439),
.Y(n_4763)
);

INVx3_ASAP7_75t_L g4764 ( 
.A(n_4609),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4671),
.Y(n_4765)
);

AND2x4_ASAP7_75t_SL g4766 ( 
.A(n_4665),
.B(n_4580),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4671),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4635),
.Y(n_4768)
);

AND2x2_ASAP7_75t_L g4769 ( 
.A(n_4609),
.B(n_4594),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4704),
.Y(n_4770)
);

HB1xp67_ASAP7_75t_L g4771 ( 
.A(n_4597),
.Y(n_4771)
);

AND2x2_ASAP7_75t_L g4772 ( 
.A(n_4640),
.B(n_4438),
.Y(n_4772)
);

OAI22xp5_ASAP7_75t_L g4773 ( 
.A1(n_4591),
.A2(n_4578),
.B1(n_4588),
.B2(n_4586),
.Y(n_4773)
);

AOI22xp33_ASAP7_75t_L g4774 ( 
.A1(n_4618),
.A2(n_4515),
.B1(n_4542),
.B2(n_4502),
.Y(n_4774)
);

OR2x2_ASAP7_75t_L g4775 ( 
.A(n_4633),
.B(n_4453),
.Y(n_4775)
);

OR2x2_ASAP7_75t_L g4776 ( 
.A(n_4663),
.B(n_4463),
.Y(n_4776)
);

INVx2_ASAP7_75t_SL g4777 ( 
.A(n_4585),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4671),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_L g4779 ( 
.A(n_4669),
.B(n_4476),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4699),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4699),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4686),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4639),
.B(n_4463),
.Y(n_4783)
);

BUFx2_ASAP7_75t_L g4784 ( 
.A(n_4680),
.Y(n_4784)
);

AND2x4_ASAP7_75t_L g4785 ( 
.A(n_4697),
.B(n_4445),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4604),
.B(n_4470),
.Y(n_4786)
);

INVx2_ASAP7_75t_L g4787 ( 
.A(n_4634),
.Y(n_4787)
);

INVx2_ASAP7_75t_L g4788 ( 
.A(n_4634),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4602),
.B(n_4477),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4593),
.Y(n_4790)
);

INVx2_ASAP7_75t_L g4791 ( 
.A(n_4680),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4606),
.Y(n_4792)
);

AOI222xp33_ASAP7_75t_L g4793 ( 
.A1(n_4583),
.A2(n_4481),
.B1(n_4470),
.B2(n_4462),
.C1(n_4559),
.C2(n_4436),
.Y(n_4793)
);

INVx2_ASAP7_75t_L g4794 ( 
.A(n_4651),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4587),
.B(n_4481),
.Y(n_4795)
);

INVx2_ASAP7_75t_L g4796 ( 
.A(n_4684),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4581),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4576),
.B(n_4548),
.Y(n_4798)
);

INVx2_ASAP7_75t_SL g4799 ( 
.A(n_4647),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4660),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_4662),
.Y(n_4801)
);

AOI22xp33_ASAP7_75t_L g4802 ( 
.A1(n_4598),
.A2(n_4515),
.B1(n_4542),
.B2(n_4570),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4667),
.Y(n_4803)
);

OR2x2_ASAP7_75t_L g4804 ( 
.A(n_4691),
.B(n_4480),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4596),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4613),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4692),
.B(n_4445),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4591),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4607),
.B(n_4548),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4599),
.B(n_4439),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4629),
.Y(n_4811)
);

OAI221xp5_ASAP7_75t_L g4812 ( 
.A1(n_4773),
.A2(n_4629),
.B1(n_4703),
.B2(n_4655),
.C(n_4689),
.Y(n_4812)
);

INVxp67_ASAP7_75t_SL g4813 ( 
.A(n_4771),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4723),
.Y(n_4814)
);

AOI22xp33_ASAP7_75t_L g4815 ( 
.A1(n_4797),
.A2(n_4622),
.B1(n_4675),
.B2(n_4641),
.Y(n_4815)
);

AOI22xp33_ASAP7_75t_SL g4816 ( 
.A1(n_4798),
.A2(n_4636),
.B1(n_4661),
.B2(n_4648),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4711),
.Y(n_4817)
);

OAI33xp33_ASAP7_75t_L g4818 ( 
.A1(n_4805),
.A2(n_4645),
.A3(n_4682),
.B1(n_4664),
.B2(n_4619),
.B3(n_4630),
.Y(n_4818)
);

AND2x4_ASAP7_75t_L g4819 ( 
.A(n_4711),
.B(n_4480),
.Y(n_4819)
);

AO21x2_ASAP7_75t_L g4820 ( 
.A1(n_4707),
.A2(n_4625),
.B(n_4703),
.Y(n_4820)
);

INVxp67_ASAP7_75t_L g4821 ( 
.A(n_4784),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4808),
.A2(n_4801),
.B1(n_4811),
.B2(n_4735),
.Y(n_4822)
);

AOI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4808),
.A2(n_4677),
.B1(n_4638),
.B2(n_4646),
.Y(n_4823)
);

AND2x4_ASAP7_75t_L g4824 ( 
.A(n_4727),
.B(n_4441),
.Y(n_4824)
);

O2A1O1Ixp5_ASAP7_75t_L g4825 ( 
.A1(n_4727),
.A2(n_4654),
.B(n_4653),
.C(n_4617),
.Y(n_4825)
);

NAND3xp33_ASAP7_75t_L g4826 ( 
.A(n_4741),
.B(n_4809),
.C(n_4793),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4713),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_4715),
.A2(n_4623),
.B1(n_4603),
.B2(n_4643),
.Y(n_4828)
);

INVx3_ASAP7_75t_L g4829 ( 
.A(n_4724),
.Y(n_4829)
);

AOI221xp5_ASAP7_75t_L g4830 ( 
.A1(n_4803),
.A2(n_4615),
.B1(n_4614),
.B2(n_4605),
.C(n_4681),
.Y(n_4830)
);

INVx1_ASAP7_75t_SL g4831 ( 
.A(n_4766),
.Y(n_4831)
);

AOI22xp33_ASAP7_75t_SL g4832 ( 
.A1(n_4759),
.A2(n_4542),
.B1(n_4451),
.B2(n_4487),
.Y(n_4832)
);

OAI211xp5_ASAP7_75t_L g4833 ( 
.A1(n_4802),
.A2(n_4690),
.B(n_4673),
.C(n_4674),
.Y(n_4833)
);

AOI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4735),
.A2(n_4451),
.B(n_4656),
.Y(n_4834)
);

HB1xp67_ASAP7_75t_L g4835 ( 
.A(n_4746),
.Y(n_4835)
);

AOI22xp33_ASAP7_75t_L g4836 ( 
.A1(n_4801),
.A2(n_4571),
.B1(n_4570),
.B2(n_4487),
.Y(n_4836)
);

OR2x2_ASAP7_75t_L g4837 ( 
.A(n_4789),
.B(n_4548),
.Y(n_4837)
);

INVx2_ASAP7_75t_SL g4838 ( 
.A(n_4724),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4746),
.B(n_4548),
.Y(n_4839)
);

AND2x2_ASAP7_75t_L g4840 ( 
.A(n_4766),
.B(n_4657),
.Y(n_4840)
);

AOI22xp33_ASAP7_75t_L g4841 ( 
.A1(n_4792),
.A2(n_4571),
.B1(n_4487),
.B2(n_4696),
.Y(n_4841)
);

NOR2xp33_ASAP7_75t_L g4842 ( 
.A(n_4752),
.B(n_4758),
.Y(n_4842)
);

NAND3xp33_ASAP7_75t_SL g4843 ( 
.A(n_4774),
.B(n_4644),
.C(n_4702),
.Y(n_4843)
);

OAI21xp5_ASAP7_75t_SL g4844 ( 
.A1(n_4800),
.A2(n_4701),
.B(n_4441),
.Y(n_4844)
);

NOR3xp33_ASAP7_75t_L g4845 ( 
.A(n_4727),
.B(n_4489),
.C(n_4483),
.Y(n_4845)
);

OAI222xp33_ASAP7_75t_L g4846 ( 
.A1(n_4790),
.A2(n_4489),
.B1(n_4469),
.B2(n_4471),
.C1(n_4483),
.C2(n_4465),
.Y(n_4846)
);

INVxp67_ASAP7_75t_SL g4847 ( 
.A(n_4724),
.Y(n_4847)
);

AOI22xp33_ASAP7_75t_L g4848 ( 
.A1(n_4806),
.A2(n_4471),
.B1(n_4469),
.B2(n_4467),
.Y(n_4848)
);

OAI22xp5_ASAP7_75t_L g4849 ( 
.A1(n_4715),
.A2(n_4762),
.B1(n_4784),
.B2(n_4724),
.Y(n_4849)
);

AOI211xp5_ASAP7_75t_L g4850 ( 
.A1(n_4733),
.A2(n_4467),
.B(n_4465),
.C(n_305),
.Y(n_4850)
);

AND2x2_ASAP7_75t_L g4851 ( 
.A(n_4751),
.B(n_4471),
.Y(n_4851)
);

OAI22xp33_ASAP7_75t_L g4852 ( 
.A1(n_4762),
.A2(n_306),
.B1(n_303),
.B2(n_304),
.Y(n_4852)
);

OAI33xp33_ASAP7_75t_L g4853 ( 
.A1(n_4781),
.A2(n_303),
.A3(n_307),
.B1(n_308),
.B2(n_309),
.B3(n_310),
.Y(n_4853)
);

OAI22xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4768),
.A2(n_311),
.B1(n_307),
.B2(n_308),
.Y(n_4854)
);

OAI221xp5_ASAP7_75t_L g4855 ( 
.A1(n_4768),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.C(n_315),
.Y(n_4855)
);

OAI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4791),
.A2(n_316),
.B1(n_312),
.B2(n_315),
.Y(n_4856)
);

OAI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4791),
.A2(n_322),
.B1(n_316),
.B2(n_318),
.Y(n_4857)
);

HB1xp67_ASAP7_75t_L g4858 ( 
.A(n_4729),
.Y(n_4858)
);

BUFx6f_ASAP7_75t_L g4859 ( 
.A(n_4752),
.Y(n_4859)
);

OR2x2_ASAP7_75t_L g4860 ( 
.A(n_4770),
.B(n_318),
.Y(n_4860)
);

INVx2_ASAP7_75t_L g4861 ( 
.A(n_4717),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4717),
.Y(n_4862)
);

OAI221xp5_ASAP7_75t_L g4863 ( 
.A1(n_4777),
.A2(n_4799),
.B1(n_4770),
.B2(n_4764),
.C(n_4717),
.Y(n_4863)
);

OAI22xp5_ASAP7_75t_L g4864 ( 
.A1(n_4729),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_4864)
);

OAI211xp5_ASAP7_75t_L g4865 ( 
.A1(n_4804),
.A2(n_323),
.B(n_326),
.C(n_328),
.Y(n_4865)
);

INVxp67_ASAP7_75t_SL g4866 ( 
.A(n_4737),
.Y(n_4866)
);

OR2x2_ASAP7_75t_L g4867 ( 
.A(n_4776),
.B(n_328),
.Y(n_4867)
);

AO21x2_ASAP7_75t_L g4868 ( 
.A1(n_4780),
.A2(n_4788),
.B(n_4787),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4751),
.B(n_330),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4776),
.Y(n_4870)
);

OA222x2_ASAP7_75t_L g4871 ( 
.A1(n_4786),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.C1(n_336),
.C2(n_337),
.Y(n_4871)
);

NAND4xp25_ASAP7_75t_L g4872 ( 
.A(n_4810),
.B(n_331),
.C(n_336),
.D(n_338),
.Y(n_4872)
);

AOI221xp5_ASAP7_75t_L g4873 ( 
.A1(n_4810),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.C(n_342),
.Y(n_4873)
);

NOR2x1p5_ASAP7_75t_L g4874 ( 
.A(n_4782),
.B(n_339),
.Y(n_4874)
);

AOI22xp33_ASAP7_75t_L g4875 ( 
.A1(n_4745),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4795),
.B(n_4783),
.Y(n_4876)
);

AOI221xp5_ASAP7_75t_SL g4877 ( 
.A1(n_4765),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.C(n_347),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4769),
.B(n_345),
.Y(n_4878)
);

INVx2_ASAP7_75t_L g4879 ( 
.A(n_4737),
.Y(n_4879)
);

OA21x2_ASAP7_75t_L g4880 ( 
.A1(n_4780),
.A2(n_346),
.B(n_347),
.Y(n_4880)
);

OAI22xp5_ASAP7_75t_L g4881 ( 
.A1(n_4777),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_4881)
);

INVx3_ASAP7_75t_L g4882 ( 
.A(n_4737),
.Y(n_4882)
);

HB1xp67_ASAP7_75t_L g4883 ( 
.A(n_4835),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4829),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4858),
.Y(n_4885)
);

HB1xp67_ASAP7_75t_L g4886 ( 
.A(n_4821),
.Y(n_4886)
);

BUFx2_ASAP7_75t_SL g4887 ( 
.A(n_4859),
.Y(n_4887)
);

HB1xp67_ASAP7_75t_L g4888 ( 
.A(n_4868),
.Y(n_4888)
);

NOR2xp33_ASAP7_75t_L g4889 ( 
.A(n_4859),
.B(n_4799),
.Y(n_4889)
);

AND2x2_ASAP7_75t_L g4890 ( 
.A(n_4831),
.B(n_4769),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4868),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4814),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4822),
.B(n_4795),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4827),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4867),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4870),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4880),
.Y(n_4897)
);

OR2x2_ASAP7_75t_L g4898 ( 
.A(n_4876),
.B(n_4761),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4829),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_L g4900 ( 
.A(n_4816),
.B(n_4760),
.Y(n_4900)
);

INVx2_ASAP7_75t_L g4901 ( 
.A(n_4882),
.Y(n_4901)
);

INVx1_ASAP7_75t_L g4902 ( 
.A(n_4880),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4847),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4840),
.B(n_4716),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_4817),
.B(n_4716),
.Y(n_4905)
);

NOR2xp33_ASAP7_75t_L g4906 ( 
.A(n_4859),
.B(n_4760),
.Y(n_4906)
);

AND2x2_ASAP7_75t_L g4907 ( 
.A(n_4838),
.B(n_4764),
.Y(n_4907)
);

NAND2x1p5_ASAP7_75t_L g4908 ( 
.A(n_4882),
.B(n_4737),
.Y(n_4908)
);

OR2x2_ASAP7_75t_L g4909 ( 
.A(n_4820),
.B(n_4709),
.Y(n_4909)
);

AND2x2_ASAP7_75t_L g4910 ( 
.A(n_4866),
.B(n_4764),
.Y(n_4910)
);

INVx2_ASAP7_75t_L g4911 ( 
.A(n_4861),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4860),
.Y(n_4912)
);

AND2x4_ASAP7_75t_L g4913 ( 
.A(n_4862),
.B(n_4719),
.Y(n_4913)
);

AND2x2_ASAP7_75t_L g4914 ( 
.A(n_4842),
.B(n_4748),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4813),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4879),
.Y(n_4916)
);

OR2x2_ASAP7_75t_L g4917 ( 
.A(n_4820),
.B(n_4706),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4878),
.Y(n_4918)
);

NAND4xp25_ASAP7_75t_L g4919 ( 
.A(n_4826),
.B(n_4755),
.C(n_4745),
.D(n_4804),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4839),
.Y(n_4920)
);

INVxp67_ASAP7_75t_L g4921 ( 
.A(n_4869),
.Y(n_4921)
);

OR2x2_ASAP7_75t_L g4922 ( 
.A(n_4837),
.B(n_4734),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4819),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4819),
.Y(n_4924)
);

AND2x4_ASAP7_75t_SL g4925 ( 
.A(n_4823),
.B(n_4748),
.Y(n_4925)
);

HB1xp67_ASAP7_75t_L g4926 ( 
.A(n_4874),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4863),
.Y(n_4927)
);

OR2x2_ASAP7_75t_L g4928 ( 
.A(n_4844),
.B(n_4718),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4914),
.B(n_4849),
.Y(n_4929)
);

AND2x4_ASAP7_75t_L g4930 ( 
.A(n_4910),
.B(n_4824),
.Y(n_4930)
);

HB1xp67_ASAP7_75t_L g4931 ( 
.A(n_4883),
.Y(n_4931)
);

INVx1_ASAP7_75t_L g4932 ( 
.A(n_4883),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4886),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4908),
.Y(n_4934)
);

NAND4xp25_ASAP7_75t_L g4935 ( 
.A(n_4919),
.B(n_4815),
.C(n_4812),
.D(n_4825),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4886),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4926),
.B(n_4830),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4888),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4888),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_4908),
.Y(n_4940)
);

OAI221xp5_ASAP7_75t_L g4941 ( 
.A1(n_4909),
.A2(n_4850),
.B1(n_4832),
.B2(n_4873),
.C(n_4865),
.Y(n_4941)
);

INVx3_ASAP7_75t_L g4942 ( 
.A(n_4913),
.Y(n_4942)
);

AO21x2_ASAP7_75t_L g4943 ( 
.A1(n_4891),
.A2(n_4871),
.B(n_4852),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4885),
.Y(n_4944)
);

AND2x4_ASAP7_75t_L g4945 ( 
.A(n_4910),
.B(n_4824),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4915),
.Y(n_4946)
);

NAND5xp2_ASAP7_75t_L g4947 ( 
.A(n_4927),
.B(n_4877),
.C(n_4875),
.D(n_4855),
.E(n_4834),
.Y(n_4947)
);

AND2x2_ASAP7_75t_L g4948 ( 
.A(n_4926),
.B(n_4890),
.Y(n_4948)
);

INVx2_ASAP7_75t_L g4949 ( 
.A(n_4917),
.Y(n_4949)
);

NAND4xp25_ASAP7_75t_L g4950 ( 
.A(n_4900),
.B(n_4872),
.C(n_4828),
.D(n_4841),
.Y(n_4950)
);

AOI322xp5_ASAP7_75t_L g4951 ( 
.A1(n_4893),
.A2(n_4843),
.A3(n_4871),
.B1(n_4836),
.B2(n_4848),
.C1(n_4788),
.C2(n_4787),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4925),
.B(n_4854),
.Y(n_4952)
);

INVx2_ASAP7_75t_L g4953 ( 
.A(n_4913),
.Y(n_4953)
);

AOI22xp33_ASAP7_75t_L g4954 ( 
.A1(n_4925),
.A2(n_4818),
.B1(n_4845),
.B2(n_4763),
.Y(n_4954)
);

AND2x2_ASAP7_75t_L g4955 ( 
.A(n_4907),
.B(n_4719),
.Y(n_4955)
);

AOI22xp33_ASAP7_75t_L g4956 ( 
.A1(n_4889),
.A2(n_4928),
.B1(n_4904),
.B2(n_4918),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4912),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4903),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4897),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_4948),
.B(n_4921),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4931),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4932),
.Y(n_4962)
);

AND2x2_ASAP7_75t_L g4963 ( 
.A(n_4948),
.B(n_4887),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4955),
.B(n_4889),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4959),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4959),
.Y(n_4966)
);

OAI21xp33_ASAP7_75t_SL g4967 ( 
.A1(n_4951),
.A2(n_4902),
.B(n_4906),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4933),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4936),
.Y(n_4969)
);

INVx2_ASAP7_75t_SL g4970 ( 
.A(n_4942),
.Y(n_4970)
);

HB1xp67_ASAP7_75t_L g4971 ( 
.A(n_4943),
.Y(n_4971)
);

AND2x6_ASAP7_75t_SL g4972 ( 
.A(n_4937),
.B(n_4906),
.Y(n_4972)
);

INVxp67_ASAP7_75t_L g4973 ( 
.A(n_4942),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4929),
.B(n_4921),
.Y(n_4974)
);

OR2x2_ASAP7_75t_L g4975 ( 
.A(n_4952),
.B(n_4898),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4942),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4930),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4929),
.B(n_4956),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4930),
.B(n_4884),
.Y(n_4979)
);

OAI31xp33_ASAP7_75t_L g4980 ( 
.A1(n_4971),
.A2(n_4941),
.A3(n_4935),
.B(n_4947),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4970),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4971),
.B(n_4943),
.Y(n_4982)
);

OR2x2_ASAP7_75t_L g4983 ( 
.A(n_4974),
.B(n_4943),
.Y(n_4983)
);

OR2x2_ASAP7_75t_L g4984 ( 
.A(n_4960),
.B(n_4895),
.Y(n_4984)
);

NAND3xp33_ASAP7_75t_L g4985 ( 
.A(n_4967),
.B(n_4949),
.C(n_4954),
.Y(n_4985)
);

AND2x2_ASAP7_75t_L g4986 ( 
.A(n_4963),
.B(n_4905),
.Y(n_4986)
);

INVx2_ASAP7_75t_L g4987 ( 
.A(n_4970),
.Y(n_4987)
);

AND2x2_ASAP7_75t_L g4988 ( 
.A(n_4964),
.B(n_4930),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4977),
.B(n_4945),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4973),
.B(n_4949),
.Y(n_4990)
);

OR2x2_ASAP7_75t_L g4991 ( 
.A(n_4975),
.B(n_4958),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4976),
.Y(n_4992)
);

AOI211xp5_ASAP7_75t_SL g4993 ( 
.A1(n_4973),
.A2(n_4938),
.B(n_4939),
.C(n_4864),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4977),
.B(n_4945),
.Y(n_4994)
);

AND2x2_ASAP7_75t_SL g4995 ( 
.A(n_4978),
.B(n_4945),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4961),
.B(n_4953),
.Y(n_4996)
);

AOI22xp33_ASAP7_75t_L g4997 ( 
.A1(n_4968),
.A2(n_4950),
.B1(n_4955),
.B2(n_4944),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4976),
.B(n_4953),
.Y(n_4998)
);

INVx2_ASAP7_75t_L g4999 ( 
.A(n_4979),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4998),
.Y(n_5000)
);

OR2x2_ASAP7_75t_L g5001 ( 
.A(n_4983),
.B(n_4946),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_L g5002 ( 
.A(n_4995),
.B(n_4969),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4994),
.B(n_4962),
.Y(n_5003)
);

NOR2xp33_ASAP7_75t_SL g5004 ( 
.A(n_4988),
.B(n_4934),
.Y(n_5004)
);

OR2x2_ASAP7_75t_L g5005 ( 
.A(n_4989),
.B(n_4957),
.Y(n_5005)
);

AND2x4_ASAP7_75t_L g5006 ( 
.A(n_4981),
.B(n_4965),
.Y(n_5006)
);

OR2x2_ASAP7_75t_L g5007 ( 
.A(n_4996),
.B(n_4916),
.Y(n_5007)
);

INVx3_ASAP7_75t_SL g5008 ( 
.A(n_4987),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4990),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4991),
.B(n_4984),
.Y(n_5010)
);

AND2x2_ASAP7_75t_L g5011 ( 
.A(n_4986),
.B(n_4884),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4999),
.B(n_4899),
.Y(n_5012)
);

HB1xp67_ASAP7_75t_L g5013 ( 
.A(n_4982),
.Y(n_5013)
);

AND2x2_ASAP7_75t_L g5014 ( 
.A(n_5011),
.B(n_4997),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_5008),
.B(n_4993),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_5000),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_5004),
.B(n_4993),
.Y(n_5017)
);

XOR2xp5_ASAP7_75t_L g5018 ( 
.A(n_5010),
.B(n_4985),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_5012),
.B(n_4980),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_5006),
.B(n_4980),
.Y(n_5020)
);

HB1xp67_ASAP7_75t_L g5021 ( 
.A(n_5006),
.Y(n_5021)
);

OR2x2_ASAP7_75t_L g5022 ( 
.A(n_5003),
.B(n_4990),
.Y(n_5022)
);

HB1xp67_ASAP7_75t_L g5023 ( 
.A(n_5002),
.Y(n_5023)
);

AND2x2_ASAP7_75t_L g5024 ( 
.A(n_5009),
.B(n_4992),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_5021),
.Y(n_5025)
);

INVx1_ASAP7_75t_SL g5026 ( 
.A(n_5015),
.Y(n_5026)
);

OAI332xp33_ASAP7_75t_L g5027 ( 
.A1(n_5020),
.A2(n_4982),
.A3(n_5005),
.B1(n_5001),
.B2(n_4985),
.B3(n_4966),
.C1(n_4972),
.C2(n_5007),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_5023),
.Y(n_5028)
);

AOI22xp5_ASAP7_75t_L g5029 ( 
.A1(n_5018),
.A2(n_4899),
.B1(n_4940),
.B2(n_4934),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_5014),
.B(n_5013),
.Y(n_5030)
);

INVxp67_ASAP7_75t_L g5031 ( 
.A(n_5017),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_5019),
.A2(n_5016),
.B(n_5022),
.Y(n_5032)
);

OAI22xp5_ASAP7_75t_L g5033 ( 
.A1(n_5024),
.A2(n_4940),
.B1(n_4901),
.B2(n_4911),
.Y(n_5033)
);

OR2x2_ASAP7_75t_L g5034 ( 
.A(n_5021),
.B(n_4896),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_5021),
.Y(n_5035)
);

AND2x2_ASAP7_75t_L g5036 ( 
.A(n_5014),
.B(n_4901),
.Y(n_5036)
);

OAI22xp33_ASAP7_75t_L g5037 ( 
.A1(n_5017),
.A2(n_4922),
.B1(n_4911),
.B2(n_4923),
.Y(n_5037)
);

AND2x2_ASAP7_75t_L g5038 ( 
.A(n_5036),
.B(n_4913),
.Y(n_5038)
);

NOR2x1_ASAP7_75t_L g5039 ( 
.A(n_5035),
.B(n_4938),
.Y(n_5039)
);

NAND2x1p5_ASAP7_75t_L g5040 ( 
.A(n_5028),
.B(n_5025),
.Y(n_5040)
);

OR2x2_ASAP7_75t_L g5041 ( 
.A(n_5034),
.B(n_4892),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_5029),
.B(n_4894),
.Y(n_5042)
);

OAI32xp33_ASAP7_75t_L g5043 ( 
.A1(n_5030),
.A2(n_4939),
.A3(n_4924),
.B1(n_4920),
.B2(n_4881),
.Y(n_5043)
);

NAND2x1_ASAP7_75t_L g5044 ( 
.A(n_5033),
.B(n_4721),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_5037),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_5027),
.B(n_4755),
.Y(n_5046)
);

O2A1O1Ixp33_ASAP7_75t_L g5047 ( 
.A1(n_5032),
.A2(n_4857),
.B(n_4856),
.C(n_4853),
.Y(n_5047)
);

AND2x2_ASAP7_75t_L g5048 ( 
.A(n_5038),
.B(n_5026),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_5039),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_5044),
.B(n_5031),
.Y(n_5050)
);

AOI31xp33_ASAP7_75t_L g5051 ( 
.A1(n_5040),
.A2(n_4778),
.A3(n_4767),
.B(n_4833),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_5041),
.Y(n_5052)
);

OAI22xp33_ASAP7_75t_SL g5053 ( 
.A1(n_5046),
.A2(n_5045),
.B1(n_5042),
.B2(n_5043),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_5047),
.Y(n_5054)
);

AND2x2_ASAP7_75t_L g5055 ( 
.A(n_5038),
.B(n_4721),
.Y(n_5055)
);

INVxp67_ASAP7_75t_SL g5056 ( 
.A(n_5039),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_5055),
.B(n_5048),
.Y(n_5057)
);

INVxp67_ASAP7_75t_L g5058 ( 
.A(n_5056),
.Y(n_5058)
);

AOI22xp5_ASAP7_75t_SL g5059 ( 
.A1(n_5049),
.A2(n_4785),
.B1(n_4725),
.B2(n_4743),
.Y(n_5059)
);

OA21x2_ASAP7_75t_L g5060 ( 
.A1(n_5050),
.A2(n_4851),
.B(n_4738),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_5052),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5051),
.B(n_4763),
.Y(n_5062)
);

AOI221xp5_ASAP7_75t_L g5063 ( 
.A1(n_5051),
.A2(n_4846),
.B1(n_4763),
.B2(n_4785),
.C(n_4708),
.Y(n_5063)
);

OAI211xp5_ASAP7_75t_SL g5064 ( 
.A1(n_5054),
.A2(n_5053),
.B(n_4739),
.C(n_4786),
.Y(n_5064)
);

XNOR2xp5_ASAP7_75t_L g5065 ( 
.A(n_5048),
.B(n_348),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_L g5066 ( 
.A(n_5055),
.B(n_4744),
.Y(n_5066)
);

INVxp67_ASAP7_75t_L g5067 ( 
.A(n_5056),
.Y(n_5067)
);

INVx1_ASAP7_75t_L g5068 ( 
.A(n_5056),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_5055),
.B(n_4744),
.Y(n_5069)
);

XNOR2xp5_ASAP7_75t_L g5070 ( 
.A(n_5048),
.B(n_349),
.Y(n_5070)
);

NOR3xp33_ASAP7_75t_L g5071 ( 
.A(n_5057),
.B(n_5061),
.C(n_5064),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_5065),
.B(n_4708),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5070),
.Y(n_5073)
);

XNOR2x1_ASAP7_75t_L g5074 ( 
.A(n_5068),
.B(n_351),
.Y(n_5074)
);

INVxp33_ASAP7_75t_L g5075 ( 
.A(n_5066),
.Y(n_5075)
);

AOI21xp5_ASAP7_75t_L g5076 ( 
.A1(n_5058),
.A2(n_4779),
.B(n_4731),
.Y(n_5076)
);

NAND3xp33_ASAP7_75t_L g5077 ( 
.A(n_5067),
.B(n_4796),
.C(n_4794),
.Y(n_5077)
);

NOR3xp33_ASAP7_75t_L g5078 ( 
.A(n_5069),
.B(n_4785),
.C(n_4794),
.Y(n_5078)
);

AOI211xp5_ASAP7_75t_L g5079 ( 
.A1(n_5062),
.A2(n_4796),
.B(n_4749),
.C(n_4754),
.Y(n_5079)
);

NOR3xp33_ASAP7_75t_L g5080 ( 
.A(n_5063),
.B(n_4726),
.C(n_4720),
.Y(n_5080)
);

NAND4xp75_ASAP7_75t_SL g5081 ( 
.A(n_5060),
.B(n_4807),
.C(n_4772),
.D(n_4732),
.Y(n_5081)
);

NOR2xp33_ASAP7_75t_L g5082 ( 
.A(n_5059),
.B(n_5060),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_5065),
.Y(n_5083)
);

NOR3xp33_ASAP7_75t_L g5084 ( 
.A(n_5057),
.B(n_4726),
.C(n_4720),
.Y(n_5084)
);

OAI211xp5_ASAP7_75t_SL g5085 ( 
.A1(n_5058),
.A2(n_4747),
.B(n_353),
.C(n_354),
.Y(n_5085)
);

NOR2x1_ASAP7_75t_L g5086 ( 
.A(n_5064),
.B(n_4725),
.Y(n_5086)
);

AOI22xp33_ASAP7_75t_L g5087 ( 
.A1(n_5064),
.A2(n_4725),
.B1(n_4742),
.B2(n_4807),
.Y(n_5087)
);

NAND3xp33_ASAP7_75t_L g5088 ( 
.A(n_5064),
.B(n_4730),
.C(n_4714),
.Y(n_5088)
);

OA22x2_ASAP7_75t_L g5089 ( 
.A1(n_5068),
.A2(n_4742),
.B1(n_4730),
.B2(n_4712),
.Y(n_5089)
);

AOI21xp5_ASAP7_75t_L g5090 ( 
.A1(n_5057),
.A2(n_4714),
.B(n_4712),
.Y(n_5090)
);

NAND3xp33_ASAP7_75t_L g5091 ( 
.A(n_5064),
.B(n_4740),
.C(n_4736),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_5057),
.A2(n_4740),
.B(n_4736),
.Y(n_5092)
);

HB1xp67_ASAP7_75t_L g5093 ( 
.A(n_5065),
.Y(n_5093)
);

NOR4xp25_ASAP7_75t_L g5094 ( 
.A(n_5064),
.B(n_4753),
.C(n_4750),
.D(n_4757),
.Y(n_5094)
);

OAI22xp33_ASAP7_75t_L g5095 ( 
.A1(n_5075),
.A2(n_4710),
.B1(n_4775),
.B2(n_4750),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_5082),
.A2(n_4757),
.B(n_4753),
.Y(n_5096)
);

AOI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_5071),
.A2(n_4783),
.B(n_4756),
.Y(n_5097)
);

XNOR2xp5_ASAP7_75t_L g5098 ( 
.A(n_5074),
.B(n_352),
.Y(n_5098)
);

AOI21xp5_ASAP7_75t_L g5099 ( 
.A1(n_5093),
.A2(n_4756),
.B(n_4742),
.Y(n_5099)
);

OAI211xp5_ASAP7_75t_L g5100 ( 
.A1(n_5085),
.A2(n_352),
.B(n_355),
.C(n_356),
.Y(n_5100)
);

AOI32xp33_ASAP7_75t_L g5101 ( 
.A1(n_5086),
.A2(n_4772),
.A3(n_4722),
.B1(n_4732),
.B2(n_4728),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5089),
.Y(n_5102)
);

INVxp67_ASAP7_75t_SL g5103 ( 
.A(n_5073),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5072),
.Y(n_5104)
);

AOI21xp5_ASAP7_75t_L g5105 ( 
.A1(n_5083),
.A2(n_4710),
.B(n_4728),
.Y(n_5105)
);

INVx1_ASAP7_75t_SL g5106 ( 
.A(n_5081),
.Y(n_5106)
);

NOR2xp33_ASAP7_75t_L g5107 ( 
.A(n_5076),
.B(n_4728),
.Y(n_5107)
);

AOI321xp33_ASAP7_75t_L g5108 ( 
.A1(n_5094),
.A2(n_4722),
.A3(n_4775),
.B1(n_358),
.B2(n_360),
.C(n_362),
.Y(n_5108)
);

NAND3xp33_ASAP7_75t_SL g5109 ( 
.A(n_5084),
.B(n_356),
.C(n_357),
.Y(n_5109)
);

AO22x1_ASAP7_75t_L g5110 ( 
.A1(n_5078),
.A2(n_362),
.B1(n_364),
.B2(n_366),
.Y(n_5110)
);

AOI22xp5_ASAP7_75t_L g5111 ( 
.A1(n_5080),
.A2(n_366),
.B1(n_367),
.B2(n_369),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_5088),
.Y(n_5112)
);

OAI31xp33_ASAP7_75t_L g5113 ( 
.A1(n_5077),
.A2(n_367),
.A3(n_370),
.B(n_371),
.Y(n_5113)
);

AOI21xp33_ASAP7_75t_L g5114 ( 
.A1(n_5079),
.A2(n_370),
.B(n_372),
.Y(n_5114)
);

AOI21xp33_ASAP7_75t_SL g5115 ( 
.A1(n_5091),
.A2(n_373),
.B(n_374),
.Y(n_5115)
);

NAND3xp33_ASAP7_75t_L g5116 ( 
.A(n_5090),
.B(n_5092),
.C(n_5087),
.Y(n_5116)
);

NOR2xp33_ASAP7_75t_L g5117 ( 
.A(n_5075),
.B(n_373),
.Y(n_5117)
);

OAI21xp33_ASAP7_75t_L g5118 ( 
.A1(n_5075),
.A2(n_375),
.B(n_376),
.Y(n_5118)
);

HB1xp67_ASAP7_75t_L g5119 ( 
.A(n_5082),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_5086),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_5086),
.B(n_376),
.Y(n_5121)
);

AND3x1_ASAP7_75t_L g5122 ( 
.A(n_5113),
.B(n_377),
.C(n_378),
.Y(n_5122)
);

NOR3xp33_ASAP7_75t_SL g5123 ( 
.A(n_5109),
.B(n_377),
.C(n_379),
.Y(n_5123)
);

NOR2xp33_ASAP7_75t_L g5124 ( 
.A(n_5118),
.B(n_379),
.Y(n_5124)
);

AND5x1_ASAP7_75t_L g5125 ( 
.A(n_5108),
.B(n_380),
.C(n_383),
.D(n_386),
.E(n_387),
.Y(n_5125)
);

NOR3xp33_ASAP7_75t_L g5126 ( 
.A(n_5119),
.B(n_380),
.C(n_383),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_5099),
.B(n_387),
.Y(n_5127)
);

NOR2x1_ASAP7_75t_L g5128 ( 
.A(n_5120),
.B(n_389),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_5121),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_L g5130 ( 
.A(n_5110),
.B(n_389),
.Y(n_5130)
);

NOR3xp33_ASAP7_75t_SL g5131 ( 
.A(n_5116),
.B(n_390),
.C(n_391),
.Y(n_5131)
);

NOR3xp33_ASAP7_75t_L g5132 ( 
.A(n_5103),
.B(n_390),
.C(n_392),
.Y(n_5132)
);

NOR2xp33_ASAP7_75t_L g5133 ( 
.A(n_5100),
.B(n_392),
.Y(n_5133)
);

NOR3xp33_ASAP7_75t_L g5134 ( 
.A(n_5117),
.B(n_393),
.C(n_394),
.Y(n_5134)
);

OAI322xp33_ASAP7_75t_L g5135 ( 
.A1(n_5106),
.A2(n_393),
.A3(n_394),
.B1(n_396),
.B2(n_397),
.C1(n_398),
.C2(n_401),
.Y(n_5135)
);

NOR2x1_ASAP7_75t_L g5136 ( 
.A(n_5098),
.B(n_397),
.Y(n_5136)
);

NAND3xp33_ASAP7_75t_L g5137 ( 
.A(n_5111),
.B(n_401),
.C(n_402),
.Y(n_5137)
);

NOR3xp33_ASAP7_75t_L g5138 ( 
.A(n_5104),
.B(n_402),
.C(n_412),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_5097),
.B(n_413),
.Y(n_5139)
);

NOR2x1_ASAP7_75t_L g5140 ( 
.A(n_5102),
.B(n_414),
.Y(n_5140)
);

O2A1O1Ixp33_ASAP7_75t_L g5141 ( 
.A1(n_5114),
.A2(n_416),
.B(n_417),
.C(n_420),
.Y(n_5141)
);

NOR4xp75_ASAP7_75t_L g5142 ( 
.A(n_5115),
.B(n_5112),
.C(n_5107),
.D(n_5096),
.Y(n_5142)
);

NAND4xp75_ASAP7_75t_L g5143 ( 
.A(n_5105),
.B(n_421),
.C(n_428),
.D(n_435),
.Y(n_5143)
);

AOI211xp5_ASAP7_75t_SL g5144 ( 
.A1(n_5095),
.A2(n_438),
.B(n_439),
.C(n_443),
.Y(n_5144)
);

NAND3xp33_ASAP7_75t_L g5145 ( 
.A(n_5101),
.B(n_2239),
.C(n_2236),
.Y(n_5145)
);

O2A1O1Ixp33_ASAP7_75t_SL g5146 ( 
.A1(n_5130),
.A2(n_444),
.B(n_446),
.C(n_449),
.Y(n_5146)
);

AOI221xp5_ASAP7_75t_L g5147 ( 
.A1(n_5122),
.A2(n_2239),
.B1(n_2236),
.B2(n_2226),
.C(n_2222),
.Y(n_5147)
);

NOR2x1p5_ASAP7_75t_L g5148 ( 
.A(n_5127),
.B(n_454),
.Y(n_5148)
);

NOR3xp33_ASAP7_75t_L g5149 ( 
.A(n_5136),
.B(n_456),
.C(n_460),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_5128),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5133),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_5132),
.B(n_463),
.Y(n_5152)
);

INVx2_ASAP7_75t_L g5153 ( 
.A(n_5143),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5140),
.Y(n_5154)
);

AOI211xp5_ASAP7_75t_L g5155 ( 
.A1(n_5137),
.A2(n_468),
.B(n_469),
.C(n_474),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_5126),
.B(n_475),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_5131),
.Y(n_5157)
);

OAI211xp5_ASAP7_75t_SL g5158 ( 
.A1(n_5123),
.A2(n_477),
.B(n_478),
.C(n_479),
.Y(n_5158)
);

OAI221xp5_ASAP7_75t_L g5159 ( 
.A1(n_5125),
.A2(n_482),
.B1(n_484),
.B2(n_485),
.C(n_487),
.Y(n_5159)
);

OAI221xp5_ASAP7_75t_L g5160 ( 
.A1(n_5124),
.A2(n_489),
.B1(n_491),
.B2(n_495),
.C(n_497),
.Y(n_5160)
);

OAI22xp5_ASAP7_75t_L g5161 ( 
.A1(n_5139),
.A2(n_2158),
.B1(n_2181),
.B2(n_2239),
.Y(n_5161)
);

O2A1O1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_5141),
.A2(n_498),
.B(n_501),
.C(n_508),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_5134),
.Y(n_5163)
);

NOR2xp33_ASAP7_75t_L g5164 ( 
.A(n_5159),
.B(n_5129),
.Y(n_5164)
);

OR2x2_ASAP7_75t_L g5165 ( 
.A(n_5150),
.B(n_5138),
.Y(n_5165)
);

NOR2xp67_ASAP7_75t_L g5166 ( 
.A(n_5154),
.B(n_5157),
.Y(n_5166)
);

INVxp67_ASAP7_75t_L g5167 ( 
.A(n_5152),
.Y(n_5167)
);

NAND3xp33_ASAP7_75t_L g5168 ( 
.A(n_5149),
.B(n_5144),
.C(n_5145),
.Y(n_5168)
);

NAND2xp5_ASAP7_75t_SL g5169 ( 
.A(n_5155),
.B(n_5142),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_5148),
.B(n_5135),
.Y(n_5170)
);

NAND5xp2_ASAP7_75t_L g5171 ( 
.A(n_5151),
.B(n_512),
.C(n_513),
.D(n_514),
.E(n_515),
.Y(n_5171)
);

NAND2xp5_ASAP7_75t_L g5172 ( 
.A(n_5146),
.B(n_518),
.Y(n_5172)
);

AND3x4_ASAP7_75t_L g5173 ( 
.A(n_5153),
.B(n_521),
.C(n_523),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_5156),
.Y(n_5174)
);

OAI322xp33_ASAP7_75t_L g5175 ( 
.A1(n_5163),
.A2(n_528),
.A3(n_529),
.B1(n_530),
.B2(n_531),
.C1(n_532),
.C2(n_534),
.Y(n_5175)
);

OR2x2_ASAP7_75t_L g5176 ( 
.A(n_5160),
.B(n_535),
.Y(n_5176)
);

NAND3xp33_ASAP7_75t_SL g5177 ( 
.A(n_5147),
.B(n_537),
.C(n_538),
.Y(n_5177)
);

CKINVDCx6p67_ASAP7_75t_R g5178 ( 
.A(n_5158),
.Y(n_5178)
);

NAND3x1_ASAP7_75t_L g5179 ( 
.A(n_5161),
.B(n_543),
.C(n_545),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_5166),
.B(n_5172),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5178),
.B(n_5162),
.Y(n_5181)
);

AOI22xp5_ASAP7_75t_L g5182 ( 
.A1(n_5164),
.A2(n_2239),
.B1(n_2236),
.B2(n_2226),
.Y(n_5182)
);

NOR5xp2_ASAP7_75t_SL g5183 ( 
.A(n_5169),
.B(n_546),
.C(n_548),
.D(n_550),
.E(n_552),
.Y(n_5183)
);

OAI211xp5_ASAP7_75t_SL g5184 ( 
.A1(n_5165),
.A2(n_554),
.B(n_557),
.C(n_559),
.Y(n_5184)
);

OR2x2_ASAP7_75t_L g5185 ( 
.A(n_5170),
.B(n_560),
.Y(n_5185)
);

NOR3x1_ASAP7_75t_SL g5186 ( 
.A(n_5175),
.B(n_561),
.C(n_562),
.Y(n_5186)
);

OAI221xp5_ASAP7_75t_L g5187 ( 
.A1(n_5168),
.A2(n_564),
.B1(n_570),
.B2(n_572),
.C(n_574),
.Y(n_5187)
);

AND2x2_ASAP7_75t_L g5188 ( 
.A(n_5174),
.B(n_577),
.Y(n_5188)
);

NAND3xp33_ASAP7_75t_L g5189 ( 
.A(n_5167),
.B(n_2236),
.C(n_2226),
.Y(n_5189)
);

OAI22xp5_ASAP7_75t_L g5190 ( 
.A1(n_5173),
.A2(n_2226),
.B1(n_2222),
.B2(n_2218),
.Y(n_5190)
);

NAND5xp2_ASAP7_75t_L g5191 ( 
.A(n_5177),
.B(n_580),
.C(n_581),
.D(n_585),
.E(n_592),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5179),
.B(n_593),
.Y(n_5192)
);

OA22x2_ASAP7_75t_L g5193 ( 
.A1(n_5171),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_5193)
);

NAND3xp33_ASAP7_75t_L g5194 ( 
.A(n_5176),
.B(n_1988),
.C(n_2218),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5166),
.B(n_597),
.Y(n_5195)
);

AOI22xp5_ASAP7_75t_L g5196 ( 
.A1(n_5166),
.A2(n_1988),
.B1(n_2218),
.B2(n_2211),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_5166),
.B(n_599),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_5188),
.Y(n_5198)
);

OR2x2_ASAP7_75t_L g5199 ( 
.A(n_5192),
.B(n_600),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_5186),
.Y(n_5200)
);

AND2x2_ASAP7_75t_L g5201 ( 
.A(n_5193),
.B(n_601),
.Y(n_5201)
);

INVx2_ASAP7_75t_L g5202 ( 
.A(n_5185),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5195),
.Y(n_5203)
);

OAI22xp5_ASAP7_75t_L g5204 ( 
.A1(n_5197),
.A2(n_602),
.B1(n_607),
.B2(n_612),
.Y(n_5204)
);

OAI221xp5_ASAP7_75t_L g5205 ( 
.A1(n_5180),
.A2(n_614),
.B1(n_616),
.B2(n_619),
.C(n_620),
.Y(n_5205)
);

INVx1_ASAP7_75t_SL g5206 ( 
.A(n_5181),
.Y(n_5206)
);

XOR2x1_ASAP7_75t_L g5207 ( 
.A(n_5190),
.B(n_621),
.Y(n_5207)
);

AOI221xp5_ASAP7_75t_L g5208 ( 
.A1(n_5194),
.A2(n_5191),
.B1(n_5189),
.B2(n_5184),
.C(n_5182),
.Y(n_5208)
);

XNOR2xp5_ASAP7_75t_L g5209 ( 
.A(n_5187),
.B(n_622),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_5196),
.A2(n_2222),
.B(n_2218),
.Y(n_5210)
);

NAND3xp33_ASAP7_75t_SL g5211 ( 
.A(n_5206),
.B(n_5183),
.C(n_629),
.Y(n_5211)
);

OAI222xp33_ASAP7_75t_L g5212 ( 
.A1(n_5200),
.A2(n_1528),
.B1(n_1581),
.B2(n_1605),
.C1(n_1637),
.C2(n_1646),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_5201),
.B(n_2222),
.Y(n_5213)
);

AOI21xp5_ASAP7_75t_L g5214 ( 
.A1(n_5209),
.A2(n_2211),
.B(n_2177),
.Y(n_5214)
);

NAND2xp5_ASAP7_75t_L g5215 ( 
.A(n_5207),
.B(n_5198),
.Y(n_5215)
);

OAI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_5199),
.A2(n_2211),
.B1(n_2177),
.B2(n_2169),
.Y(n_5216)
);

NOR3xp33_ASAP7_75t_L g5217 ( 
.A(n_5203),
.B(n_2211),
.C(n_2177),
.Y(n_5217)
);

AOI22x1_ASAP7_75t_L g5218 ( 
.A1(n_5214),
.A2(n_5202),
.B1(n_5210),
.B2(n_5215),
.Y(n_5218)
);

INVx1_ASAP7_75t_SL g5219 ( 
.A(n_5213),
.Y(n_5219)
);

BUFx2_ASAP7_75t_L g5220 ( 
.A(n_5216),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_5211),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_5217),
.B(n_5208),
.Y(n_5222)
);

HB1xp67_ASAP7_75t_L g5223 ( 
.A(n_5212),
.Y(n_5223)
);

OAI22xp5_ASAP7_75t_SL g5224 ( 
.A1(n_5215),
.A2(n_5205),
.B1(n_5204),
.B2(n_2177),
.Y(n_5224)
);

AOI22xp5_ASAP7_75t_L g5225 ( 
.A1(n_5221),
.A2(n_2169),
.B1(n_2166),
.B2(n_2163),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_5218),
.Y(n_5226)
);

NOR2xp67_ASAP7_75t_L g5227 ( 
.A(n_5223),
.B(n_2169),
.Y(n_5227)
);

XOR2xp5_ASAP7_75t_L g5228 ( 
.A(n_5224),
.B(n_2169),
.Y(n_5228)
);

AOI21xp5_ASAP7_75t_L g5229 ( 
.A1(n_5222),
.A2(n_5219),
.B(n_5220),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5224),
.Y(n_5230)
);

CKINVDCx20_ASAP7_75t_R g5231 ( 
.A(n_5229),
.Y(n_5231)
);

OAI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_5226),
.A2(n_2166),
.B1(n_2163),
.B2(n_2160),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_5228),
.Y(n_5233)
);

AOI22x1_ASAP7_75t_L g5234 ( 
.A1(n_5230),
.A2(n_2166),
.B1(n_2163),
.B2(n_2160),
.Y(n_5234)
);

OAI22xp5_ASAP7_75t_L g5235 ( 
.A1(n_5225),
.A2(n_2166),
.B1(n_2163),
.B2(n_2160),
.Y(n_5235)
);

OAI22xp5_ASAP7_75t_L g5236 ( 
.A1(n_5231),
.A2(n_5227),
.B1(n_2160),
.B2(n_2152),
.Y(n_5236)
);

OAI22x1_ASAP7_75t_L g5237 ( 
.A1(n_5233),
.A2(n_1528),
.B1(n_1581),
.B2(n_1605),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5232),
.Y(n_5238)
);

INVx4_ASAP7_75t_L g5239 ( 
.A(n_5234),
.Y(n_5239)
);

OAI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_5238),
.A2(n_5235),
.B(n_1581),
.Y(n_5240)
);

OAI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_5236),
.A2(n_1528),
.B(n_1581),
.Y(n_5241)
);

AOI22xp33_ASAP7_75t_L g5242 ( 
.A1(n_5237),
.A2(n_2152),
.B1(n_2094),
.B2(n_2087),
.Y(n_5242)
);

NOR3xp33_ASAP7_75t_L g5243 ( 
.A(n_5239),
.B(n_2152),
.C(n_2094),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_5241),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5240),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_5243),
.Y(n_5246)
);

INVxp33_ASAP7_75t_SL g5247 ( 
.A(n_5242),
.Y(n_5247)
);

AOI21xp5_ASAP7_75t_L g5248 ( 
.A1(n_5241),
.A2(n_2087),
.B(n_2070),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5241),
.Y(n_5249)
);

INVxp67_ASAP7_75t_SL g5250 ( 
.A(n_5241),
.Y(n_5250)
);

INVx1_ASAP7_75t_L g5251 ( 
.A(n_5241),
.Y(n_5251)
);

AOI22xp33_ASAP7_75t_L g5252 ( 
.A1(n_5247),
.A2(n_1988),
.B1(n_1984),
.B2(n_2070),
.Y(n_5252)
);

AND2x2_ASAP7_75t_L g5253 ( 
.A(n_5250),
.B(n_2070),
.Y(n_5253)
);

AOI22xp5_ASAP7_75t_L g5254 ( 
.A1(n_5245),
.A2(n_2042),
.B1(n_2041),
.B2(n_1988),
.Y(n_5254)
);

INVxp33_ASAP7_75t_SL g5255 ( 
.A(n_5244),
.Y(n_5255)
);

AOI22xp33_ASAP7_75t_L g5256 ( 
.A1(n_5249),
.A2(n_1984),
.B1(n_1965),
.B2(n_2042),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5246),
.Y(n_5257)
);

OAI21xp5_ASAP7_75t_L g5258 ( 
.A1(n_5251),
.A2(n_1528),
.B(n_1581),
.Y(n_5258)
);

AND2x2_ASAP7_75t_L g5259 ( 
.A(n_5248),
.B(n_2041),
.Y(n_5259)
);

INVxp67_ASAP7_75t_L g5260 ( 
.A(n_5253),
.Y(n_5260)
);

BUFx2_ASAP7_75t_L g5261 ( 
.A(n_5257),
.Y(n_5261)
);

AOI22x1_ASAP7_75t_L g5262 ( 
.A1(n_5258),
.A2(n_2041),
.B1(n_1984),
.B2(n_1965),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5259),
.Y(n_5263)
);

OAI31xp33_ASAP7_75t_L g5264 ( 
.A1(n_5255),
.A2(n_1965),
.A3(n_2142),
.B(n_2027),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_5254),
.Y(n_5265)
);

AOI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_5252),
.A2(n_2018),
.B1(n_2115),
.B2(n_2040),
.Y(n_5266)
);

OR2x6_ASAP7_75t_L g5267 ( 
.A(n_5261),
.B(n_5260),
.Y(n_5267)
);

OR2x6_ASAP7_75t_L g5268 ( 
.A(n_5263),
.B(n_5256),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_5265),
.B(n_2142),
.Y(n_5269)
);

AOI21xp5_ASAP7_75t_L g5270 ( 
.A1(n_5267),
.A2(n_5264),
.B(n_5262),
.Y(n_5270)
);

AOI211xp5_ASAP7_75t_L g5271 ( 
.A1(n_5270),
.A2(n_5269),
.B(n_5268),
.C(n_5266),
.Y(n_5271)
);


endmodule