module fake_jpeg_29910_n_273 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_273);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_227;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_69),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_18),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_24),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_89),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_31),
.B1(n_20),
.B2(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_31),
.B1(n_38),
.B2(n_43),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_52),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_63),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_37),
.Y(n_129)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_81),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_106),
.A2(n_120),
.B1(n_121),
.B2(n_128),
.Y(n_133)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_30),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_64),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_66),
.B1(n_67),
.B2(n_59),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_127),
.Y(n_132)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_71),
.A2(n_68),
.B1(n_62),
.B2(n_53),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_84),
.A2(n_49),
.B1(n_48),
.B2(n_41),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_105),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_100),
.A2(n_97),
.B1(n_56),
.B2(n_82),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_115),
.B1(n_105),
.B2(n_97),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_146),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_138),
.B1(n_133),
.B2(n_55),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_146),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_110),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_40),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_40),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_28),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_183),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_143),
.B(n_145),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_149),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_143),
.B1(n_133),
.B2(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_170),
.A2(n_153),
.B1(n_107),
.B2(n_101),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_178),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_146),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_177),
.C(n_136),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_141),
.C(n_131),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_28),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_150),
.B1(n_152),
.B2(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_192),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_173),
.B1(n_183),
.B2(n_166),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_153),
.B1(n_23),
.B2(n_37),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_171),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_140),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_179),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_102),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_200),
.A2(n_177),
.B1(n_180),
.B2(n_171),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_179),
.B1(n_135),
.B2(n_127),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_23),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_175),
.B1(n_174),
.B2(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_208),
.A2(n_200),
.B1(n_186),
.B2(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_182),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_193),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_208),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_187),
.B(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_215),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_204),
.B1(n_212),
.B2(n_114),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_198),
.C(n_191),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_216),
.C(n_227),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_207),
.B1(n_203),
.B2(n_201),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_135),
.B1(n_93),
.B2(n_137),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_225),
.B1(n_119),
.B2(n_124),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_137),
.B1(n_131),
.B2(n_118),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_122),
.B(n_102),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_88),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_89),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_41),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_217),
.A2(n_47),
.B1(n_104),
.B2(n_116),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_219),
.C(n_218),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_15),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_245),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_225),
.C(n_223),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_244),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_42),
.C(n_76),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_248),
.B(n_243),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_9),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_228),
.B(n_238),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_250),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_233),
.B1(n_230),
.B2(n_91),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_254),
.C(n_32),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_242),
.A2(n_230),
.B1(n_70),
.B2(n_91),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_45),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_45),
.B1(n_88),
.B2(n_9),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_255),
.B(n_15),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_SL g262 ( 
.A(n_259),
.B(n_13),
.C(n_11),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_258),
.A2(n_13),
.B(n_32),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_0),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_266),
.B(n_264),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B(n_3),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_3),
.C(n_4),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_4),
.B(n_5),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_5),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_6),
.Y(n_273)
);


endmodule