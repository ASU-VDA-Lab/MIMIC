module fake_jpeg_26396_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_10),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_33),
.B1(n_30),
.B2(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_45),
.B1(n_43),
.B2(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_42),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_20),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_33),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_62),
.B(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_56),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_69),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_31),
.B1(n_24),
.B2(n_14),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_66),
.B1(n_51),
.B2(n_43),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_63),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_23),
.B(n_19),
.C(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_40),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_31),
.B1(n_19),
.B2(n_26),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_48),
.B1(n_14),
.B2(n_40),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_86),
.B1(n_66),
.B2(n_51),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_44),
.B1(n_45),
.B2(n_25),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_82),
.B(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_88),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_44),
.B1(n_25),
.B2(n_17),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_16),
.C(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_13),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_104),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_102),
.Y(n_120)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_51),
.B1(n_61),
.B2(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_99),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_72),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_50),
.B1(n_57),
.B2(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_106),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_62),
.B(n_67),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_54),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_62),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_12),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_85),
.C(n_89),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_98),
.B(n_96),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_105),
.C(n_97),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_119),
.C(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_107),
.B1(n_93),
.B2(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_88),
.C(n_75),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_75),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_84),
.C(n_80),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_121),
.C(n_117),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_109),
.C(n_94),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_136),
.C(n_124),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_29),
.B(n_4),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_106),
.C(n_74),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_127),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_120),
.B1(n_126),
.B2(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_148),
.B1(n_130),
.B2(n_133),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_113),
.B1(n_48),
.B2(n_29),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_128),
.Y(n_147)
);

AOI21x1_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_3),
.B(n_5),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.C(n_131),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_137),
.B1(n_128),
.B2(n_139),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_141),
.C(n_147),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_131),
.C(n_148),
.Y(n_158)
);

NOR2x1_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_140),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_161),
.A3(n_162),
.B1(n_158),
.B2(n_157),
.C1(n_3),
.C2(n_8),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_6),
.B(n_7),
.Y(n_166)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_11),
.CI(n_5),
.CON(n_162),
.SN(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_149),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_9),
.B(n_6),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_8),
.C(n_9),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_164),
.C(n_9),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_170),
.Y(n_172)
);


endmodule