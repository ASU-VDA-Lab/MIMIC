module real_jpeg_24319_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_258;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_257;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_37),
.B1(n_48),
.B2(n_50),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_22),
.B1(n_26),
.B2(n_37),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_54),
.B1(n_69),
.B2(n_83),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_6),
.A2(n_22),
.B1(n_26),
.B2(n_69),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_40),
.B1(n_54),
.B2(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_40),
.B1(n_48),
.B2(n_50),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_40),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_47),
.C(n_50),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_8),
.B(n_46),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_8),
.B(n_35),
.C(n_72),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_8),
.B(n_22),
.C(n_32),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_8),
.B(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_8),
.B(n_63),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_75),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_47),
.B1(n_51),
.B2(n_54),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_11),
.Y(n_162)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_116),
.B1(n_257),
.B2(n_258),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_14),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_115),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_97),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_16),
.B(n_97),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_58),
.Y(n_16)
);

AOI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B(n_43),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_18),
.A2(n_43),
.B1(n_44),
.B2(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_18),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_18),
.A2(n_29),
.B1(n_100),
.B2(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_20),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_21),
.A2(n_25),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_21),
.B(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_21),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_22),
.B(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_24),
.A2(n_105),
.B(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_24),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_28),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_29),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B(n_38),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_30),
.B(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_30),
.A2(n_38),
.B(n_132),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

OA22x2_ASAP7_75t_SL g74 ( 
.A1(n_34),
.A2(n_35),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_35),
.B(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_39),
.A2(n_41),
.B1(n_63),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_39),
.B(n_90),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_46),
.A2(n_52),
.B1(n_56),
.B2(n_112),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_50),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_50),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_56),
.Y(n_84)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_77),
.B2(n_78),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_61),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_66),
.A2(n_111),
.B1(n_121),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_66),
.B(n_175),
.C(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_66),
.A2(n_165),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_66),
.B(n_111),
.C(n_152),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_74),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_70),
.B(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_93),
.B(n_95),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_74),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_76),
.Y(n_135)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_113),
.C(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_79),
.A2(n_80),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_79),
.A2(n_80),
.B1(n_133),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_125),
.C(n_133),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_92),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.C(n_102),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_101),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_111),
.C(n_113),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_104),
.Y(n_248)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_108),
.A2(n_109),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_108),
.A2(n_109),
.B1(n_188),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_109),
.B(n_182),
.C(n_188),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_109),
.B(n_158),
.C(n_219),
.Y(n_223)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_113),
.A2(n_114),
.B1(n_148),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_113),
.A2(n_114),
.B1(n_131),
.B2(n_145),
.Y(n_225)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_114),
.B(n_131),
.C(n_226),
.Y(n_229)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_116),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_138),
.B(n_256),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_136),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_118),
.B(n_136),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_119),
.B(n_122),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_124),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_125),
.A2(n_126),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_131),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_160),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_131),
.A2(n_145),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_205),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_133),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_251),
.B(n_255),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_178),
.B(n_237),
.C(n_250),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_167),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_141),
.B(n_167),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_151),
.B2(n_166),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_144),
.B(n_150),
.C(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_164),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_157),
.A2(n_158),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_211),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_158)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_174),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_169),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_176),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_176),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_236),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_197),
.B(n_235),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_194),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_181),
.B(n_194),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_183),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_228),
.B(n_234),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_222),
.B(n_227),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_214),
.B(n_221),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_206),
.B(n_213),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_203),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_210),
.B(n_212),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_216),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_249),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_246),
.B2(n_247),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_247),
.C(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);


endmodule