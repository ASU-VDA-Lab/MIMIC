module fake_ariane_2811_n_1907 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1907);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1907;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_83),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_28),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_91),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_18),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_88),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_122),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_67),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_3),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_22),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_108),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_148),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_120),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_46),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_143),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_7),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_129),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_43),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_153),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_12),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_68),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_121),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_10),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_139),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_46),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_20),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_1),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_154),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_117),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_168),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_82),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_102),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_10),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_32),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_99),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_85),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_89),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_131),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_61),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_137),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_28),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_101),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_69),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_105),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_64),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_104),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_118),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_164),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_37),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_58),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_95),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_0),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_43),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_92),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_100),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_78),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_74),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_79),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_5),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_58),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_158),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_51),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_34),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_37),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_169),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_138),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_173),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_132),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_93),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_124),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_72),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_151),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_145),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_22),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_172),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_127),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_163),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_29),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_178),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_52),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_38),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_94),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_156),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_128),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_111),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_96),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_44),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_84),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_149),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_8),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_76),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_32),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_80),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_112),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_123),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_57),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_176),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_7),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_13),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_77),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_39),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_59),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_125),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_71),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_14),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_47),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_8),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_19),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_87),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_86),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_116),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_81),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_119),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_12),
.Y(n_339)
);

HB1xp67_ASAP7_75t_SL g340 ( 
.A(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_150),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_2),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_0),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_49),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_126),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_51),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_42),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_152),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_35),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_106),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_9),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_15),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_2),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_55),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_352),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_213),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_184),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_334),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_258),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_180),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_331),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_182),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_184),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_345),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_258),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_340),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_209),
.B(n_4),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_185),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_191),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_267),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_185),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_192),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_193),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_193),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_200),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_200),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_206),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_256),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_206),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_279),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_196),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_218),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_218),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_222),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_209),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_223),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_R g392 ( 
.A(n_223),
.B(n_177),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_222),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_241),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_197),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_241),
.B(n_6),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_244),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_186),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_186),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_244),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_205),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_245),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_183),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_245),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_246),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_246),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_247),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_247),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_352),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_189),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_250),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_208),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_250),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_186),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_220),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_252),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_252),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_258),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_269),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_269),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_282),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_258),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_224),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_225),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_227),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_276),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_282),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_283),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_283),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_287),
.B(n_6),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_230),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_219),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_231),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_232),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_287),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_237),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_292),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_219),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_238),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_243),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_251),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_219),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_292),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_309),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_257),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_368),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_419),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_398),
.B(n_294),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_398),
.B(n_294),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_361),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_371),
.B(n_258),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_423),
.A2(n_300),
.B(n_298),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_410),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_368),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_362),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_362),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_408),
.B(n_298),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_362),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_359),
.B(n_300),
.Y(n_468)
);

NAND2x1_ASAP7_75t_L g469 ( 
.A(n_359),
.B(n_228),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_366),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_366),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_372),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_427),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_376),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_378),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_390),
.A2(n_391),
.B1(n_367),
.B2(n_364),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_378),
.B(n_302),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_379),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_380),
.A2(n_382),
.B(n_381),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_408),
.B(n_384),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_387),
.A2(n_305),
.B(n_302),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_363),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_383),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_389),
.B(n_393),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_369),
.A2(n_315),
.B1(n_248),
.B2(n_239),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_394),
.B(n_305),
.Y(n_501)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_394),
.A2(n_312),
.B(n_306),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_358),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_402),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_404),
.B(n_279),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_306),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_404),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_365),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_405),
.B(n_279),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_310),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g518 ( 
.A(n_392),
.B(n_310),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_412),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_464),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_461),
.B(n_414),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_464),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_461),
.B(n_497),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_464),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_453),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_451),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_414),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_513),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_513),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_473),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_513),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_518),
.A2(n_396),
.B1(n_431),
.B2(n_262),
.Y(n_540)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_451),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_473),
.B(n_370),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_484),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_417),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g545 ( 
.A(n_496),
.B(n_374),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_513),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_482),
.B(n_373),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_493),
.B(n_377),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_489),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_418),
.C(n_417),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_513),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_513),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_513),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_L g557 ( 
.A(n_520),
.B(n_420),
.C(n_418),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_489),
.B(n_395),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_511),
.A2(n_433),
.B1(n_445),
.B2(n_415),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_497),
.B(n_420),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_459),
.A2(n_318),
.B(n_312),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_482),
.B(n_401),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_457),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_497),
.B(n_413),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_511),
.A2(n_439),
.B1(n_399),
.B2(n_443),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_497),
.B(n_228),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_523),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_497),
.B(n_421),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_490),
.B(n_416),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_486),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_457),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_523),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_486),
.B(n_421),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_457),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_457),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_510),
.B(n_422),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_484),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_523),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_453),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_523),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_479),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_490),
.B(n_425),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_514),
.B(n_426),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_523),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_453),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_523),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_523),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_496),
.B(n_440),
.Y(n_597)
);

OR2x6_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_385),
.Y(n_598)
);

BUFx8_ASAP7_75t_SL g599 ( 
.A(n_504),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_514),
.B(n_432),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_498),
.B(n_442),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_510),
.B(n_422),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_457),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_428),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_523),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_465),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_486),
.B(n_428),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_478),
.Y(n_613)
);

AOI21x1_ASAP7_75t_L g614 ( 
.A1(n_469),
.A2(n_430),
.B(n_429),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_465),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_505),
.B(n_429),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_465),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_465),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_492),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_520),
.B(n_434),
.Y(n_620)
);

INVx4_ASAP7_75t_SL g621 ( 
.A(n_505),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_465),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_492),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_465),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_510),
.B(n_515),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_462),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_505),
.B(n_435),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_498),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_478),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_484),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_484),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_462),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_459),
.A2(n_320),
.B1(n_261),
.B2(n_263),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_462),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_448),
.Y(n_636)
);

OAI21xp33_ASAP7_75t_L g637 ( 
.A1(n_470),
.A2(n_436),
.B(n_430),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_436),
.Y(n_638)
);

BUFx6f_ASAP7_75t_SL g639 ( 
.A(n_522),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_448),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_448),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_450),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_452),
.A2(n_278),
.B1(n_313),
.B2(n_265),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_450),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_450),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_520),
.B(n_441),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_515),
.B(n_438),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_522),
.B(n_446),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_520),
.B(n_438),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_522),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_454),
.B(n_403),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_468),
.A2(n_323),
.B1(n_355),
.B2(n_354),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_452),
.B(n_360),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_522),
.B(n_444),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_520),
.B(n_444),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_494),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_494),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_494),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_494),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_458),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_454),
.Y(n_663)
);

AND3x1_ASAP7_75t_L g664 ( 
.A(n_515),
.B(n_187),
.C(n_183),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_458),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_517),
.A2(n_353),
.B1(n_273),
.B2(n_350),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_468),
.B(n_187),
.Y(n_667)
);

BUFx4f_ASAP7_75t_L g668 ( 
.A(n_491),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_520),
.B(n_274),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_346),
.Y(n_670)
);

BUFx4f_ASAP7_75t_L g671 ( 
.A(n_491),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_458),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_508),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_508),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_508),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_456),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_562),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_626),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_562),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_663),
.B(n_508),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_526),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_L g682 ( 
.A(n_533),
.B(n_480),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_606),
.B(n_508),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_528),
.B(n_508),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_533),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_526),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_541),
.B(n_579),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_527),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_620),
.B(n_509),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_648),
.B(n_509),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_584),
.B(n_509),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_537),
.B(n_579),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_632),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_584),
.B(n_509),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_546),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_602),
.B(n_509),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_606),
.B(n_611),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_572),
.B(n_470),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_606),
.B(n_509),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_606),
.B(n_519),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_572),
.B(n_470),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_543),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_602),
.B(n_519),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_529),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_611),
.B(n_519),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_649),
.B(n_519),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_542),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_543),
.B(n_519),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_R g711 ( 
.A(n_545),
.B(n_519),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_540),
.A2(n_512),
.B1(n_469),
.B2(n_517),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_529),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_649),
.B(n_471),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_531),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_531),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_530),
.B(n_653),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_540),
.A2(n_524),
.B1(n_521),
.B2(n_474),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_632),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_558),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_611),
.B(n_471),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_645),
.A2(n_480),
.B1(n_501),
.B2(n_471),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_550),
.A2(n_517),
.B1(n_521),
.B2(n_524),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_611),
.B(n_474),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_635),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_653),
.B(n_474),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_566),
.B(n_475),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_SL g728 ( 
.A(n_552),
.B(n_475),
.Y(n_728)
);

AO21x2_ASAP7_75t_L g729 ( 
.A1(n_553),
.A2(n_501),
.B(n_336),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_589),
.B(n_475),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_552),
.B(n_481),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_544),
.B(n_481),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_628),
.A2(n_491),
.B1(n_502),
.B2(n_460),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_544),
.B(n_481),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_625),
.B(n_485),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_558),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_560),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_625),
.B(n_485),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_570),
.B(n_485),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_559),
.B(n_488),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_546),
.B(n_488),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_534),
.A2(n_524),
.B(n_521),
.C(n_516),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_589),
.B(n_488),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_651),
.B(n_495),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_546),
.B(n_495),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_609),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_546),
.B(n_495),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_670),
.B(n_499),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_560),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_664),
.B(n_499),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_543),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_563),
.A2(n_516),
.B(n_507),
.C(n_506),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_667),
.B(n_499),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_664),
.B(n_645),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_666),
.B(n_500),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_627),
.B(n_650),
.Y(n_758)
);

BUFx5_ASAP7_75t_L g759 ( 
.A(n_572),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_601),
.B(n_597),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_655),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_578),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_610),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_572),
.B(n_500),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_597),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_578),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_667),
.B(n_500),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_553),
.A2(n_516),
.B1(n_507),
.B2(n_506),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_578),
.A2(n_506),
.B1(n_503),
.B2(n_507),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_619),
.B(n_503),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_574),
.B(n_619),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_567),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_572),
.A2(n_502),
.B1(n_491),
.B2(n_460),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_561),
.B(n_503),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_599),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_619),
.B(n_472),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_610),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_619),
.B(n_472),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_668),
.A2(n_472),
.B(n_487),
.C(n_483),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_623),
.B(n_472),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_623),
.B(n_476),
.Y(n_781)
);

O2A1O1Ixp5_ASAP7_75t_L g782 ( 
.A1(n_669),
.A2(n_476),
.B(n_477),
.C(n_487),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_666),
.B(n_476),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_662),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_623),
.B(n_476),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_575),
.B(n_477),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_590),
.Y(n_787)
);

NAND2x1_ASAP7_75t_L g788 ( 
.A(n_592),
.B(n_477),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_623),
.B(n_477),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_634),
.B(n_483),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_601),
.A2(n_322),
.B1(n_310),
.B2(n_487),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_668),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_634),
.B(n_483),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_634),
.B(n_483),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_634),
.B(n_487),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_491),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_571),
.B(n_491),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_640),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_629),
.B(n_256),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_654),
.B(n_668),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_576),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_658),
.B(n_502),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_658),
.B(n_277),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_640),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_658),
.B(n_502),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_673),
.B(n_502),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_644),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_673),
.B(n_281),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_662),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_644),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_671),
.B(n_285),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_673),
.B(n_502),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_673),
.B(n_460),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_671),
.B(n_318),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_662),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_675),
.B(n_661),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_675),
.B(n_460),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_671),
.B(n_295),
.Y(n_818)
);

OAI221xp5_ASAP7_75t_L g819 ( 
.A1(n_633),
.A2(n_290),
.B1(n_304),
.B2(n_212),
.C(n_280),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_551),
.B(n_214),
.C(n_212),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_675),
.B(n_296),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_659),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_576),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_598),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_675),
.B(n_299),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_585),
.B(n_336),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_581),
.B(n_460),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_660),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_660),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_591),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_604),
.B(n_460),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_SL g833 ( 
.A1(n_629),
.A2(n_303),
.B1(n_301),
.B2(n_317),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_665),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_665),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_572),
.B(n_535),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_576),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_612),
.B(n_289),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_674),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_616),
.A2(n_322),
.B(n_239),
.C(n_249),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_661),
.B(n_326),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_638),
.B(n_308),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_572),
.B(n_535),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_535),
.B(n_330),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_775),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_687),
.B(n_598),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_759),
.B(n_585),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_747),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_717),
.B(n_726),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_697),
.B(n_639),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_759),
.B(n_585),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_756),
.A2(n_639),
.B1(n_600),
.B2(n_598),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_759),
.B(n_585),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_677),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_689),
.A2(n_532),
.B(n_525),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_677),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_796),
.A2(n_630),
.B(n_607),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_691),
.A2(n_532),
.B(n_525),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_802),
.A2(n_630),
.B(n_607),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_656),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_710),
.A2(n_817),
.B(n_813),
.Y(n_861)
);

NOR2x1p5_ASAP7_75t_L g862 ( 
.A(n_730),
.B(n_557),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_731),
.B(n_661),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_763),
.Y(n_864)
);

NAND2x1_ASAP7_75t_L g865 ( 
.A(n_801),
.B(n_592),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_777),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_731),
.A2(n_637),
.B(n_557),
.C(n_674),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_755),
.B(n_767),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_805),
.A2(n_630),
.B(n_607),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_685),
.B(n_652),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_680),
.B(n_652),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_739),
.A2(n_637),
.B(n_322),
.C(n_665),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_711),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_710),
.A2(n_532),
.B(n_525),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_824),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_694),
.B(n_613),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_787),
.B(n_652),
.Y(n_877)
);

O2A1O1Ixp5_ASAP7_75t_L g878 ( 
.A1(n_727),
.A2(n_800),
.B(n_818),
.C(n_811),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_679),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_831),
.B(n_607),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_760),
.B(n_598),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_806),
.A2(n_532),
.B(n_525),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_812),
.A2(n_587),
.B(n_549),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_722),
.B(n_630),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_786),
.A2(n_631),
.B(n_657),
.C(n_614),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_740),
.B(n_631),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_739),
.A2(n_740),
.B(n_841),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_837),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_683),
.A2(n_592),
.B1(n_631),
.B2(n_594),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_711),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_824),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_743),
.B(n_749),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_759),
.B(n_631),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_723),
.B(n_549),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_732),
.B(n_549),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_824),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_684),
.A2(n_587),
.B(n_549),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_765),
.B(n_598),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_744),
.A2(n_594),
.B(n_587),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_779),
.A2(n_538),
.B(n_536),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_683),
.A2(n_592),
.B1(n_594),
.B2(n_587),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_758),
.A2(n_639),
.B1(n_583),
.B2(n_582),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_827),
.A2(n_614),
.B(n_538),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_770),
.A2(n_304),
.B(n_325),
.C(n_329),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_776),
.A2(n_594),
.B(n_547),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_774),
.B(n_582),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_734),
.B(n_582),
.Y(n_907)
);

O2A1O1Ixp5_ASAP7_75t_L g908 ( 
.A1(n_721),
.A2(n_596),
.B(n_536),
.C(n_554),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_827),
.A2(n_782),
.B(n_769),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_681),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_681),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_797),
.B(n_583),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_761),
.B(n_583),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_778),
.A2(n_554),
.B(n_547),
.Y(n_914)
);

AOI33xp33_ASAP7_75t_L g915 ( 
.A1(n_791),
.A2(n_266),
.A3(n_339),
.B1(n_329),
.B2(n_325),
.B3(n_290),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_837),
.B(n_792),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_693),
.A2(n_577),
.B(n_608),
.C(n_615),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_825),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_735),
.B(n_568),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_738),
.B(n_568),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_686),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_798),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_780),
.A2(n_556),
.B(n_555),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_758),
.B(n_569),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_799),
.B(n_569),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_714),
.B(n_577),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_833),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_696),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_698),
.B(n_603),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_705),
.A2(n_603),
.B1(n_608),
.B2(n_615),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_781),
.A2(n_556),
.B(n_555),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_708),
.B(n_617),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_841),
.B(n_617),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_816),
.A2(n_618),
.B1(n_622),
.B2(n_624),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_709),
.B(n_618),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_792),
.Y(n_937)
);

HB1xp67_ASAP7_75t_SL g938 ( 
.A(n_820),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_686),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_741),
.B(n_621),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_699),
.B(n_622),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_751),
.A2(n_624),
.B(n_214),
.C(n_339),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_804),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_785),
.A2(n_573),
.B(n_564),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_759),
.B(n_535),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_814),
.A2(n_351),
.B(n_341),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_783),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_688),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_757),
.B(n_712),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_688),
.Y(n_950)
);

BUFx12f_ASAP7_75t_L g951 ( 
.A(n_792),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_814),
.A2(n_573),
.B(n_564),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_771),
.A2(n_819),
.B(n_718),
.C(n_724),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_807),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_803),
.B(n_808),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_790),
.A2(n_586),
.B(n_580),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_690),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_770),
.A2(n_586),
.B(n_580),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_803),
.A2(n_821),
.B(n_808),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_701),
.A2(n_249),
.B(n_266),
.C(n_280),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_746),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_793),
.A2(n_593),
.B(n_588),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_748),
.B(n_565),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_704),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_838),
.B(n_636),
.Y(n_965)
);

BUFx4f_ASAP7_75t_L g966 ( 
.A(n_792),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_794),
.A2(n_593),
.B(n_588),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_795),
.A2(n_596),
.B(n_595),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_801),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_842),
.B(n_636),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_690),
.Y(n_971)
);

AOI21xp33_ASAP7_75t_L g972 ( 
.A1(n_821),
.A2(n_565),
.B(n_641),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_706),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_759),
.B(n_535),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_810),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_702),
.A2(n_605),
.B(n_595),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_706),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_707),
.A2(n_605),
.B(n_548),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_704),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_826),
.B(n_816),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_704),
.B(n_752),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_789),
.A2(n_548),
.B(n_539),
.Y(n_982)
);

NAND2x1p5_ASAP7_75t_L g983 ( 
.A(n_704),
.B(n_641),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_752),
.B(n_539),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_789),
.A2(n_548),
.B(n_539),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_826),
.B(n_642),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_784),
.B(n_809),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_752),
.B(n_539),
.Y(n_988)
);

OAI321xp33_ASAP7_75t_L g989 ( 
.A1(n_840),
.A2(n_351),
.A3(n_341),
.B1(n_327),
.B2(n_203),
.C(n_335),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_828),
.A2(n_643),
.B(n_672),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_752),
.B(n_565),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_784),
.B(n_809),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_822),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_762),
.B(n_766),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_815),
.B(n_642),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_762),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_788),
.A2(n_548),
.B(n_539),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_823),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_548),
.B(n_676),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_700),
.A2(n_676),
.B(n_672),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_829),
.A2(n_643),
.B1(n_647),
.B2(n_646),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_729),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_762),
.B(n_256),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_SL g1004 ( 
.A1(n_830),
.A2(n_327),
.B(n_203),
.C(n_335),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_733),
.B(n_729),
.Y(n_1005)
);

AOI21xp33_ASAP7_75t_L g1006 ( 
.A1(n_742),
.A2(n_646),
.B(n_647),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_762),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_713),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_839),
.A2(n_348),
.B(n_332),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_815),
.B(n_621),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_834),
.B(n_621),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_678),
.A2(n_343),
.B1(n_347),
.B2(n_344),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_692),
.Y(n_1013)
);

NAND2x1p5_ASAP7_75t_L g1014 ( 
.A(n_766),
.B(n_621),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_695),
.A2(n_455),
.B(n_447),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_703),
.A2(n_676),
.B(n_455),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_764),
.A2(n_676),
.B(n_455),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_773),
.A2(n_676),
.B(n_455),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_719),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_766),
.B(n_621),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_728),
.A2(n_338),
.B1(n_356),
.B2(n_349),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_725),
.A2(n_260),
.B(n_228),
.C(n_235),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_834),
.A2(n_676),
.B(n_449),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_766),
.B(n_235),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_835),
.A2(n_843),
.B(n_836),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_768),
.B(n_309),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_835),
.A2(n_447),
.B(n_449),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_773),
.A2(n_449),
.B(n_447),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_733),
.A2(n_745),
.B1(n_844),
.B2(n_753),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_713),
.A2(n_447),
.B(n_449),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_772),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_SL g1032 ( 
.A(n_754),
.B(n_256),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_848),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_849),
.B(n_715),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_980),
.A2(n_772),
.B(n_753),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_887),
.A2(n_750),
.B(n_737),
.C(n_736),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_892),
.B(n_715),
.Y(n_1037)
);

AND2x2_ASAP7_75t_SL g1038 ( 
.A(n_949),
.B(n_235),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_928),
.A2(n_750),
.B1(n_737),
.B2(n_736),
.C(n_720),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_901),
.A2(n_720),
.B(n_716),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_876),
.B(n_716),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_868),
.A2(n_959),
.B(n_904),
.C(n_955),
.Y(n_1042)
);

O2A1O1Ixp5_ASAP7_75t_L g1043 ( 
.A1(n_878),
.A2(n_260),
.B(n_195),
.C(n_255),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_873),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_929),
.B(n_11),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_951),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_846),
.B(n_309),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_864),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_863),
.A2(n_260),
.B1(n_255),
.B2(n_195),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_986),
.A2(n_463),
.B(n_456),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_964),
.B(n_845),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_1007),
.B(n_456),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_929),
.B(n_11),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_1009),
.B(n_194),
.C(n_342),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_904),
.A2(n_953),
.B(n_1032),
.C(n_1004),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_866),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_939),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_939),
.Y(n_1058)
);

OR2x6_ASAP7_75t_SL g1059 ( 
.A(n_1012),
.B(n_179),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_948),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_862),
.B(n_13),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_966),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_909),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1007),
.B(n_456),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_966),
.B(n_181),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_1007),
.B(n_902),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_850),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_884),
.A2(n_199),
.B(n_337),
.C(n_333),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_890),
.B(n_16),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_881),
.B(n_19),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_906),
.B(n_21),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_877),
.B(n_21),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_877),
.B(n_24),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_846),
.B(n_24),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1026),
.A2(n_1005),
.B1(n_1019),
.B2(n_1013),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_937),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_925),
.B(n_25),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_894),
.A2(n_202),
.B1(n_328),
.B2(n_324),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_891),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1004),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_925),
.B(n_26),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_SL g1082 ( 
.A(n_852),
.B(n_201),
.C(n_321),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_880),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_1083)
);

AO21x1_ASAP7_75t_L g1084 ( 
.A1(n_963),
.A2(n_175),
.B(n_166),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_861),
.A2(n_210),
.B(n_319),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_870),
.B(n_33),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_922),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_899),
.A2(n_207),
.B(n_316),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_1007),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_846),
.B(n_33),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_870),
.B(n_34),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_898),
.B(n_35),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_994),
.B(n_456),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_918),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_913),
.B(n_36),
.Y(n_1095)
);

BUFx2_ASAP7_75t_L g1096 ( 
.A(n_918),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_889),
.A2(n_211),
.B(n_314),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_L g1098 ( 
.A1(n_984),
.A2(n_36),
.B(n_40),
.C(n_41),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_943),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_948),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_850),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_954),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_994),
.B(n_456),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_915),
.A2(n_215),
.B(n_311),
.C(n_307),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_975),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_915),
.B(n_40),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_957),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_886),
.A2(n_204),
.B1(n_297),
.B2(n_293),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_855),
.A2(n_198),
.B(n_291),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_936),
.B(n_45),
.Y(n_1110)
);

AOI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_880),
.A2(n_190),
.B(n_288),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_924),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_957),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_885),
.A2(n_188),
.B(n_286),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_936),
.B(n_47),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_867),
.A2(n_217),
.B(n_284),
.C(n_275),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_971),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_934),
.A2(n_48),
.B(n_50),
.C(n_53),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_926),
.B(n_48),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_858),
.A2(n_253),
.B(n_226),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_924),
.B(n_996),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_891),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_867),
.A2(n_254),
.B(n_229),
.C(n_272),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_924),
.B(n_456),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_938),
.A2(n_268),
.B1(n_233),
.B2(n_234),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1031),
.Y(n_1126)
);

NOR2x1_ASAP7_75t_L g1127 ( 
.A(n_896),
.B(n_463),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_926),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_961),
.B(n_50),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_993),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_937),
.B(n_463),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_896),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_924),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_895),
.A2(n_259),
.B(n_236),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_996),
.B(n_456),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_856),
.Y(n_1136)
);

CKINVDCx6p67_ASAP7_75t_R g1137 ( 
.A(n_1026),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_SL g1138 ( 
.A1(n_941),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_979),
.B(n_456),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_998),
.B(n_54),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1014),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_979),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_888),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_971),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_960),
.A2(n_56),
.B(n_59),
.C(n_61),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_888),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_958),
.A2(n_56),
.B(n_66),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_875),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_965),
.B(n_271),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1003),
.B(n_270),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_947),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_875),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_984),
.A2(n_463),
.B(n_264),
.C(n_242),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_856),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_907),
.A2(n_240),
.B1(n_221),
.B2(n_463),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_860),
.B(n_463),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_970),
.B(n_463),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_919),
.B(n_463),
.Y(n_1158)
);

BUFx12f_ASAP7_75t_L g1159 ( 
.A(n_916),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_969),
.B(n_463),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_SL g1161 ( 
.A1(n_1024),
.A2(n_90),
.B(n_98),
.C(n_103),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_910),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_941),
.B(n_107),
.C(n_130),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_969),
.B(n_134),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_916),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_911),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_882),
.A2(n_136),
.B(n_141),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_942),
.A2(n_142),
.B(n_155),
.C(n_160),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1025),
.B(n_161),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1006),
.A2(n_1001),
.B(n_872),
.C(n_920),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_872),
.A2(n_989),
.B(n_963),
.C(n_990),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1021),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_927),
.A2(n_935),
.B(n_930),
.C(n_933),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_921),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_912),
.B(n_879),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_950),
.B(n_973),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_883),
.A2(n_897),
.B(n_999),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_879),
.B(n_854),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_983),
.B(n_869),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_871),
.A2(n_859),
.B1(n_857),
.B2(n_1029),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_977),
.B(n_1008),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_991),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_983),
.B(n_991),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_987),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_1020),
.B(n_903),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_981),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_995),
.A2(n_992),
.B1(n_865),
.B2(n_931),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_940),
.B(n_1028),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1014),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1062),
.B(n_1079),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_1062),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1073),
.A2(n_1038),
.B1(n_1081),
.B2(n_1077),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1180),
.A2(n_985),
.B(n_982),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1079),
.B(n_940),
.Y(n_1194)
);

NAND3x1_ASAP7_75t_L g1195 ( 
.A(n_1090),
.B(n_1074),
.C(n_1061),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_L g1196 ( 
.A1(n_1042),
.A2(n_972),
.B1(n_1022),
.B2(n_946),
.C(n_917),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1177),
.A2(n_974),
.B(n_945),
.Y(n_1197)
);

NAND2x1_ASAP7_75t_L g1198 ( 
.A(n_1143),
.B(n_997),
.Y(n_1198)
);

AO32x2_ASAP7_75t_L g1199 ( 
.A1(n_1049),
.A2(n_1002),
.A3(n_1024),
.B1(n_1015),
.B2(n_900),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1173),
.A2(n_945),
.B(n_974),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1073),
.A2(n_874),
.B(n_908),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1051),
.Y(n_1202)
);

A2O1A1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1055),
.A2(n_1020),
.B(n_981),
.C(n_1000),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1036),
.A2(n_1010),
.A3(n_1011),
.B(n_1023),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1033),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_SL g1206 ( 
.A1(n_1116),
.A2(n_988),
.B(n_851),
.C(n_853),
.Y(n_1206)
);

AOI31xp67_ASAP7_75t_L g1207 ( 
.A1(n_1169),
.A2(n_988),
.A3(n_851),
.B(n_853),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1036),
.A2(n_962),
.A3(n_967),
.B(n_956),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1050),
.A2(n_968),
.B(n_914),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_SL g1210 ( 
.A1(n_1083),
.A2(n_952),
.B(n_978),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_893),
.C(n_847),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1172),
.A2(n_847),
.B1(n_893),
.B2(n_905),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1187),
.A2(n_923),
.B(n_932),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1187),
.A2(n_1169),
.B(n_1040),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1179),
.A2(n_944),
.B(n_976),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_SL g1216 ( 
.A(n_1051),
.B(n_1119),
.C(n_1118),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1179),
.A2(n_1170),
.B(n_1035),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1111),
.A2(n_1027),
.B(n_1030),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1171),
.A2(n_1016),
.A3(n_1017),
.B(n_1084),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1138),
.A2(n_1110),
.B(n_1115),
.C(n_1116),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1046),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_1044),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1138),
.A2(n_1123),
.B(n_1068),
.C(n_1129),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1189),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1123),
.A2(n_1068),
.B(n_1129),
.C(n_1072),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1034),
.A2(n_1037),
.B(n_1092),
.C(n_1171),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1034),
.A2(n_1158),
.B(n_1085),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1046),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1066),
.A2(n_1183),
.B(n_1103),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1147),
.B(n_1054),
.C(n_1145),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_1122),
.B(n_1041),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1128),
.B(n_1059),
.Y(n_1232)
);

AOI221x1_ASAP7_75t_L g1233 ( 
.A1(n_1114),
.A2(n_1104),
.B1(n_1086),
.B2(n_1091),
.C(n_1090),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1161),
.A2(n_1043),
.B(n_1167),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1124),
.A2(n_1037),
.B(n_1157),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1151),
.B(n_1182),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1066),
.A2(n_1183),
.B(n_1103),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1093),
.A2(n_1124),
.B(n_1127),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1126),
.B(n_1092),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1141),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1157),
.A2(n_1164),
.B(n_1160),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1168),
.A2(n_1080),
.B(n_1104),
.C(n_1082),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1069),
.A2(n_1045),
.B(n_1053),
.C(n_1063),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1071),
.A2(n_1095),
.B(n_1039),
.C(n_1097),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1065),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1093),
.A2(n_1064),
.B(n_1052),
.Y(n_1246)
);

AO22x2_ASAP7_75t_L g1247 ( 
.A1(n_1047),
.A2(n_1188),
.B1(n_1174),
.B2(n_1166),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1159),
.B(n_1101),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1126),
.B(n_1137),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1052),
.A2(n_1064),
.B(n_1175),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1136),
.A2(n_1156),
.A3(n_1117),
.B(n_1100),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1125),
.A2(n_1150),
.B1(n_1070),
.B2(n_1186),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1048),
.B(n_1099),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1163),
.A2(n_1149),
.B(n_1106),
.C(n_1098),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1164),
.A2(n_1160),
.B(n_1156),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_1153),
.B(n_1139),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1108),
.A2(n_1078),
.B(n_1134),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1139),
.A2(n_1135),
.B(n_1155),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1047),
.A2(n_1162),
.B1(n_1184),
.B2(n_1102),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1065),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1056),
.A2(n_1130),
.B(n_1105),
.C(n_1087),
.Y(n_1261)
);

AO32x2_ASAP7_75t_L g1262 ( 
.A1(n_1146),
.A2(n_1089),
.A3(n_1143),
.B1(n_1075),
.B2(n_1152),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1121),
.A2(n_1135),
.B(n_1131),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1067),
.A2(n_1140),
.B1(n_1075),
.B2(n_1132),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1136),
.A2(n_1057),
.A3(n_1058),
.B(n_1060),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_1107),
.A2(n_1144),
.B1(n_1113),
.B2(n_1154),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1088),
.A2(n_1120),
.B(n_1109),
.C(n_1148),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1122),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_SL g1269 ( 
.A1(n_1148),
.A2(n_1076),
.B(n_1165),
.C(n_1178),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1112),
.A2(n_1133),
.B(n_1131),
.Y(n_1270)
);

AND2x6_ASAP7_75t_L g1271 ( 
.A(n_1141),
.B(n_1076),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_R g1272 ( 
.A(n_1142),
.B(n_1152),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1112),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1185),
.A2(n_1176),
.B(n_1181),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1133),
.B(n_1142),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1133),
.A2(n_1142),
.B(n_1141),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1185),
.A2(n_756),
.B(n_887),
.C(n_566),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1142),
.A2(n_887),
.B(n_1042),
.C(n_1055),
.Y(n_1279)
);

CKINVDCx9p33_ASAP7_75t_R g1280 ( 
.A(n_1141),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1041),
.B(n_876),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1094),
.B(n_876),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_849),
.B2(n_892),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_849),
.B2(n_892),
.Y(n_1284)
);

AO32x2_ASAP7_75t_L g1285 ( 
.A1(n_1180),
.A2(n_1002),
.A3(n_1049),
.B1(n_718),
.B2(n_498),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1073),
.A2(n_887),
.B(n_959),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1126),
.Y(n_1289)
);

AOI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1050),
.A2(n_1177),
.B(n_1180),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1291)
);

AOI221x1_ASAP7_75t_L g1292 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_1123),
.B2(n_1116),
.C(n_1171),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1073),
.A2(n_756),
.B(n_887),
.C(n_566),
.Y(n_1293)
);

AOI31xp67_ASAP7_75t_L g1294 ( 
.A1(n_1169),
.A2(n_1179),
.A3(n_1103),
.B(n_1093),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1172),
.A2(n_928),
.B1(n_566),
.B2(n_550),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1051),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1041),
.B(n_876),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1180),
.A2(n_1036),
.A3(n_1171),
.B(n_991),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1033),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1041),
.B(n_876),
.Y(n_1301)
);

INVx4_ASAP7_75t_L g1302 ( 
.A(n_1062),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1172),
.B(n_504),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1062),
.B(n_1046),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1034),
.A2(n_887),
.B(n_1042),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1073),
.A2(n_887),
.B(n_959),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1041),
.B(n_876),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1073),
.A2(n_887),
.B(n_959),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1096),
.Y(n_1309)
);

OA22x2_ASAP7_75t_L g1310 ( 
.A1(n_1172),
.A2(n_478),
.B1(n_358),
.B2(n_928),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_SL g1311 ( 
.A(n_1062),
.B(n_687),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1046),
.B(n_846),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1062),
.B(n_1079),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1116),
.A2(n_699),
.B(n_1123),
.C(n_887),
.Y(n_1314)
);

OAI22x1_ASAP7_75t_L g1315 ( 
.A1(n_1090),
.A2(n_628),
.B1(n_756),
.B2(n_1182),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_849),
.B2(n_892),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1094),
.B(n_876),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1051),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1041),
.B(n_876),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_849),
.B2(n_892),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1172),
.B(n_504),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1073),
.A2(n_887),
.B(n_959),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1177),
.A2(n_1050),
.B(n_1169),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1177),
.A2(n_1050),
.B(n_1169),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1325)
);

OA21x2_ASAP7_75t_L g1326 ( 
.A1(n_1177),
.A2(n_1171),
.B(n_959),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1177),
.A2(n_1050),
.B(n_1169),
.Y(n_1327)
);

AO32x2_ASAP7_75t_L g1328 ( 
.A1(n_1180),
.A2(n_1002),
.A3(n_1049),
.B1(n_718),
.B2(n_498),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1096),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1177),
.A2(n_1050),
.B(n_1169),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1033),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1059),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1055),
.A2(n_1042),
.B(n_1119),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1062),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1073),
.A2(n_887),
.B1(n_849),
.B2(n_892),
.Y(n_1336)
);

NAND2x1_ASAP7_75t_L g1337 ( 
.A(n_1143),
.B(n_1089),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1073),
.A2(n_887),
.B(n_959),
.Y(n_1338)
);

AO32x2_ASAP7_75t_L g1339 ( 
.A1(n_1180),
.A2(n_1002),
.A3(n_1049),
.B1(n_718),
.B2(n_498),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1177),
.A2(n_1050),
.B(n_1169),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1051),
.Y(n_1341)
);

BUFx8_ASAP7_75t_L g1342 ( 
.A(n_1096),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1172),
.B(n_504),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1180),
.A2(n_959),
.B(n_980),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1033),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1192),
.A2(n_1316),
.B1(n_1320),
.B2(n_1283),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1237),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1310),
.A2(n_1315),
.B1(n_1336),
.B2(n_1284),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1191),
.B(n_1334),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1281),
.B(n_1297),
.Y(n_1350)
);

INVx6_ASAP7_75t_L g1351 ( 
.A(n_1191),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1289),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1282),
.B(n_1317),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1295),
.A2(n_1287),
.B1(n_1322),
.B2(n_1306),
.Y(n_1354)
);

INVx8_ASAP7_75t_L g1355 ( 
.A(n_1271),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1332),
.A2(n_1338),
.B1(n_1308),
.B2(n_1319),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1222),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1301),
.A2(n_1307),
.B1(n_1216),
.B2(n_1230),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1205),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1342),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1296),
.Y(n_1361)
);

BUFx8_ASAP7_75t_SL g1362 ( 
.A(n_1202),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1333),
.A2(n_1252),
.B1(n_1232),
.B2(n_1239),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1293),
.A2(n_1226),
.B1(n_1254),
.B2(n_1278),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1341),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1334),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1303),
.A2(n_1321),
.B1(n_1343),
.B2(n_1242),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1248),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1318),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1273),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1342),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1300),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1236),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1331),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1249),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1345),
.Y(n_1376)
);

CKINVDCx11_ASAP7_75t_R g1377 ( 
.A(n_1245),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1260),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1261),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1259),
.A2(n_1247),
.B1(n_1326),
.B2(n_1195),
.Y(n_1380)
);

INVx1_ASAP7_75t_SL g1381 ( 
.A(n_1309),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1259),
.A2(n_1247),
.B1(n_1326),
.B2(n_1285),
.Y(n_1382)
);

AOI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1264),
.A2(n_1311),
.B1(n_1231),
.B2(n_1312),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1265),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1285),
.A2(n_1328),
.B1(n_1339),
.B2(n_1292),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1221),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1265),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1228),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1225),
.A2(n_1344),
.B1(n_1335),
.B2(n_1286),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_SL g1390 ( 
.A1(n_1285),
.A2(n_1339),
.B1(n_1328),
.B2(n_1298),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1231),
.A2(n_1312),
.B1(n_1313),
.B2(n_1190),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1329),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1268),
.Y(n_1393)
);

INVx6_ASAP7_75t_L g1394 ( 
.A(n_1302),
.Y(n_1394)
);

CKINVDCx14_ASAP7_75t_R g1395 ( 
.A(n_1248),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1271),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1190),
.Y(n_1397)
);

INVxp67_ASAP7_75t_L g1398 ( 
.A(n_1276),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1196),
.A2(n_1257),
.B1(n_1291),
.B2(n_1288),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1325),
.A2(n_1274),
.B1(n_1194),
.B2(n_1227),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1328),
.A2(n_1339),
.B1(n_1305),
.B2(n_1201),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1266),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1266),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1224),
.Y(n_1404)
);

BUFx10_ASAP7_75t_L g1405 ( 
.A(n_1194),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1214),
.A2(n_1235),
.B1(n_1212),
.B2(n_1217),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1233),
.A2(n_1223),
.B1(n_1299),
.B2(n_1279),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1271),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1280),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1251),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1271),
.B1(n_1302),
.B2(n_1255),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1299),
.A2(n_1262),
.B1(n_1314),
.B2(n_1244),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_L g1413 ( 
.A(n_1304),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1262),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1299),
.A2(n_1262),
.B1(n_1200),
.B2(n_1213),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1240),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1272),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1241),
.A2(n_1258),
.B1(n_1218),
.B2(n_1250),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1243),
.A2(n_1220),
.B1(n_1193),
.B2(n_1215),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1275),
.B(n_1277),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1337),
.B(n_1263),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1211),
.A2(n_1210),
.B1(n_1269),
.B2(n_1206),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1270),
.B(n_1229),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1238),
.B(n_1246),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1256),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1198),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1234),
.A2(n_1197),
.B1(n_1209),
.B2(n_1199),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1323),
.B(n_1340),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1294),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1203),
.B(n_1219),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1199),
.A2(n_1327),
.B1(n_1324),
.B2(n_1330),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1267),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1290),
.A2(n_1207),
.B1(n_1219),
.B2(n_1199),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1204),
.A2(n_1038),
.B1(n_478),
.B2(n_1192),
.Y(n_1434)
);

INVx8_ASAP7_75t_L g1435 ( 
.A(n_1208),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1253),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1295),
.A2(n_1283),
.B1(n_1316),
.B2(n_1284),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1253),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1192),
.A2(n_1038),
.B1(n_478),
.B2(n_1310),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1273),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1281),
.B(n_1297),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1332),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1332),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1332),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1192),
.A2(n_1038),
.B1(n_628),
.B2(n_360),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1192),
.A2(n_1038),
.B1(n_478),
.B2(n_1310),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1192),
.A2(n_1038),
.B1(n_478),
.B2(n_1310),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1192),
.A2(n_1038),
.B1(n_478),
.B2(n_1310),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1224),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_1202),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1253),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1253),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1253),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1342),
.Y(n_1454)
);

CKINVDCx6p67_ASAP7_75t_R g1455 ( 
.A(n_1332),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1253),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1282),
.B(n_1317),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1253),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1202),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1202),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1273),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1295),
.A2(n_1343),
.B1(n_1321),
.B2(n_1303),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1295),
.A2(n_1192),
.B1(n_1284),
.B2(n_1283),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1191),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1342),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1237),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1295),
.A2(n_1192),
.B1(n_1284),
.B2(n_1283),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1342),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1295),
.A2(n_1293),
.B(n_1192),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1281),
.B(n_1297),
.Y(n_1470)
);

CKINVDCx9p33_ASAP7_75t_R g1471 ( 
.A(n_1280),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1384),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1387),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1426),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1410),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1426),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1389),
.A2(n_1433),
.B(n_1364),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1428),
.A2(n_1419),
.B(n_1431),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1426),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1429),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1420),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1424),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1347),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1353),
.B(n_1457),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1428),
.A2(n_1419),
.B(n_1431),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1352),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1396),
.B(n_1408),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1466),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1352),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1466),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1423),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1359),
.Y(n_1492)
);

INVx5_ASAP7_75t_L g1493 ( 
.A(n_1355),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1425),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1372),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1432),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1427),
.A2(n_1418),
.B(n_1406),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1374),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1376),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1435),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1430),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1414),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1401),
.B(n_1390),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1402),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1403),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1398),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1398),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1379),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1382),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1382),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1437),
.A2(n_1463),
.B(n_1467),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1421),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_SL g1513 ( 
.A1(n_1346),
.A2(n_1469),
.B(n_1399),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1415),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1415),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1390),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1436),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1357),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1438),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1427),
.A2(n_1406),
.B(n_1418),
.Y(n_1520)
);

INVx1_ASAP7_75t_SL g1521 ( 
.A(n_1361),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1471),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1462),
.B(n_1367),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1385),
.B(n_1346),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1351),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1416),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1451),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1445),
.A2(n_1446),
.B1(n_1439),
.B2(n_1447),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1456),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1458),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1437),
.A2(n_1422),
.B(n_1354),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1416),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1412),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1354),
.A2(n_1399),
.B(n_1356),
.C(n_1348),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1412),
.Y(n_1536)
);

AO21x2_ASAP7_75t_L g1537 ( 
.A1(n_1383),
.A2(n_1385),
.B(n_1350),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1373),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1400),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1400),
.B(n_1391),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1407),
.B(n_1434),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1380),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1411),
.A2(n_1349),
.B(n_1363),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1380),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1411),
.A2(n_1363),
.B(n_1358),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1369),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1393),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1375),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1441),
.B(n_1470),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_SL g1550 ( 
.A(n_1366),
.B(n_1417),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1407),
.Y(n_1551)
);

CKINVDCx6p67_ASAP7_75t_R g1552 ( 
.A(n_1442),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1392),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1358),
.B(n_1381),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1356),
.B(n_1440),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1397),
.B(n_1448),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1501),
.B(n_1445),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1501),
.B(n_1417),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1449),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1484),
.B(n_1440),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1484),
.B(n_1440),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1541),
.B(n_1461),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1511),
.B(n_1368),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1480),
.B(n_1461),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1404),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1480),
.B(n_1461),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1486),
.B(n_1370),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1511),
.B(n_1370),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1535),
.A2(n_1409),
.B(n_1413),
.C(n_1395),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1496),
.B(n_1370),
.Y(n_1570)
);

AO32x2_ASAP7_75t_L g1571 ( 
.A1(n_1481),
.A2(n_1479),
.A3(n_1474),
.B1(n_1476),
.B2(n_1525),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1513),
.A2(n_1360),
.B(n_1468),
.C(n_1465),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1541),
.A2(n_1455),
.B1(n_1443),
.B2(n_1444),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1529),
.A2(n_1413),
.B(n_1454),
.C(n_1386),
.Y(n_1574)
);

AOI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1524),
.A2(n_1513),
.B1(n_1503),
.B2(n_1551),
.C(n_1496),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1489),
.B(n_1460),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1477),
.A2(n_1460),
.B(n_1371),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1540),
.B(n_1464),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1524),
.A2(n_1459),
.B(n_1365),
.C(n_1450),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_SL g1580 ( 
.A1(n_1550),
.A2(n_1377),
.B(n_1378),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1518),
.B(n_1388),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1545),
.A2(n_1394),
.B1(n_1464),
.B2(n_1405),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1489),
.B(n_1362),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1532),
.B(n_1394),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1553),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1522),
.B(n_1394),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1547),
.Y(n_1587)
);

CKINVDCx6p67_ASAP7_75t_R g1588 ( 
.A(n_1552),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1503),
.A2(n_1551),
.B1(n_1532),
.B2(n_1514),
.C(n_1515),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1552),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1555),
.A2(n_1540),
.B(n_1514),
.C(n_1515),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1521),
.B(n_1546),
.Y(n_1592)
);

AO21x1_ASAP7_75t_L g1593 ( 
.A1(n_1554),
.A2(n_1536),
.B(n_1534),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1508),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1481),
.B(n_1506),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1492),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1555),
.B(n_1548),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1540),
.A2(n_1539),
.B(n_1543),
.C(n_1542),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1532),
.B(n_1522),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1540),
.A2(n_1543),
.B(n_1544),
.C(n_1516),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1507),
.B(n_1500),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1491),
.B(n_1517),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1545),
.A2(n_1537),
.B1(n_1509),
.B2(n_1510),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1526),
.A2(n_1533),
.B(n_1538),
.C(n_1495),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1545),
.B(n_1477),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1549),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1487),
.Y(n_1607)
);

O2A1O1Ixp33_ASAP7_75t_SL g1608 ( 
.A1(n_1526),
.A2(n_1533),
.B(n_1499),
.C(n_1498),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1487),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1545),
.A2(n_1497),
.B(n_1520),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1509),
.A2(n_1510),
.B1(n_1491),
.B2(n_1527),
.C(n_1519),
.Y(n_1611)
);

CKINVDCx20_ASAP7_75t_R g1612 ( 
.A(n_1549),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1497),
.A2(n_1485),
.B(n_1478),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1556),
.A2(n_1512),
.B(n_1478),
.C(n_1485),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1594),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1594),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1482),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1596),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1483),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1609),
.B(n_1520),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1575),
.A2(n_1520),
.B1(n_1556),
.B2(n_1493),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1571),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1605),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1605),
.B(n_1599),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1610),
.B(n_1520),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1580),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1530),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1595),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1494),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1613),
.B(n_1494),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1602),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1571),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1559),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1571),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1565),
.B(n_1512),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1575),
.A2(n_1537),
.B1(n_1504),
.B2(n_1505),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1559),
.B(n_1488),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1557),
.A2(n_1505),
.B1(n_1504),
.B2(n_1528),
.Y(n_1639)
);

AND2x4_ASAP7_75t_SL g1640 ( 
.A(n_1578),
.B(n_1583),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1571),
.B(n_1490),
.Y(n_1641)
);

INVxp67_ASAP7_75t_SL g1642 ( 
.A(n_1584),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1589),
.A2(n_1537),
.B1(n_1531),
.B2(n_1502),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1563),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1601),
.B(n_1597),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1558),
.B(n_1502),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1629),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1644),
.B(n_1565),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1644),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1629),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1614),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1622),
.B(n_1598),
.Y(n_1655)
);

AOI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1623),
.A2(n_1589),
.B1(n_1557),
.B2(n_1593),
.C(n_1611),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1631),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1558),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1624),
.A2(n_1611),
.B1(n_1563),
.B2(n_1579),
.C(n_1600),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1606),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1633),
.B(n_1585),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1629),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1640),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1630),
.B(n_1603),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1633),
.A2(n_1582),
.B(n_1577),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1633),
.B(n_1576),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1620),
.B(n_1617),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1640),
.Y(n_1669)
);

AO21x2_ASAP7_75t_L g1670 ( 
.A1(n_1621),
.A2(n_1591),
.B(n_1582),
.Y(n_1670)
);

AO21x2_ASAP7_75t_L g1671 ( 
.A1(n_1621),
.A2(n_1472),
.B(n_1473),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1560),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1631),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1626),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1637),
.A2(n_1612),
.B1(n_1562),
.B2(n_1569),
.Y(n_1676)
);

OAI31xp33_ASAP7_75t_L g1677 ( 
.A1(n_1637),
.A2(n_1574),
.A3(n_1572),
.B(n_1564),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1561),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1625),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1618),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1641),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1635),
.B(n_1577),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1635),
.B(n_1566),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1632),
.B(n_1567),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1618),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1638),
.B(n_1475),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1680),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1657),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1664),
.B(n_1646),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1650),
.B(n_1615),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1651),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1657),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1664),
.B(n_1646),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1673),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1664),
.B(n_1646),
.Y(n_1696)
);

OR2x6_ASAP7_75t_L g1697 ( 
.A(n_1654),
.B(n_1578),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1669),
.B(n_1628),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1650),
.B(n_1615),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1680),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1659),
.B(n_1616),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1680),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1685),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1667),
.B(n_1638),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1667),
.B(n_1638),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1659),
.B(n_1616),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1651),
.B(n_1640),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1667),
.B(n_1627),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1651),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1656),
.A2(n_1643),
.B1(n_1625),
.B2(n_1562),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1685),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1659),
.B(n_1627),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1661),
.B(n_1588),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1658),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1686),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1656),
.A2(n_1643),
.B1(n_1642),
.B2(n_1639),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1686),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1662),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1684),
.B(n_1647),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1662),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1679),
.B(n_1619),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1688),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1688),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1695),
.B(n_1673),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1722),
.B(n_1709),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1653),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1711),
.A2(n_1573),
.B1(n_1590),
.B2(n_1583),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1687),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1716),
.B(n_1661),
.Y(n_1734)
);

NOR2xp67_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1700),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1700),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1710),
.B(n_1653),
.Y(n_1740)
);

NOR2x1_ASAP7_75t_R g1741 ( 
.A(n_1692),
.B(n_1626),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1691),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1702),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1687),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1708),
.B(n_1675),
.Y(n_1746)
);

AOI21xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1724),
.A2(n_1669),
.B(n_1648),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1724),
.B(n_1675),
.Y(n_1748)
);

OAI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1697),
.A2(n_1676),
.B1(n_1660),
.B2(n_1655),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1697),
.B(n_1676),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1692),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1703),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1724),
.B(n_1675),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1703),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1706),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1706),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1713),
.Y(n_1758)
);

OR2x6_ASAP7_75t_L g1759 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1713),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1711),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1718),
.B(n_1655),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1692),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1718),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1690),
.B(n_1675),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1720),
.B(n_1655),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1720),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1725),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1755),
.B(n_1729),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1726),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1726),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1751),
.B(n_1690),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1751),
.B(n_1694),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1730),
.B(n_1704),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1694),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1761),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1733),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1748),
.B(n_1696),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1728),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1730),
.B(n_1762),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1749),
.B(n_1675),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1654),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1728),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1753),
.B(n_1696),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1763),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1753),
.B(n_1698),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1766),
.B(n_1679),
.Y(n_1787)
);

INVxp33_ASAP7_75t_L g1788 ( 
.A(n_1741),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1727),
.B(n_1738),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1736),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1768),
.B(n_1704),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1763),
.B(n_1679),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1679),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1705),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1736),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1675),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1727),
.B(n_1698),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1738),
.B(n_1668),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1746),
.B(n_1765),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1764),
.B(n_1705),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1732),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1734),
.B(n_1581),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_L g1803 ( 
.A(n_1731),
.B(n_1592),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1764),
.B(n_1682),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1769),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1774),
.B(n_1709),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1772),
.Y(n_1807)
);

NAND2x1_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1731),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1772),
.B(n_1746),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1803),
.A2(n_1750),
.B1(n_1719),
.B2(n_1759),
.C(n_1712),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1801),
.B(n_1750),
.C(n_1677),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1773),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1776),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1776),
.B(n_1735),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1802),
.B(n_1747),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1782),
.A2(n_1750),
.B1(n_1759),
.B2(n_1677),
.C(n_1665),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1781),
.A2(n_1750),
.B1(n_1759),
.B2(n_1681),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1770),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1796),
.A2(n_1765),
.B(n_1681),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1773),
.B(n_1740),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1774),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1777),
.A2(n_1671),
.B1(n_1670),
.B2(n_1759),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1804),
.A2(n_1697),
.B1(n_1665),
.B2(n_1791),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1788),
.A2(n_1697),
.B1(n_1648),
.B2(n_1682),
.Y(n_1824)
);

NAND2x1_ASAP7_75t_L g1825 ( 
.A(n_1796),
.B(n_1740),
.Y(n_1825)
);

AOI211xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1780),
.A2(n_1740),
.B(n_1758),
.C(n_1737),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1780),
.A2(n_1682),
.B1(n_1707),
.B2(n_1701),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1770),
.Y(n_1828)
);

NOR4xp25_ASAP7_75t_SL g1829 ( 
.A(n_1771),
.B(n_1760),
.C(n_1737),
.D(n_1758),
.Y(n_1829)
);

A2O1A1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1787),
.A2(n_1666),
.B(n_1634),
.C(n_1662),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1813),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1813),
.A2(n_1815),
.B1(n_1811),
.B2(n_1816),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1821),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1806),
.B(n_1807),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1818),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1812),
.B(n_1805),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_1805),
.B(n_1785),
.Y(n_1837)
);

NOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1785),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1809),
.B(n_1791),
.Y(n_1839)
);

XOR2x2_ASAP7_75t_L g1840 ( 
.A(n_1810),
.B(n_1670),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1820),
.B(n_1789),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1826),
.B(n_1794),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1827),
.B(n_1794),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1827),
.B(n_1800),
.Y(n_1844)
);

CKINVDCx16_ASAP7_75t_R g1845 ( 
.A(n_1829),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1822),
.B(n_1800),
.Y(n_1846)
);

OAI32xp33_ASAP7_75t_L g1847 ( 
.A1(n_1819),
.A2(n_1793),
.A3(n_1792),
.B1(n_1790),
.B2(n_1795),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1828),
.Y(n_1848)
);

OAI31xp33_ASAP7_75t_L g1849 ( 
.A1(n_1824),
.A2(n_1777),
.A3(n_1771),
.B(n_1783),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1814),
.Y(n_1850)
);

AOI32xp33_ASAP7_75t_L g1851 ( 
.A1(n_1842),
.A2(n_1843),
.A3(n_1844),
.B1(n_1837),
.B2(n_1838),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1839),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1845),
.A2(n_1817),
.B1(n_1824),
.B2(n_1823),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1836),
.Y(n_1854)
);

AOI322xp5_ASAP7_75t_L g1855 ( 
.A1(n_1846),
.A2(n_1830),
.A3(n_1777),
.B1(n_1825),
.B2(n_1779),
.C1(n_1783),
.C2(n_1795),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1837),
.B(n_1775),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1831),
.Y(n_1857)
);

INVx2_ASAP7_75t_SL g1858 ( 
.A(n_1841),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1849),
.A2(n_1847),
.B(n_1840),
.C(n_1848),
.Y(n_1859)
);

AOI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1832),
.A2(n_1779),
.B1(n_1790),
.B2(n_1745),
.C(n_1733),
.Y(n_1860)
);

INVxp33_ASAP7_75t_L g1861 ( 
.A(n_1833),
.Y(n_1861)
);

OA21x2_ASAP7_75t_SL g1862 ( 
.A1(n_1840),
.A2(n_1715),
.B(n_1668),
.Y(n_1862)
);

NAND4xp25_ASAP7_75t_L g1863 ( 
.A(n_1851),
.B(n_1856),
.C(n_1852),
.D(n_1853),
.Y(n_1863)
);

AOI21xp33_ASAP7_75t_L g1864 ( 
.A1(n_1861),
.A2(n_1833),
.B(n_1848),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1858),
.B(n_1834),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1857),
.Y(n_1866)
);

NAND4xp75_ASAP7_75t_SL g1867 ( 
.A(n_1862),
.B(n_1841),
.C(n_1789),
.D(n_1799),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1857),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1854),
.B(n_1835),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1859),
.A2(n_1850),
.B1(n_1745),
.B2(n_1739),
.Y(n_1870)
);

O2A1O1Ixp5_ASAP7_75t_L g1871 ( 
.A1(n_1855),
.A2(n_1799),
.B(n_1786),
.C(n_1797),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_SL g1872 ( 
.A(n_1860),
.B(n_1570),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1851),
.B(n_1797),
.Y(n_1873)
);

NOR3xp33_ASAP7_75t_L g1874 ( 
.A(n_1859),
.B(n_1572),
.C(n_1739),
.Y(n_1874)
);

AOI211xp5_ASAP7_75t_L g1875 ( 
.A1(n_1864),
.A2(n_1786),
.B(n_1784),
.C(n_1778),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1873),
.A2(n_1760),
.B(n_1754),
.C(n_1743),
.Y(n_1876)
);

AOI321xp33_ASAP7_75t_L g1877 ( 
.A1(n_1870),
.A2(n_1874),
.A3(n_1869),
.B1(n_1866),
.B2(n_1868),
.C(n_1865),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_SL g1878 ( 
.A1(n_1872),
.A2(n_1671),
.B1(n_1784),
.B2(n_1778),
.Y(n_1878)
);

NAND3xp33_ASAP7_75t_L g1879 ( 
.A(n_1863),
.B(n_1775),
.C(n_1752),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1871),
.A2(n_1757),
.B1(n_1756),
.B2(n_1744),
.C(n_1671),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1876),
.A2(n_1867),
.B(n_1798),
.Y(n_1881)
);

CKINVDCx16_ASAP7_75t_R g1882 ( 
.A(n_1877),
.Y(n_1882)
);

NOR4xp25_ASAP7_75t_L g1883 ( 
.A(n_1879),
.B(n_1880),
.C(n_1875),
.D(n_1878),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1723),
.B1(n_1721),
.B2(n_1798),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1880),
.A2(n_1671),
.B1(n_1670),
.B2(n_1666),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_L g1886 ( 
.A(n_1879),
.B(n_1721),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1886),
.B(n_1723),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_L g1888 ( 
.A(n_1884),
.B(n_1669),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1882),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1881),
.B(n_1683),
.Y(n_1890)
);

OR2x6_ASAP7_75t_L g1891 ( 
.A(n_1883),
.B(n_1689),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_SL g1892 ( 
.A(n_1889),
.B(n_1890),
.C(n_1891),
.Y(n_1892)
);

OAI321xp33_ASAP7_75t_L g1893 ( 
.A1(n_1891),
.A2(n_1885),
.A3(n_1634),
.B1(n_1645),
.B2(n_1714),
.C(n_1717),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1888),
.A2(n_1689),
.B(n_1717),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1892),
.B(n_1887),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1895),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1896),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1896),
.A2(n_1894),
.B1(n_1893),
.B2(n_1689),
.Y(n_1898)
);

OAI22x1_ASAP7_75t_L g1899 ( 
.A1(n_1897),
.A2(n_1898),
.B1(n_1693),
.B2(n_1717),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1897),
.B(n_1693),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1714),
.B(n_1693),
.Y(n_1901)
);

AO21x2_ASAP7_75t_L g1902 ( 
.A1(n_1899),
.A2(n_1714),
.B(n_1683),
.Y(n_1902)
);

OAI22x1_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1636),
.B1(n_1725),
.B2(n_1683),
.Y(n_1903)
);

NAND3xp33_ASAP7_75t_L g1904 ( 
.A(n_1903),
.B(n_1901),
.C(n_1674),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1652),
.B1(n_1649),
.B2(n_1663),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_R g1906 ( 
.A1(n_1905),
.A2(n_1550),
.B1(n_1668),
.B2(n_1672),
.C(n_1678),
.Y(n_1906)
);

AOI211xp5_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1636),
.B(n_1586),
.C(n_1666),
.Y(n_1907)
);


endmodule